

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FySm6LQkQ1pXmnt9db9MDo1J0Y0sgfI6V37f+hOhdxXb0uRZEBUgQPHWGnkCx5p2UWv+d6Fd1giy
AUbI3MIMmA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZJche/Nz1jLSHFht4bxHZL+FzmEM4py5IivDzuIGqOtvcXdIogSKR/Qh+CMHHKg167REa07CQTeF
q+om4CFjJPw4usqHU6vWkbuhhqUl9tXU9z404UCeJWg3ng7UfxajdZdGumQ9Ota9MB8vPmPh2bKX
OmqNcPXFu5C40aFaYq0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RO86T5wZ2Pmnkz4qWRNv9HcEdDv5BE05sSzauVNR0Wug0nNMcDDDQx9znRGaflmIl8D2zQqqi7UY
mX2vrPlgl8qYZ9e/c7KysVfjNx/nWYKOt7t+LWKXJEDBCIMrgoFahGqvqnPZKJ5RpueodLA6Cwvz
Toii5JNhp6PJGQ2EUHmI9AVBo1njntlaZccvdYOympPmjsMDUJvcDy0Adq1AynMhoR97wiRH5xDr
tsbyU3BmnJw+1Q3dWyu7HfoArNmQL9hAGRpFhfq9nDMxZ3gmZ35y8IAjfhIcW+rhZDrYxtxMD3p+
xozzeXkjjgfbI7uy+/gsE+tFGyNaQVDOuDKR7A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dV/KWISc9xGeCOltVPF2Pb9Iw8SR+1BYfCcxiT61SkgRi8GTMwdR69SRZ6wVdC48GyT7C8ARpvXF
OWkAYhP4J2TgnbwKhSPn6ct2cqclGK0gDpEbjybSGmukDgqdFzBmiaRqD74fE3UekSSBUq63xYuk
/R7S5lGWxUhCKxpC3DNgQuNBmKJ2v2mDc3iRkjj2QvyU3p9rKMpLugQALbcooKz5Hg3sOPSgC2+r
+uEqaxRpFjyI/69itxB4OWVuwR0XtG9KZ7scjdSMvT30Rklpx+oRzIvkw834fcqLOzlVY0K2xN0S
CSs2vp/wmS9sBq6GAWYNgM3rn0lCfhBXEOWUQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nrWsRH4rMlzB1P+CLGnKDWDKNFOZaNP7zMYSXnyazRQ599AFY17MT3Qto45Ob/RaXWc6VK5zHASp
VJsw1yclaoUBz2jTtYoBLh9+MXRbt3L/Z3xBrweXruJFcnKK5kSjR0YosPG6uDYf9xyHdCeHjSAx
TsJx2uZ7jsDGTMQSFywIrSMzwMDr/GiSPKo/B1uE3GVCWzRUsOyLEdAY7zjzIIi7Xb+2C8buut36
aa8EYS5W/86fYzOea7KUprx+MY5/zJKevWX9/P9W9vywhRSEN6jjmntAYbxTcAV1XFeXPQ1WYT+v
6dqqzaB5yBMZjal5g4r3frBDp3J5HCiP43eXlA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g9fGcDFap7buvVmXkEct8AjKzpCrKIQE2LT1UKu84GxZG/guH3M26I8ynda0idhFABD5Wy9mvPDZ
ZhZB1TiNs5DFq35tCzL3uOEQU+70keod9JF45idCaq0ziiS5FGF9Kkvaow4RUxcwzIBQXryMZu+z
YgNIlOCjEqAKQk1TEZE=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ik3rJlzUoAxI0+INws7w9B9QSkZVhGMhbc4TvgQ/6GlUsAHD6mxSmW5OtnZ37fQfRqQFLSOfUMaJ
LnJTYem8uc/7seaifZWsfyO6jawQ6dQHA913p6AVTqA8qVSgAnpSQAlgUGyUF+9jLj/AnhHWeRIx
tedySnQTai1xfKWIK2LhZw6gE+h/3SQ5l5hNfKvIPMvQrmU0fBP35YE9ebZ3IS18bMuAtd8tFN/h
t9NSBN4J6j0mQRMWt4uFv5UH2B+4w2LIAD3u7yD3/y0122iCxNKIWIhGsCbjl7zUEoaswqCATg4O
Xn6qFvMzH+VFUtMapZM5XLuXKhagCcXDyIdDXA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RvzR1yfzS8587OwTygm++9bAnFwkZrqwGwqMgxnQMX+pouDhihx4vS7qQeV0rPPvgRrum2vAZxFC
cawDHAC0bW5K3u+FCGC0TwMYiz5fX4PRO6MLzwb3Ccqtc2+U48wKaQP+80ac6U8UCb9jD1j6gyNM
6w+G3hiDAqcA5C7vDxNuRvYI5HIKx72o2ZQY1lyqnT4MVgMAMJnvciACsmhJefKoXt0UmYlg3eq0
3NYsHfUd4o5zplRP78PigWD1xAkkspz+Q2uSvqVCTWTZkoCKmjM6P8s8ZRHvWhUq1OPqJG014U1Z
W9eswTkc6YVxYKZg0IxIm6jEaajI0n5ip1HZNA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
TbOw584tzXkaUyYU4/Lg4MF/E59+8GeFs6iODoG6P601SDA10L+razH/CVflMhKyRJFHU/mPzhIv
/78oCc3N1uDrOsbXpDec9e39cC8qSk4dm58z1RgZEEcCNdPhBGZzuiVURcu0ySi2p8rtYiIlCL+k
E07bFOuHQN/DLSt12+M/tdeLnnLPahYWsRM+XVJpz35LLPDmpVGm7k6jBIYjLw6iBzPP33srWdM9
EbB3ZBLah+uL72sgmN26iFFtKiwo8OpeiSoQ55mGJKaHghG+sXEQMwakdxXkDVXUt1kPSDQ2v0jk
Hlk3p6kZV5nngvVgeg/KtZzXK7GKyKZCUXRYflbN6EUUZFLz3s05STlHf8fyUtvU74PEzXt7C50+
/nDP6UtP/WjyIuz9nwxCLWQ7Om6PhFBDjiNG5C1iPv2A5+vF4DLkaveqIBtM4PgMWnG0IkQIPTdP
VeoXumIbX1Slc092J4qBbatotuh0suUuLqY8dvmUIeiojg0KvIOKCn+d/hYkU5Cit1Z98zbU+TDP
QMQnSWYLNR3Z/xrU3wDdifPdJWGnoQ6A/czvMsZYzctClnjTypj9cJiTH5VSwzjLqscf9NHGEYpj
b3Js7XryTyFPQIWG9Y/XRbs+1O16+C/dR2WCtWf6qeT44PlK/cm1AL8KF8k8XPVZdb8mS8KQ1gMU
Jwsq4ly15EGZETogJW2spoR086RTT/4QvpFD0+QyRgmG/lI2PtTFV6xnHUHGowJDjy28j98k3KQC
AMV5PTuIBV87Lk18PAhJKem834V3SyxXxGMr63l7f/3X0R2xe8UhNx94OyeBv2ErkjTc7FJnY+0i
M35SnWwxZD/v+tNgOlKNuWhBllA/t85cL5S0zo6+eW4WN/VQFdqkVyFa2GBywZYlhjykY6x7oxBw
zGGYAV3rdc5XLSqaWsx9xZcx+eWQGXhKhMQd5k9mYQUKQ4laVN9einVSLvorW292rk/Z5+WgqKxK
Sq26aC/YqLCNnqlYeG/sFGS2CI1Y35SjgPce6+YdTyl1+fx9hZmh4dmOvtNsc0qyE8FDI7vIYP5b
Lo6UQLVM78oaGnR84s50XGjHtgxV7rPsaU7MteP7e3OSgrSlC+/Zr9/qF5QCZ9Qn4cj5ejQFnZTE
de2ymnlDaKkleHdp28MqreOWrloTJukVgHk4ZZzfq054cMJ0OSsFE02eZJqB4FphaCKaANXhQxYn
j8+HzpWwzf+uJcL/6kTAzMtJQo5E2tXZ4RR5D9+XzuFxJ67eZ1Zr3dm1gJoGcOIT327Q46BzdLfH
i2nx2D5OlAqUjwmQCdP99G3gg9635EUtnjGPCGMZUeGFGcN5fmZEk1iLbTpBFgJa9Iiedk+kZHm8
h5FSL5XtFoiqAP79VKzw62XTN0xuPU03M9xHp07Nt0o8sNvCiclf5K9R1xN0xrg2O7VJgBLjQIp2
CIYFa2dnqhOa6PIs9rolWmv/u55Y77/Tbyw0tYklcbjAWT0NyiA/3MfyelyKmcf61M1OWS6iO1ky
IwBTnHeEBfeNHqI+VNswlIsBB30c58BFDVpJ8d+fJ6muYv3wYj7khla9enqL1aCOiT0+y0/m6paI
6Sd0L33KGM9fiaRUmYx6D9a1/xgPiD8EN3Dc1o8k+mQnPZg8yi0rbOHrZ/NKShxq7VWblHGhfeb7
CvQJl6hu8mgwg/yz0qpe+FkfnoUi08tedpQZZckDW0V2+feM3pKW2XsQwuERzTH/3n9lhuX2duEp
f1zFW4ntZB94lCxzGuKM1yHcS9ScI/Soi6aDwV43JTxkvDeJbOrx5hg1/W++BijG0SNioSMIHOhu
edYC5JraM4WS05BRS1hjWk8MLg+11u4cKU0HpihHdD0fSITezaMBJMtGW+V1JQrgHq9AsGye31v7
t5HDtY0zefXvIij4sl3XuF6bXBZmZjszOrIfswJlnvq+wByqZ5ekb7w5U4wMPH/JeZ/cldO3kHYk
nmU825UqcnCJwoKOWXT3AnmZCgEa0gwKZfnTmYGTq1jNU/F7+MQFMKWhbj9wYpkZxJbpnTgAS4if
WC9S9fV/vWVLOkXVqxpOohinkhh9/zNWHbhZZC1atnRpCCMq/1LEjtEMnQdmLNdF2Iv7e+QQg7SF
39zuafBRk5M9acFgyTrAEJ1mRU2eCiOLv97sJjpbPyPE6Hk/CUT09J1KRc5BQburpchEoxnBn3VG
o4DdFP5XYgaO9CBQc09xF4Ez/r33Vr6T5L9ozWeiVopUUKDJwDJ7t1uAzSjeVR1yiWCv+Sfe0qIG
OV11g/VBWVuV4pB16ILs4sGA15S0rq4XDslUxgZ0j5YzTOWWD2AKuBDHsGI57hwxmb1ERjYGg/9S
XU3JpFK4Hzs9Q/6OSqbiHzalMdS+odleRkLP1h9YWd7Qdoeue6r67oruXTlTsWm0LD7OnbshIBZx
tLBqQHiwSFM55JS2fm8s/i5qiqVS9J5B2gCYHmXEmXfQd6PeBU6hUxhunOHxsn/d2kjC9xA2VLSF
h8331sSeISAFWMyCSElHS0l/sIIXL3g9kyH37DRjuT21LmyyXd6/bn/Dos0eogdqAVFkM6cD2w5r
UWVeC3g1YJa/6FnviHeb23jYd34OWZauSPkzN52aMyZgwNpL7BS7ZnPA65F1Qgh4vxyRiK0B5gxJ
DGZX5QzJ+EJu1UP6Y6MS0GA3nkAdpUlfzomgN2M6zeqgxEOvnkEknT36Ikzy+DlEWMzJcOYrLlX9
maDDBkJ6vd8xCuouVFLT4R1k0APgnIhb3VLJKaynyAHGs8scndeilBKwh2/PJbAMiML/sDVv0jew
zy0DpHi0B1TTDcjF1/haWtudWTFdojKdMWSs2BLAldv8+MQkIgSO4UG1OPrpyWfAEpGukXrOMd/g
ik40WfsAbqwVrtKir+p4z+COxasg8TiLqP97RXSUg66SO6JoPbAMUymsVyWV1l36FMo/xt+7DUPG
IgQgak7FcEbDTUVl03OlutZ7knXgckE19CU7Uzcm/UigMAV10jOZ0wUQVTJiEVMWR2Kqoq6a6igI
X54/VAL7EFgIJxymT0ziKaHvFdesA+3hzMgh6605o1Kz51aigd8GSr4WQkb/3TZ45tIoA7KIeWwd
hSxHnTcOs2Qx9Lmn76zqJ4higxUgXvdyM7DxsPoucFxJXD7tOgMfQ/Ye0A9nr8Sg/BAqKLEsWPrD
KeGgilRQLaZXzxtuHKOdtSQCfjC0kw0NMuTfA81X6xyIUJskjQU/Y6GpUECet/PFqQeCCnEsxHL4
ckeCA+eiQ1ImB0yLm117LPDRD0eNJkay9S/+2p1Nc0Vp0zd5rtIiTOSfaY0S/24kkIv2d1hdiqlt
N2apW8ZR19QeQdVLow01EmxBM33jkAnYi+9p3bEfZ9qFkFR8ICfx9D8flijDwOrQvUCXA+dZKqxJ
KBEwrWvZApFxrl+FKxKsQxFp6nxvbNxoaTsGcBLc/hexyspu42VRpBCaF/X+PXq6RAXaIiwqpWw0
40SrdfNsAIoes4yQFPY7Qc3ItV3wi2uXG3pmH0ldZ5ZhmVB885Ouw5QRy8WxVAvE5OhAAIeO24Tz
nccugLccE17T5zw+0y06MAa/DgGcVBK4fsinoH8NYIlty09782O6ZATKiytVZIy6A2Jyi3NspQDK
aAUKWFSqO95QgBLZT7xS/ya8QYe8zdZiBH/SwjGk0rYtTgxes4eKhIqBHnuCigyy3meEky1Y7DC0
/je/MVCt/NSqtdo/LFnhFo8pUS7N6PRXQQ5vRjKgdmmQEuUfhfBOREz2tVMPsDehYuFd/ipQzkGk
T56vD+8FKKF4CCwhbHuJQnm37YV18tiMVLdGCtUSKUzhHw10LWJ42X5i4I+NJ5i2Gs2kr7cLDres
p7B7lADpbAr0oIedyGbCNHtQazBxjswont7EA9JDNHA8JOqLKqJ8Yh8PoTApJAZUT3kmwISuiLp+
Lv4zRoetjxsE4AnBRnm9l9CEmbuypUjMxLRAzCmImctfyLqlPuOo7qCjRCCvHF/lsxxSkmYiyDEF
C4ksGlFUpdu1kV58kfgdjCv1OM8luKm0V972/aPzpuXSESlVvFfa5FZ+pwAMwIfm8sMCzr+pc5Gl
vPz3uyT8dS4tcELD+i34FFu1Yoik7U+eX7BIu10ctsZ0aed0wggh7eXsJ0JJAxHCenNrsYV2ixdC
4OQaZ8V88z3yykkzt9DmGCpSAztLo6ABTMvxDitQ+hjgTp0TfbDdSPDj/yer15NDq01xuUffJuc1
ABfsXI0Jza37GnNNfBhqnnBkZrX49ixJ3LA4ix4jifka/gSIgma1LgUeo8rCe/xT7trV0M9CRj5S
VkkDd5sFo0BE+dTPyBGWeefQ7JmuJyy/bPVwdMu4iQZMej8NzkMlYcqK5G/VJRqWvuQWh7d/dabL
7v6GQjaamxp6K1yvVcy3mHwfbqb+EQRjMV1zv1YC4y6KO/6kRKe3iH933EmcHqH4NsxeeBv6xkzI
tMBD7NY/zDyLoX8hlhHnqjC6W+p6PXccbFjbIkj4OiiE4L2yNfWwiHfNxBtcTZcgw+j//FQfvtwL
TO1sNySp/BQcSYDEK48nGpywYPjLkuSJ7SjuS2Sn0nQ4ODmrKZpV12h6q71f/dEtb/wXBbfl7XaX
V8d/nC/4m5EPelg/bU2ZmVVEC0OO5B3AzScvn0ePs63BLAR2ouuk9uoCvKJjnno6g/QZdAXGkN8o
bxwZa14aWt59jPXju9vReppr2SkpV7W/FVedP+a2EngT6MabCaIf7rpl9PcfFgQ6MpXApUD21WlY
zsHCT5qpdeoTpXOYmwSW6/JtxcpZhESvEZq7VRTnEvBm7WHMEhgQcTcSBRaPVIoqwx8ds1SVFMip
kL8LR/3PIQcXV02focRu5LU+65KxaRO2mNnZGtMKPH9RycAfIufiz8KmzOThEov+vfvseu5Mht8R
gYxnNrKTD17c1wexNoaFy70ZeD8JUeNjj1knlXkVn2H1V0EnMvjmoY6hdXiv1H3pKFghH4MH3ckW
julrS7vkDGK26cwp7iUGMh52xbdLe+iIcnkOyk+8L3Vf5NEpkP1wBWACTXsRTJfec9l0wdJ+ANyw
ReFAq/K1YBinCLPDKnRguF0DF4dKd27X+b6lGSKhnAofUYaty931DCC97stZBADZr4P4MDTsGGzv
wNgOl0RqV76fTTREvgj2OXvrsWeqofcb9i9QpEJp8QYRFyvPjvnbrY98gQkUrcXqG6Dr7yNx3VQu
D0zn/WpiPwOiW2gL91RX7Iao1W/QwEB/m05W9mK85i+oHsIcnaPagjt6QkAVa1a5/9yhhFMV7p7I
3+wyo4PKU/Nk1HMiISPDzfGvHCtpLWlgaH20vzLvixoTWldjcoa0KbNkX4BclrlZFHyr3347JvgX
uy3ANgCtAj6bqz1fkD4J+aiOGB3/47BhNOl4iiP/s+xadGNTSKfahV0sI1NIh+Bsd5tYWciGCSLw
eQTUm8BBQMgl3F4CXJGw6KBvaAoOet30OCI1N+P79HC4vbPLAvzjLqQfUElvkV7V/sjAsVOdAikD
rJQo7MrQU79V0+4Wvpa8rOaDMpja/ihV40GgDeA/D97pkZYj3niXOhmrKPfHiooXKhFSM9JuBjOW
gsce5NFObbi9FvvBtfTbzhiQE1wGJcoob0HjPwJ2s3L3g3JWyaRXUqeOlR8bh0YHg6geoYQsOM5a
TRVx1/DQOByCd5B+4l1nFlk7HK2MbTR48MxVODS3UwarJ0VyhM4mXofrZOqo2pfF3+yH01Ve/MV3
/H/vr8XYS3nTeheUinwcZDCx2mORbOHtQcSeFwuUTIMC9DORnV3LClcFYcV+gUM1mRSm+OYs0x2F
gBiqJ+n8HuPPrub3//3HEXPpaw1I8Ya8ag17Y/iJ18jac7/iQoajxDVbnM1FhAcqTGGG7M+aGKVo
kuQGtXAXp7AVFJtjddeihHN2Tn39GbvbnlDRzVJenMSOrTPh9rlYuIi8X+UQAs2WyAujPuJhskEw
rF0UkHSdXVvHwqCkwBP3LTxwXVF4Vz0M8h4F+0yXAHPF9v6BMrvS7HFv1nV203MH82S/uiUdLt6X
YEBp4La4NVR+cKgifhFZEfptO5guW8bK/MMlKOFn1hydyK8FzjO9olejUvbCnJgGecddcjFkRnD4
JbWyVEX+lr5JXLr2CW97Edyrv8w9ZmWGdcbNyzQSm+2+M12d64ZOAXYsb+LEpdndoo1q3Y28JCVw
a631oyWxXViQNEBbbhk2yvDnRCYfmYWWdPoJcQp0S696zHE1YLX4v0eYBsH8kJj+nfr0fahm/zPs
1asZZAKM1eMfufu/35CYCb8BHHU69n5bITK6vwYhVQTUTxNHxfv/nGiaycN1Av9CemMqKTV994g4
JnnWZOBFPTe1QpiUnFfnLFoQtvVz0I/EDttc9omH68BHXWIFLqPcff81kTW43VthL3ocDe4Wg3w2
8aZtvJlJPB/sv1p1rEorjxmBuWOPhL+rxlVshaq6V0aYqLfPhW4mDHmQlKCyuVtbw/LZtHAKFfPB
tpx9m8WEQfmeIfVv8iyX7Vjzw60VCTCJ1Ottr++V5/5BTJ8RWyZk6pOP1pVgFjUL1TarX8l7IMm2
GRCrK9/Lo+y27JfRudkA37kHiuvFABRgT4S3f0ZOYK4OmaCmg7L3XolkBwg1lIZE8tfDH7jyWV9h
44BqmtujeB3cs9YRfaCme7xL3/+5gayzuet8dZS1Wc4ek+GlR2TJTDVOX3EWfr3JnV1bT/BeWfVh
Hufv7sEe9iXh1b4MnKBQozMfRUf9UYi1NpkYO2m6JWe8zaj+0Ma4x05F0dVHoX8qjIPgc/yq4wov
jZGvGmTv7Pp2jcTZTJgKr8kGcX2BXW63X4ReCW99/suNs+6tB4mzHTeyClDLMBfxrIvvqiu1C5Mp
jfWWRNt8bQ2S8m/gZqS7yAKLYqwkEgvc+EI0JwSXg8ueTWIP6LC9CxIKfNmPM9FH8XUOJnyhH1qX
pZQP6NTCvJbNPnZowVza30oci8hDft7Dqn7xtiwfdHZHZ2b6INVCEu4ykGgstMdDHd+Rc6GatQxR
Rijz6qXE/F14nvGJhopkhjBa83AWO9Nim3NeV9KyHna4Tp8iNnBGQtneqbL9CRPln8C9D2H5R0ty
HlBoHeAlTMx7Q3idNUH3L4lUtFI6jJiv2/5wYZfNLQ0qK5dHgCKGJuvkeqrMieoEqn7wptYzuzib
1v9+UeNXjlI5VpGGFfh/lYqo2CbZmvjw+crtUuqq7LzniIDRDJcVJU59QHfXi/DbUeawQGIzhNaG
0BS+b1bFm9FJiTQz5IDgIJCLLxvW056j+WNsyH4QETE+EKUtBFIGQQo4zfYk/0slDkAK7F4fWApw
wTi0Dys1LOLCk6Us7Xl9LrmRXWgvM21YQL1sIVU2dKholoHLFYi17uJ6UX472lnGPzcqj2FE7pxl
3tzLGJdapZfrq7jMxWA+mVinjmUup4DF2/nWEAmpm52P6XFKVDy88fli53Q4UEoEJMXOLhWL7Qy3
1PwrW8ZU/msgfR+D4MEyX3Rw7k6IbeByRd1NpUgABs6zqsRU4A+S2YYH8cNU54Wr24n+mp99LAPa
5ArYtkNN9RIfEinkcdqv0cP70oV+QV4bYVUPxtcgOtaWeVwNA5fvStazNnJy2B1sOQZ5ZZbAHLoS
rQ6cp8fRwDdig9ALB+vGoQMDgQ7fWIarJF7cddbXrWj24aN8yFRk0Vggg5uk0RmxPKxh9jgKr6mR
j9tEYC1/UPGuPPoHCE1V6WZSIPo6Lmitp36jkeHMLeHsAw2E0ruAv/Np6FhUFGYmh1sErXFhZjO+
VD/sxRgSJ1ON2hCHWhZnHRpXRqehREwZ16Mi/O4SOTc7kSNORjyVkLUdgWsFNQlKPNgpwW/0ixzx
XZxymgaQtSk6KG1mb+aYDlwlu5ID0+rs0KhTD6CDSvMiN6lmotphW7dWoP7w6lwgILa1Km9484XF
QLWLP8EzGMq5nLmKKk27KENsjaEVceSWFopOg2x9qi9nXosrUxpEBKVsaGKfMhNy8RyDhCn9BXGO
ZEkTEbKyPrvaOIvt42ZTGU1ubNxfhsv/Gm6msTRo29cwEUg5+HafPtRbLMwqXHiflb3fDylSKB6A
v9yDuXsbvDxTJuomjcAj0WLdYSy1YVXmvpO+jzCLDvJ2SS79TvIkrjTCS3YNvcSTVupNBM3Qh+kW
lGJuZtkY9DjchMwQlXlrZ3BYxh2NOQ6QISG9p0Slt9apzi4JR3z2oaQ6jYSvohDhXUzGxyGv5Vl0
dG7HlTSY7Ut3NvDzwnucNdo7aoeZd83nO0nQqowjwsXge0OqmGJVFXKc7WrnET0/+/8JUkyP405i
xvAAFXWYMwIUEIn9EYwYq7QxpyQlQpendWUv+/iILnT+xgDZcLMxIi3cSeINTaWj4eHjSpdwALia
qwArYCSN1lrLyaa9UbfibLWMj193TO14oVpEg6Cb8+Ggr0Z8ZjkowAj5+m7Pvd74rmnb0QFuJhWr
wqlx3ppjy9OMtjA9Q4SNQGTOkBXaW83DYi2ULytlFY9rBXeIvVbB5YwiXIulAlSGcb/hiC74lZ1e
3YE03G9hGq0jn/S8DIUVP9n/02SxTMBG8ljx848vTjvRBMZqTnOBIs58H+TaisUONQAlSoB3VW6h
bwsUDkMoKg2lQf8vlGEdmKFV1DCE/eOmiV6i1Ho5kQF7wHM8kEsxPzUuEhBbO9Z4iJh+d285xjvG
s3cXombb4paDKjvLthSQJq8XFbeedRsM08vIn3a5IahEoJbDlzte7xwhynDkD9BGsmZNpJwXnNeK
G39Oft6iuAX/B5x0zuj0skgDha6U+arkRlpYCYlgDBBJtKxFrLy7nx1jaoegkS0SGV6qxLQ1vef5
ByNZ2HHHdGQxf1HMgHnyP7smtJVaO6Uc3kNPjKfx3ufi0YM+ah6pkAgwfeQ7R5PJglWOeKu2bUa7
sdW5nm2f0JI7g7WLMyUfDgAIYkVLE6/HgxRjNJCSku4CfB26lmcXuqEec+/4lvST2Plzx4dVh/jC
Yk30wctf1x80ttj9ZcQHmGeF7rHHwyFzhUpmZeN0F9x5zn3lPSA/NAtAC0denxejqrVsslHfFkWk
orMXApyg0U+3tLmfim4QpPWcXoEAjP/CJQWmbidqGobT346mZ3dzStfkdZfCIkV+PNWfsFHe669P
9+qVD03xhR9ymOjyqvT3nj1RPkYOv9jBN/BJUFEECnLEr35yj/2v1KccBN6MjO6NpxG+/Aj2wrmf
5Pic70vdWlwlOzNHeOZBsxhQlHccEZJHgXQVb4Ga9/zwB8nY5PUJtR0nKFlU6gUHPdtwrVpVuyio
J1BFeDkiiOX85bY/Q2wdXqnO0xwJyLstNVaNt2gqSCMl2n8KERX/iNo8RWse0Sqk4jpOXgmMVlON
umEu+V4nqnBlCNww3awfLhg3X+DblFWg5i4skOLFfEhmlB1Ze8H75T8BfazAmQ5qzZ3/BJSDL/pX
z5MCwTqOxWOGWf8/atqvZng/J2YgGr18GxGHx05d9nxiq5Ibu+aVVcQPmyx+AwMHl8FvFvDsP1zP
HsXKsabhi8KXGgIhDMjs+ZEa7/jdSxljKzOtbFNeUvU8UF279/X21dgJk6Mn9hoiQBILfQhpsyHK
6RIP6yJVMb9+ZEmZBdiL5HovLXHO/sz9dENRRboHxVsLOftysg5lhSu0qkK6u0lI2DVhoJ7No0fm
eJ8I0b3IdL9izkrs1kOBDZWhbkOdp/YaGcJnV7TfbLasAWqBHpT5HJjHj2/ZoYVDhnKHUyfsmrwy
/u+7NKuWUmVp2Ac2vI/d1cLe0teRpOZAVPLRHnyYdUsuam2mdlpOV96t3KNlHRnUC+VCdUdy4Atn
gtSfR/5IgOTkZLL6GoeeUssEw1QBSHgv41bnLMkA2hTwqfdVWRlee6VqhemlwqyEwHE3p2K6Z2IA
l++dWnOzGxNXEaPqTzb+nH4XKSDxJVJoSFnFEhQo4RECJxF2btCOX6CBSP/2Qz1shigTtYBUO0dE
NFldRw7eCoskvr2y9HEkRDv6XraYtI9saPcntQUcMSMwVfJB5SPzvl16IKsVq9Qgo+EiF/L1txSH
9wxTTpJXcFFO2Egp+QBRQaeC5VUR50/mk7aJ6WsdgZCBNTQt/dPTJy2n2ekB6QmeqBOQEK/CT43r
3a2U1XcTR/fZZRTEiuLRS0DiZQVgkuAvNQsyNEetp0soRQHTAo8BwzO1/hUIAEw8cNS38Pswznll
a2kHbJzumQ8vZ530qxecrqA0MXGecXZ58MNOdsppuIdi5R1HO0Cv0ZWivMuuKa6jo62SWPfFvdTb
qJfuYkRZQ6v8vRapVcB7WG7MUoYbJ5tYxh2vO/30/yP0ERndGwDBiURstF67hCW1LHFiNTglILD1
YvBzjeCXsgn8/e5JSdTf9UGvHQqmSGa2hDh0wH49mYwMAkW9lhE5FDxZsDq+2JZn0jQQIxU8qkHX
fRChUD0RM02IHSlviacErl57C9gHPhDHn5DYjE2qUYfzFRBt1x9Ylo+B4EpFBpLrGFSDxpWWKsZ9
1u1HMaMpQdpPH2aWpkIPBDVF115cjtQwtPdYKPplbGivdcGOXXjW+sPQo+a+B9kWm2ScPsyOY2hA
ifTqqlE3Wn6essfGhQcDysvBeh2qjgm+8W8Vw2L8OSpAMFY9tGfpacCbK2bIH944DhqoLupARQ0Y
4eu6JI45Y3Dm05gRp5RvhqQUk/8ABDq3frKAvjL+Qql6ZaYEfxd5sILS30VfHPOn0i6v4d6RaV3P
vNkQDkf1HsCoeC95QIJ9JOApV/IGq0Tl2/WHKlXwi8VCq5q6TcE7yqoG2CZ5TvaFZIoduUOUMgaY
xvTvPVTN00fbNsttXZaaJV6LF0BdaX5LKmhItrVXfWTfMA9BU5ZLoMD4+t1goHh/Det00M0iIAh2
MtTlCMrxarhad/Y+IRb4H593Mx5DGVgX/45+VtZHZCE29mJimoPfHpy7a6rcKYCL/9SZo2TcdBZF
Vtg5QZliQ/uS+WnLEdKvuZZpgcSBr51MlUfLFQxURbiBFxiqZKEa8052Vl5nejP0dQIhyiRkTF7n
eXC94Rqxt/0LhzNfS36aeHYM6Y1kx0lGDwzISO+okb58Qh3wZWaDEBncljrGFBo5zF+uSuAjzVP8
2KuMo2+QNq1yKSj7+lAPlYgXBkPHhb4Ndjk71UMw8Z+lHDzRqayP+cynS/7UpqgP1WZlIWUzyB5q
RHHipxcRi2fsu1OFsEGjDnaJ7uIaF3iGkUQM94/wG4Qt5XrmXZw7WdG6so3OrvIk/lLhMDlpTiU7
Iu3kyhBhV5gpaG0T4CINkBxIieExV4RUd/LOcPUF6Zgq78T9JzUk66pE4hk7I0D+g8VJVq3sllb7
Tj57y04MoswGdiKloHwVXpv+MMUEnZS8nawvUaItu6s1tPVBnk6/p9psMuAN7Iem9W6XWGyMvWWw
saw0CDo+JJrziIWMIh7n1rsWLW4DnBWlvR7phiOcPf84Fh2VWNqCqlXt+14UNdm9eOEuT2Aud6b3
xz9yicXN729FmjXvJMHM/YEdSmKIMR81ulUYohtteu7diquOoFuBHUoukP4TY8m8lzpZDYLn262B
NjYvwWLT2YGZA6w1LMXo/DoBMKyQbr6eI98AXbZ7ynrhYjcB9ZP9eHkp/gAc+BGL5fmdU2cAu8aK
B7FrR3Zsp10U5FnNH1KjEa/BXyQj4GuTtFQoPspoXw0f+9+vdAHL4gJz1qhs+4wSvQTSkBWmCdw9
1s63XWy6RZT+1RC2CXZ7NXtj/g6ExLs2bX/h1go+qB6OTlkCNE7f5pbNHKhkQcZUJNPA4djosDFH
+1kgUrPYgZ3KN1Zy2eJ6Hn1B6U3rkvEpqhKVM3CszCdNTddySUsZ8F8dJz4xo2OoyZEqivXv9Ggh
DGX3/Jjgbab8Oglq2FVOTxaJILYfVxw2nP9sIr4Hmw7/1qE6mBLTJIvRP9mY0BS8M7iNflAWwb9F
KPEHbP/AFoYBEldc9Qp21PoN5bCnTmr8sDkqCQueC3vclusmBkV5VsgtPZYfdAZlKBu4vNeU4nPy
O2LcHBMoYci304UDXzYlpwE5kZiYwEAjn0spr5N0qUB9akZUZ1eaDJ23zi84i4r3ed1e5JA7HmC/
JcE5Dlo3TvYNVAWwSW2rMTCDdCWcJJQroBhVnZ2Nisv4+HU6Vkns5t1Di/AJnoyEnp8kD8TM2qMx
1h9GGFsuX4+03WTH11/dtee/e12K9I9sgYAnEuUxhUEe2fwastWIESKMixq1PKAmqM914cJj6svT
6LXQQ5FjpEOEd0lbNaxzket/r6iHulBWFJz10yW4sN7GtzY3pX9a3/xnsjYVzhjJVy4Isf28LxLo
hFKRYFPSHyqzT9ILz83WzkIZmqV/UPatJqiuWQmLUhU0ZDV/Z2H25YDpdvKmKWHcNjAOaEN7DdXW
iozBw8vQH9g8gDHV7vUnJorbwO0Oi+h+0kQQ/y5DpjLnhTx4SuK8ixLMDq6ZagH+uR4OSWGP9S47
p9tWa4w+qpqLaM32kAor7022QTRxNLUnH9mezXnLMy96XoeGjrTmdBNH1nTfbXCbexmUOhx6cCx3
OQ9vzd5upPoz7StaBaS6gGue4D4Ovy5kIdV2o6JrmctX6xJ82nHQbWFc/HmrseQmlNikf/NK+Y9i
Rlm6NrmPOIqul7PjheoCpK0yf1uau85H+FCofB4ZcWLcWQKJ+bb2Tj2jehj05T35L4zmt/49+dXf
DoPQfVdA9AZf3XwEWOsmB3a60mHLjO9Y5STO6ON4qpfQR/yC1iTq2uvJBa4sq5SFAF2ij3QkVbmN
iPwocqn601SubxrLVN+3uKLJaeonnSYJglm8tW6qPJwg5z5AaNe8jxiCN+OWQSAwcKcbPKhS7LGK
zmKQUBFl5PmBR+W8KwZEg6+iLHQhmySSdM1yllDWy98UrJGJxbBmcFOpgK77kIHVXu4N8KlMcpum
MQcMrHhvpYbvGBMV2BxUs0CXiHt2MYo7ogWtMsn4CcayQqhz7bNivTrk78sOzOawGo7o2CNNxx6E
08nEFW+KYS6yvJ7VtnTorf0iRIXujeZfgzqPVHF7WwgNKXWe1uS5dLTDLI7MbryTs3ReeV/163RQ
CHNtQGWWR7tNevQxrgWtd/OIXjQYg23qzVr0sC0NAjndokNTnZ0X0DD1rClJ3vqRlufGw2ynVhhi
F0bYWDkMYwfphla5dCHM6x9A2mQhYDpF1u1ri1wGe2OqJOxjI7BcDng+DMewRblduN66ipgI4tcl
/cQR4OjOwSBJs7bhqbUiTbwk1W2MzQ44tIyWpHYeJ004QSNYaVfK1XjMqschm2ggxxLPoaX686Pq
VxXKyZX7ystWZa1MFEPcPZ8S/LljaY5fSNUyv+xdYFeClC0yKDjEzJLAyMiGkqib9UeYg8L1gn2L
qhTzuQDQNRI0fYcI+4VUID3neAbXA3MGgF8q+gZL1kBny410E5nTwnBIh08iN2ksVx7y+R4nroVU
tgPsOeWE2FTpdFg10feGu7FWz81iaHOKyXR2d7CuFwRrVHA+Gk6QO8qNhdoTE6wXw+78m+IJSDhK
5iTGhua04ZOtuGgkzSpZ1wU2pEv4NOfCt/8C11rCBFgWDOd/UN97lneXk45SWRIpo9viEi+zb65v
QMvdrvXqe4U6Ywmy840mJKuamXynBiyjNensdLJWdrbTxYQJU3Af4SYhAQkgaEwiugQ24eOvFSTn
MT/dVogMlo9w1uAOJb+a8xc6w55UNmbqRoHphD6K+7u67Ng1KwKbkDP0J0XL3+3oh1z+jz7TlMIS
XzcyaNy4GBZhvdqx9jWckMW2E6SKL+QRXhvdD4iQ+BGmWqxn1SPZBh6mO1KHMlGroe7ExIypr0rb
rnhxP8rTI/TfIC9yCzbJzUsfj5P/pv/F6DrUUBP5GVsueSK7QATdq/TqbMFHURBxx5EbVNw5+8jO
gw7Tw4cve8crcXZIalGR5BqIyqP2JBdIhqx0j7Ag4tTjdkehe4ns/l5mWXwnudfhpeIxuiDsyzLt
cnysn0dp2eZyh4WI3IaDs7N1rFVUa1C5CZ5EJosR9x6McZKnNXLICHrepaVedFLZckIsirhV9Td0
TD8EvqKpI+nEoyVmSqGJzHO95/Yu1+/BHpmygdxQvitBPJPtj5mRqP/+2qlfuF7L2W23bP7rN1iv
dK41kwW+Mcao5+4QUVjuzMSLHOesq0NzIqu0MkfdzDwPRZatMvrJoQI0aH/+k6E9yx2RbITiTz4L
E2SViaS3a96M0EJxzI0AY+m9D2Vw5L7QhL053OKH02dpMSgJgb57mAAn9P+jJQC0/ehuq/GmA7Ki
UY+vvwVqaWxtVmnCX0hGtZ1q0Wvdo31FHglpdyjlz0b37iMODacpiDo9UaYK9pi1XKdUOi8I3jIR
UlUX88yDr9ExJUJn7h3LmlVnd0cnxd3z9+gSpi1uODHV27lTYNy1BheE8Rj+M1USnaRPGDVSGNat
OGmbuP9eoVOTWmeaF56KKflLH4CC60k0/GJirHFNA8WIb4Lnu7knbIf+yRwypX60PVsn0ZzRC4J5
DqsyP04owoLk/hnPVByGldMcRELcbowqGh+zkuWL1dDniDaFWQIXET6NxFY1XoCn/T3HabrDOzwu
QbIhdwmk4l93jbfvFHkX0CanwD0UUEPDnHnDrPlEU8iwG5woZH/WPINnF4KHA0YCk/ts1pB1cuZU
1q2mRZXJ62Pcl9koussZwuXj/D1EfI0moB0KT58SyhYxQyK9SXzOSGLkcV9Ld7TBQpvrnYxOUGW5
AUZwWwfE3swMbnoxQNI9Jphw8IWKnqJ+6Iw138w9MK4edZdlXiZafv5/fEeFs6a1NzLdL+nG6c3i
jVCOlXkCx3tRE64DKL3Hu303zKIRN4mlAa+0Gdtd64iywXXSdni61BnMa6057wTv1dTgFqacsK1w
+kxw5mBN00Fibmp7K4mfcTQw9v1/Zc820hosa3lBaLQrDmkP3sqJXQhH9CQbwqgrPVhyUIUUGGA+
tht7JJlMz+mGaYaULmyETHEyN9ACOQLqLOn5SJHr1UuwOJ9Abudpnn3LfX4FfVpftdlbUakD21wQ
mQ5NKQyrNLau/g9foDfA+ZlTn/K+xAdZeBv8EF08VYURUNh4PiWSqWBXG1UiYW8iE50cAjB26AQF
QiI23tQFlcRg7rNX9G00aErIlVo/g/NC70eWKlwcJqVNWlrfWDB5qy1qTU7T8u/p0kp8wdrrmqvq
Kh47PNHJvuBUehkh4yGPji20E3EIIGyQgAszIDAmYFN6Uxrlsr+STGnhSiIDF5JYsYX348BseFib
Hsg0wbc45/Be/uW35PIh8kpsvdGrxy3Uc/T79rX9tHtw9nUkndEnsYo2MK/Hg8Ny1Z3rqNAzRtvH
b6QCx4wIp6WI4vSBGNInfSXMSJ/JyCNAaZ8Ubn/g3SoYERtb1iMjWfwOBVJLaJG/pb0JFQ3SYRON
djZPNJw99XGxP5wzc9XcKSF+WVDm3wj/p/Xw3ByxOyti2eVA/cURlcO90/XEi5dTwUhvqbDzdDKB
0HSnvqobcXIj3U/M5ku5YEkudhwfpBYG9rYLS3DqbESjALeVwIjlYDo4o1fHSmPOTBgBySZGqpe8
co0R/mKMDoXL2LVSjUrooqGfSeUlHyzPrVjGL2p9Sj6dWeqLK3uhU8xtVCQPAWA1jAHUAY6k+Jnh
YyWYz1XxXoultJyHSw+BCMbAT0jDLxQg9w7JTAmYc8lfDzxMy6Ubq5K4VowjwWqZG6a6Jt97JqFa
XZRlo1GdF/acErGNyPeVYI+f+ILca9UNkwj6olFglSGNks7jSHAQHiPntESXaAPgG3hRPAXQEFnl
WXhUEBefLIiIzUdRpWgxjdfjuHKbcmGGcwiLPZ5TzTOJ9NTH/6tvhIT3frWntBbN6R2UWCkgbGpX
7HOYgX5eqym/Wh0+lx41HXpmfpY/ftEovA3/1tz714cG0xc/XfhlC4lJZPRLBMYFBBonf+C3FB7O
y9IjRq3sdUuRNXvzX51sI/hQohMITO7cLv6oMN3KCMBV/hbfbp24u0veoXC7N107kW3fVe16u9D4
YlyZOM2wnCuIQJ5U7siaCNe7oLUjg3PzfYfnI0eg3AUQIMxfKMtV6PKdAPPP3bRwLgeY2nqG89Gx
xhHj0KVZ0k4EkX9KxCxJ9Q4Yv6nD34FUkt301M12nGoJJZ+VdbqTyyIfDr+EMZTAC+D+1QXCeZG1
+IymZhyY6vvdrly45B2VZPpJRp1UZCpcsAdjBs3SVWplsVju26Wkmd4z2EClT/GGoDiq2QrscyiK
GIntBwdz/YAmrlXZp9ocrsdYCu+jjKt5T4CCStPqzIN1DXjQUI+O2fSwQnaG/70lAcbi5fHDjyR5
ArtDleBLDKzL+wZjb6815QxN+A4JG0a0pKE1mgX0N8LBLKM/iV0NaMlc5heBOvobZnjL2AQZdlOX
IamDivc+yzbTh/n3Vi+B451Hjou8PsuiNSTKyO6IZyBWuJUOKLj29wYD3e71zdQM86ljSHKUEuxO
Onlqq9PO8RYcW62K//1tF7NlZF+56EJ4GwESv8YKIDBG1gdO8QGNiyP/sH68TKFL6cESZvIGzOrD
U0/tN94sYL2AGqgoS4rDUR8RFwfGSkDuCpYMQ+iP9kqLNm/gF6oHnhyRLqtiprIRDOF8CLtpfNs1
WNx92SHmv7QtJ4NbV+u5MCkz1FdIs+F/CMd2++mrCef5oLR1J+t5fL52m1HbMEzLEquIc+CPV++y
VSlpTFJnqU8sNh/9tlqdCWllfxL5Ca/VUEGXcVOy/QJ5IkynXd43lG4LurqVbqz0KRh/C7NhT+cJ
J4VzcTNglcvjLOQhUgSqUoy8HblQNOOy3KhMLNzWYk/hZvaWJIZa03jTZSxoackkQXfLXPbNSz4W
QXpC1NGCV5M0bnSmqkYKcWBfNyznSLr3J8ATW8lvyaMyAU3SlRHMXWUKRlqc4A9b00qF2SCOWNil
wMMT3Yf16DK2VD5EXJGfSdlaf36X2WEypbODF4UdfIv1EfkQNcAhH2PEKLEaJn9kT8ZQ1NExSuFs
2BSgz4X0IPj1q5AefOpULOkMPpF9yIJtibSt0AN24EdNp7ojifj/5lfyY5GBrg48BzFGfZRHTWWh
IapL3Oy96Olb0ThKzdo+XZDGr8sF368dNOjYBbhgcfgQNhKXB+eBISzesFnInrZuLVqZ5xT1m/xo
0orcjIRBiojZLsf0HxOrNQkGlZpImmwupwyBTQv+55HtjtBjxWROTcJnujPruyRTcFJ/uxeCUSK2
142lz7dYRQHCDeSwfL4qZ2wDI46fPNmTzUrXJdk2RM2XeqToGC1JC1cK0Vshk4BxUI5SyNQDv439
RyWFAiEET712e/WORICcFknhGrBOper7b12dQWoja8xpRQuvWf/Wi/flFjUvgGeuRxJ4GXkvNjIe
JiBkqjysCFaGqZRNAKNmcxwH+aM9Ks/X/2Gb+bawDuf1PeDtAJyv3TdtQO7ThjmIRRhoo/CyuUHn
IONOJunFHIKsZtIa0bGZN0hBYCkDUoVX+n4BrWLdI5hOxIcvRAiAg0KOL2heU1tgL3zxWiTb6JEy
oxUJuEv/08lpnxXXYB1bNSIUgC4TMEalkPZM3DYrZqSIuyJbsnmweQOeo7du0eWx6d+bWYjF/Z+Y
2JNmEFSmOGbsX94gK0VRkkb8TfU/G5Qh45XcDvf6ffWotgikE4XxzIUF4kwnufUJh37gZNG7oaLS
pFHZ97UfeqyG/aG13BYJHQcObjAPTh3Zlv2x9Qm50Jb387MprJ3Q7NjV3H5O5h1ZsIvkPE2V1UV8
Ldlvazpu+SG0iyBdwfsg6+sO0CNVtkPUiQyIfSko3iXskpue8eaaXFOK5bEZY+LRq1m2sqCsARKv
LL3VytsKt4egKym0+1u8mcC47NwdADI6Ps2i3wpb2MEQgzlWM7pzjSLGPz5LEhdtPn2U0nKj4+Zp
iXFKyNMXhwJ8RuRQ6dr/p5z8RLLne+350/8m94wjIzApGXKdyty1dOciyyi8PUPB4VVBIM1xaQv3
3ME7I4F9qRbVHrezGAgwE4h/givNzbq8RB559N+aqVpFHFAQCIGps8c8BvfQYEe9P+QF1MMcGD+x
g9n9FR5owEtGL8+WN5bWPVQNEQqqF4+3L5o/QPeEqK4YHm8c2r7nhVqTUBWxgptVbGFfMomiwJpo
L6jFiyL4XywIsN/91RFZ4ZOqZGJLRv5LUf4xGcGFk5sNdn3XKBMOMmerQTosRDM25NnIug6R8k2N
xPRgmNPE+HC94QUj03RnxdhR9fWF9Vhw/JlCQ3kbtg9kujR6NOxx4eQTj5+F7YtZwVaG0Qaw+OQ+
oWn2dJGABq0ypfFOBMbYeojvgY6/cWzlYyWQQNcYMQ6Ga1afHeuyCr/Kfdx5NCsCC7JWN2RAhrn6
ybFHruRpiiksY+QJW6K8eXN6+diuCR+ksykqD4rxZAtsrZNbJMSXmgiPCeLDZFyT/iLmDSbTXPmi
3fyKb/KwJnvDa19BxZMCU2rQukY76aqtW5449UJqeiLvMX/pV/DIia+kB10FnyOwkLn904+CRqc8
+CTRnWkcwnVzmOhwb6ROVb3lh9wWKxGG7pKUvLe84Xsb/fdOWvsJif/jJV2t8Dra6lBxlPVOfX15
qB5l/aYMV6PCI6H0k6vkHGtlwY0Oe9AGdKCmSHKrCPkFGIT7ynNhqvIhOgt+yEKnPdcL9PfvEbhs
D4rWfpICDgWIsWugLepEPMlJLXP06UiXqyNX56GJgh7jNzEgVCaGQXlVoGIVkAyczH0HNYcYRbej
qn90VywesPjymHxgx4a31muDzzxxe+SgMKzbksXZtngAU16SXPSOm7BQB7c6ge5hV+h0/8aowGSO
Nkm2ehkAreu+ebtjYfaLWiC7ORICpPbpWRV/B9Q9TYYzM1P22azjJJnSMk8muGe9xwKwZqmgM58F
YVp3e5GxkbJ3NL42tlnIm+PXGP1J9362PCeN6wmW3neW6Y3uG544EKblvZ60MxrkiwdO6HmqZws2
dCq3om4N/q+GiELAAF1YkOM/xmlCfVZFBvRvlHUZwfqvJt9rcelQfly22Fv0ZVBBlRvcdUDBR/fv
L7poMF66U+Swy/GTM/ZSuTGOrG7VnozKTr8IlU/pzJBOcqs/0zzdg2aow6XCm98+GhTagqSUuxgu
F3LMQNk51OtIGPWJcYd5SCjkOiD9kh0SHrESvSJTkQPoDsU/lc3pcvZveB4bqN1ycRngOc5+jYqD
I3wPcJGyRTEwWvxn28RGIHP/zbt/kwcEdgJnjno4ZtgxM6wLgqA3ZIN/TK7XPNTN6SUirobiRDiW
BnxiTpKcIEDf5VhFquwXqnWXDn4kNKVCPbfh7qHgvvkUh4w8HE+vc0QDtx7ry6OXBAq1Q3yP0AVZ
69Sm5xGaMumWjnZ8wu2UFrmG8HMRlJaMjdKF3Qs9xj7Js7ADgeZBvKa4iZflBinK4c0VXjDRnI3V
2rtKMdFeZPzG9LdB0yzV4ARQu/7aD2KbDua+U5du6HnErnE5ibjAJ9p9RcNBBLImQVSrlmMm2wha
0P2JvHM15hePCFGBti8cNA+lJzp8B+Fo2lOzauicJMeCg/LHMCq0jBqb0bvdfi0qAuQcMSOxb3xA
WefHL4bCcXdusf8OVbyPAV3ZYtxgwcyVEWzTuOR1YeDZRmo72f8CaMobNNKHTKC5RJvcj6yDE6i9
0EqKoR2weN425H8xKsL8QWuEOBtxBPd8vbjzRjnNlcblOZelP6P3mHExFgP3Ui7wiWGha3mxK+oc
HcpEXVfzOvyp7FMxcf0vQ9FcqWfEGLx2XPKLshIPBhjZDf5ppIjDuAglibYDVBVuSdlpKxWr3LOC
l/4PYx7MV3/svERddRIn6ULhzmhISR9KKzzLV1aDrETNW0zx/VpzTHJn9m0uk4SliPd3kczU0cQZ
Di/GYLwmyhXxMZCAmCGrvOcxr2jFBLUaZiaVkyRnpTqJ0b0LWhbAdRu+ghjRRfdiPMSmq9BtHhyK
VbVGzL1tq9XcagfZLbhpEP2ir3CDpJ1aqGcO2fodyecMjoeJ/ZKN0t9t9nLDYZJK+cr+uCRKk7tv
NKgc1mvTKe2jpQ0KazQhqWcXba5PEExewSiwV/soI1zRo0N8/5tQ2ZgtRrClShqBhchnOJBsy6W4
Gj0DjcZAUYapXbY7R/DpxvZp17bZ15RsvY30kUtj0yNva7kROcY5ZuNic2Rjkqcgum3OQwdQTgxE
it/2Z9k9rDkOVNinDwZiPYPCAuMNo8OZvx7bMeoVj0wacLN6huYitIUcfEDg0s/0LT5VKtKmlKOk
X8Di8WM7VnJIKxQteSIR8z/QoHQlzzRqiQdSgTAjv4nVkUw7KccuuhE4XKpcUOb/r3P6ljG1kIZy
4W9JNninnOsXi2QRuc+2MjhTSlxhH29/O0OkuEzZZGcTsOfSSr1Zk9LvzJEvbRLTaJG2OSx/RXZg
x72M6DPWz8i/mKPEpHfzZs4lmNDSlc6UXgm9Up244z9J4DD0qZJsoHDwNpO1sut1FhsBncW5WYZX
uV6ndqvkEIkQLIew35nM629Yg/PJVV9MR00EY75BQ2UeBnYj6lmtWOD6/yRYcpFxN8Cs1G/TrLFb
ag7q3HNllXtoZFMhsH/TL+cQpaesHlOrEoMcE+zQT3ZSmsJNyyx6WorNInyI+GO1csHn6L7tdh72
GCak80uCu2h+i37dJQM7qvchME2Ju8ZSuqIKXTW5nAHHvtDBLQlQejLkaOANr4lv81WcZ7TonNYt
kb3d1uKAKBoKBeTlBId25SYv5QDw8jEOufSLPKlNCJfPa2dckEJNG4nhlHr3SeFVo7OHSnvTt1zM
q5K/ylqz/+xrxK1bCnWqvtx8JgkS78DA0w18IxPImk3YaWJZNORi124lIaaf3ci9ifvuhB9y/SFy
jFMBpyC3Rwch+H0fQEn8Afmme4ax2fkAnHrTaVno1ZukF9hKVUFO1OPyvhyNOeoVPGfXTKVu4PxX
uZv0gpwkufE5IMnDVAiv05a/SdZO/JwWOhMzjfPusuAzAJbcu2E54/MaZQab7uN5iuCise297IoC
NDyBMvSo5Ya7FMcdLkeyHm9YM2s9QwmcNzuBBlXhnjLZL8XLMF7ooZWOJcYTSyXkIDs4Aei9CPvs
91d5dZBaUvtKcKIfFczyyyy+ImUn03d3oLhJcOR5+gJcIypC/y8QqcjB27gVGUp2y4Bhxn09bjHw
k+FlwHg/GzZYv+pv65Swn+9V1wDxrUuYy/LrccReZZMCdW7jeYGDuQyk3jt+TU89BmvB0O0si0vU
0mnJmb+ZBtTu+yvIBS0LtdVOJqlOXWwtvtOUKSKj7UnSDBU3PgC1XslmX0G6rGvSb0sWIXfkPqKO
3xJoaAMrfbyXWv/z+s1vrNbA90y4ceWq0Z4QwdFLFIXy473cu92zWB2/8+OhdJE5wCwW+BPKZRcr
iYpfilLXPaJq30OgDBUXWNi8FMbuci9m9xpBrCjgB4sFwQn2MPGAxBgOr/RU+dVAMzN0JcdEiLxs
WWiyceie1K4UcGlU/MeeFg5UW4qv+EpgchVM3xsbYfK4Nt9UcN7I1TfMfJSMjyOTtvpi5x6tsyfC
QQEAp0FSVi2+mwO/zAOCCY0NJuJAYgzQ1ZAW4fpba2dTpdPdeuD70X/gtjkIJaIi2R4qXdHtbRMm
T3XwbZMbBB8/JaCzNsMFBzfDW2KL4sWDrPoVyCC1u67DFWwDCJ7KreGOmyLqHDnULs9OqsM+yUzS
eyqWKDYrs3LqzKdySNqBlK4tkVKVypoIVw1OzaXNEVL4CY2oPaj5bO3qDpOsuGnEe6UwJ9JudPa1
+hodT3h2+lQKW1ZWQlcwYLEPTceTL2exfwCHj2/DwDKiyOc/XL7YJPbqK2kunu20I47Q6IuCxUo2
pa4UeU6+ZuS/MIiQWg561Cc0+CMo0bOnKV6oZUh5ZzyOZAddu7es3IdSsUPJc6Kt4yOEnNtGoGEE
vejsD4qSOr/r0uyFmiAS4WaBGF7SNu/TPrVP7euyBKy3avE3cZACO3v/NIGQxsReGVVRb18X7cW3
52/XRgdVyQjSmerOp+ZgPwYXV+uN7X66qn4Ah17oWEUobQ0/yT6V9GtPBDv6gciNRAMFcWvzQCzb
UDRtF6M0ET9GtOhluYNk1wk9wEx5owmhUKs65talUz20a3fxxo3Kt2goUrJW8MQnE9d3SM2G4KU/
gh95V6foUnPsMyzsnv4dfjQT6+H8QNFncspAyLshbVjx6ofwBQbLhPvj6jZ7TxRKoheqzE2r7Iix
I8djSnFXLfYP6iO3EiJ/r9goDU7tr4vLz56EqD6pYZmI/7U3u8yCaBmB3PWK5mZhJ4f68BNOcUH+
tvgzdQwHtuGaql1OiKrcw3EEhisRUZoOlO7hL5EzAcvHSS6HJwrzavUeI1EnjMQP9KDBNt8RjcB8
+97LxuKZA08nTzD7ftzXtupb9sIgJ3T4nwMiBKzxeuNb6Hjrbe8M7bA8hedNZIkNkek4E8nfw/Ze
Y1becexCgpDQ0+glPF2qT1uH6f8tQaj3oPg2vs/BzKA2lDR5+Smufz9oPTPfUVPR4Y0ee9TiLjdT
DdyZh9hB0vC3HBcQ6sC4p+SxeGxHRcbLjP+TMJ8wVEZ1wOhDkl6qonC7XomTY3+hBOOYxv1nS4Ur
SIjFgcMa9UCZfZVcZ1vDyNDyRHmAS7WIc6JjLbb57uvDBndtAY1Y4aPeF3Qa1WI/tulJtvG2+oKr
jVhSJozwfj2XDpFWl5WSIJq+uHMmgbpU/3sUYkyi9OFTikd2o4se1eC5qMZHBhALdS1nCs9mEYFv
lyNVw+JBLfL32BAVNvjX+2/BxKcouoGGjGOz8LycXyICbxGsj2W9rZGEqZkWdUqfQ8fm/pMdU+j3
LeApmxY1wT+TUJ/HYlhLPyL9RgvX6Vdgxv5pAmXkhsOw7GcyBRvrJm5Yr36m1Jae862Q6eAC3DYl
fursmMA1eCQ02I7X8lzmr+3h7MjrqYgb5xoTwqHoDiFDKGzzjHvQ1LwYUXqs4C9pitI49cui/z1o
JJZXv+rsbunr1thY5Uqqo7OdXRABW85Xd0bFwGGqMrwDopychKl+/3heqP9rSVdpAiBmx178fl2U
yyaarpP2kHqxARNAXxF807myKz7zb51eQqNs08L8GP0NuNI5lIqAIeNdTz+l3tmVs+08ScswJOqq
St1ow9OzC7TO1iXJiBXoBAsty64ZgYKSo5ojNWdSmDBRiVSb1Zqyf2guN97K4ktBg93fAYUjAp/1
thU3a0TzRu+lWH2kggsvTTmhexLXFYIqTsKcdXz2URuAb0yfnWya83kngEvXZek2/5sgWNQwQMVB
e9P/MD38JZZHhO/EkAKRsIpBxwY3nqql/z5/dk/PxdfIA81Tj9bT0HwUcURslhBLV2U+j7ayZjHn
eTKm5WRmKWoL95OAS7IE7VASpDT13mj3nhquBQstYGHt+UqQwCBsdGMMs0IfV3wT1anx7RvFtubg
tbV5NfSSMkvT9Sd9f/tZALQ3xyj7ofbBPkoSsXb7N0gny/NDyzwIxJMZUQPjgDUJcjfbBvLPfrPa
TIafKadjhfLF/L199fOHq3QdbflTJ9/EsXBsD9BJMZLxdQ+pcY/zuFciafJjGRjPC+2/KA6q6jlz
QF/PW8sONkBq9GgAqhhs/8GUINsCepWBJVU2jJXhdk3PRLGiHyuNwXk7llDrHEToB/hXRDJ+q1/A
GCg9Nv5uPIdD0thckdJgjZes79o8wwv8ura3/Fa7zGiAQ4F7/4PPcKgDyMasIzPzRH0CE6//xogy
5umemPDHea1l/Er59H8XyJhEXo7XhI8ejJu3d64VMsOckgTOvTzw+xQwCj3q5fFDSCxVdIBS7PlO
STlGNmKsi7lp20DSA4piMUftYbL9DiRDnu1Uf+5eOq8gCEqvp7vP2atuUExQLsyXfsHN6hJIcAHd
KvcMYQMBUiXfBQxXvbFT6MtKvOzvkOccYmcKIR1AAqarOuKsKRkuwtWq2yBa1ctTMo/PkCgat6UL
P/9pQTZzwBTKxptdVJjlkGL9BMhZWfjaBIU3VLWSoW+eoZli71cI40FGKfh1XH7IuqPyTS5P4UoN
ZfKGnwaPjeouJRT6rAB0jiTHS4wgbkFyOtZOmBOJD40qgjAs1r1WVY7QlBTvd8qlvu6sIzsL8/XE
VlSZI2xOow9iH1avyj6EWgVFiVgDcvCT8nxo/VBBVi3ZOpdRaGevAheQF4JCj2xRHbq5pu4+guDF
jiw2mXV4wmpjDwKJLeni4WELRgsd3ZCu+FEuhMPZMgRM/nEo8fS77Qq/LtyjK9apAw4JDY6LyAin
z7+IbZiJWRlSxC4fK2qtUdBi4Whd8g7lim0whoNyHO1FrDUn+uMXZAwibJh/EWly62HSavTz8Ck+
ET/WU2oDD3IPDf4+0eu6eiznpsKjm6fmfUx8nPN2xZeVaAjdp0ShtESCzB7gzj7iyelN+pOHgKDC
Rmeh/dNI4o5yA2ER87OEczyAzuBucsnzr56nBJClMvMcmHZdoPAEAt4zsbH4FPREEAQkSM6bTg+Y
G47g5iCUHoFdwglGvd1mjPcODrX3MQJqzEr0afq1ST5IAqNm3fl2v0+jxZP0uU9mMdvKLm0J6sKb
79MKm0IpxIgenYTfamBw8pRQVnzYRQ9aP9kcuKXvrTAvHue6kCTZyBJMYZlS29p25bZeODDTzTaD
YONF057iDisGeJ5zYHvow8Fzyrgg/PCGnpWuxhqS79LJ80c9FwEoJHtVWHA7bbzClvLFpPqCSVYu
sFgKmIfQ+qEh18x7HhYculC/tpE5Y/YGr1aVfnJycW7kAEzyU3MJF1XwX6wYxsAf+4W+2PH0CEZD
pka5qzmM91ATqb2N0C0gwwNJbmtQ9kHyAnOlR7caHZEdde0yU9bKUILPCPmxsMynpq2MtPa0aO3p
zml6iF11+hng/D/7StVBYF1+Jss7fQfEaxTzeUq7+KwQ2Fu5alpRJS9auV4yB6onYPtRa7K/1/EM
3hqjbVlhmEzKjgh69E9UbqHuMtZhsVekcPqlP+vl0yYHX3dOb2PcFMNTX/XCRxAcDVym16O1xFYP
fzmB7NJCscrJcpWSbSkWkvD1y0Bo5vAXcqU4KqG0YLWrcJ0tiaBsxwBH3xB3JohlacABgEeqTjPK
VKZPSPaPpQ45jFjgnHUoGSYSeNcTqnwMPtjcJV66hr7YxCiNjSxNgv1wPF4QB/TMjtvW9qQkv2jz
XQX2ansCqV6SYhsO+TVo17vYBAxA7ZSlgkgoTOY6ffiKg97TGDKAg0fc4L0wYoOr83DO37RsyC7v
ILgwFeNUZhb2eNgBP5eFXhTusDu8WBrl1c+LSty0D+arg30aBt2n3L1EF3dNCDG6ArOddcxqrYQ+
NIld02hNLi3xQEEUXqxuuow/EFJ15F6dXHRNUK9WJuAa2CdNpveYFOqJG6cV1ZiuoGLdrO+Fq7Uf
n4oq1BtGif29/d5/TjNip9QkECTuKdzMxhQkICQ3OzLY3A+U1EcKDb3ugPqADZLttSgphGhULqBS
5o0e/qjFahoV6lg5mAfQGRIfNYX30XxCA+l+TEe9jme2dkd11J5Lt6lFsjzw3TSWjoiAgU6dtgsP
PCDGhOkPPGHJKPk8M4axnj6A62Pb0ZrkekxcCbXf39hE+cjPoo++0rwZCkWNUmyIr8fGyOVmMg4U
AFyaibwg1OuffNcvkdRrSxMwfSA63P0G9w8OIptu+wODSZ6sp1JbayCz/C+1DWNv7Sg2AwojKdNQ
3n4l+SjQEwqLrXcfzvefGn6sOH0CVlodzCw3qpagk+EJM+ff/Yq9aMAVGecZYnm92A/WzSpgqc1U
Chci/bNTjseBZmKG1JPIhG4ffpNpRTz4DcUJnYbwY8sWEzXkQTnS0e9oVrdB7qgzi4pzzxKf5q0P
Ga3ptjmjCcyxMynYM7ktWY5MccmN5BySQs4zpcFl8ypCVuxvxCiDbTVEb+azd+I8F7vSsZiCmOjR
Cx0rnUCa0WeGI4DrCh0Bas+YTKTsGKkY9c8mT1NvB8Ft++jVQUGsneoG0nL6pgYUlzFhdsnC0xrs
0JCRs/cDo6/RUq2RUJ4ezsMnHz5ZIrs3QSElf4+WOLlvpCScS8maph6knhKU0iFbO0TAUL8+5X++
LLBJDmwSlTaroY1nzMX9mc1FaYxSOYfrUrmLjKqTpBxvSrbqIeOOvlP2YHOTsiMXWO5IkgxpZ/qT
/S2mAxNW3gHfH2Hg5PZTI4ZQ+xl8nuTe6qLCeFyoJzqZgAZcIHzXCWIKHb/budaQ27ovMXzArObx
NzaGX8DY5/5sgP2x9c3HZ0gjdrZV9VbH7WyxO4JOiPITsXwZwzKq9SexoRTCM5+aU+h1isihb/u7
NOibWVlpDuBZqWer9nLmYL/k3jfbocwpQE0uqaXox/WRdk03Ob1EgI2M2HQ62fNmGwruipEOayTP
yH8j2XYMZ5gxd6f7TVdgdXMT96LlF+gyQUa8FBwR6hDIa8meZ8cEzdM4+CuBlpdC1oHJ4ta+pINq
y8rR0V8eBFB0naD0VHQURUhx8yoeZUEHVuHaAi5jGwYnj+PCBiornzbr1cx250p49Q/l/GFVAgT6
o7YFuLcWK+kkkkOL0r6vegugseprTrhnu7H/YZeUcxtakrgOJolg37e7/NJtTM6z2nDUFGWqt3y2
2GykC5WowuyMBigVmCMB45XJa/dM3K75/t96yd5JRNz1jnlroXycKw/NZxQoyDUbz1WOzE7jlx8E
TzAoCmQBFihBvfdnlq4y1DDyCnwxvk4WUkG5I9u+Br+AGA0YwtZGaBpP+xKNKTGW1i9Yw1tl0ObL
u1vPsFwaKhDdNKRIWeTCSwOr+33BMN7bDyL0JhY/sPsAiA5u+N/WfWoTwgb8HdBOKBpm0IpnLtOy
eFUdR0vil6j3Mk8eHPdNYdKtY80oeVD2bqcNa6uSNZsbZKtxG5hud14m9mhOdPhwwLYz8iQUREFd
IRNiSiNg6yYsxcVCED2xtlKRh5Gh/Vkr5UdV2Lb/sHpjdNBwkcBjhdtsyIt/0KHPSv51n10D91tb
EqEaUyQzhCzznVtPqoKOHxDLcBbQeLWQEaAh02EtOj91PesX/XzD8TcJbd8s3FHXicU4fGVN1ErO
0GPGj91+tZUEH3iMsmsth2rFqS+ifgKcRiQVUyLkhBiU1woLvZ+3wx7Y30WzmQiDAlokSAq2iSb4
E4X/tpwoeL2UUFGi3eS2KK6LT/YFv4043fdyEDsRcxwEUwusd4Am/DjO8y+LoOIPcTC5oric6ASg
rmxkhV2z0UwtRB+HLOXtqYUQ6EjZQZlCn5BJ7ktM15dUBBcGgxwuuOj+7qzW4zaS3owjMl7Nxcxj
LrlxGNaQZuRWFQkPf5FK1QlrQqU3rgKq+WHojBSI8LO83a4LlVJ3EJibph1tiF7sjNfYFqOSuV9U
qHMQ5lxFV46nQMYDBHa14AC04wIrR2BigDtQgx92gF6uG/aMd4a3ab/L2yzvBMyZlvYvX9K+jkLk
1toy739I9lFmwYNAq6vgIeO2f01b93qwGCRh3UUhwnyCsfpyVBcm5u9qDBVHbsTg4WKcrRhrsnCF
PQm9OrriQUnrPvwxFeLJwznyAXN21xmcwsewl0e4Y665I6FKkn9/fmD54lPkxDjYrp/OylwKOSrE
36q1zK0ExhujmZ7muSTUmolz6vBsnQffMpPBQOmx2u1vcqSorg0kgoFGrMhCv0uGE7B1sBQjmShD
LIzIraLlYc3XI7Xy0M6tT8uVlf3O1rApgXI6K6SwTzzR0Em6fBSBuGPJ+hlmpApNf8kg/ysx+Isg
sPDlBrE/jpISooph8J3AAGrFqauJgT+A3CtvzKpoI8keIWekhW94Qj4c/oBkILWn3b6kz+J9CIfc
j555mkaj2F3AzWacWWS0ZPKuqmybMsRaL5gnXI6XyKU6qxckaQso48ddFjMUXmJlg1tUDLjxJdtx
ndR/gc+G1oJ6Ml7t0pMRvO7ArNzheGHsQ+gXUV4RMjBK5uiEoY2gzWM7zwBV+w/z6xbT617jvef9
tFxfv9dBKHFsk3eUrOd30qlLzp2TjmQxOje6pPsByQVhGCQD988d0N+8ZE8Pdgp+CNYsrTacuXpW
VYfchEKUCZ2YrVygTijCfKKboOcUhKy9FkwVqUXtvyboknl7shBpcOz1fprMFn6xU1DfooxwjkFP
BhQXy3OJ4dsm2RKJRpYJdruE0iqZ1FGU1ivJf/kJCFk8cjcnwhdlQSN0s22mbe/XKEsIPEfgRU1x
AdoO5cpZsUt1w+21SabMksGJ3LVz3XKb9ysU8Qs+Z6k4a36TAB9F31S6vkRfKl0RN7lgGXT17TCX
Hg2sj2qdTcBbYLo0ZZ5P/sgR9CPtUcdTeqK746NFIErhanhmUcq5wUBbSla5bj/A+sFkktFYuvty
YDWQr02dwmYljfAHhEPbJT9dyC2UVBWvN9AySNYpYLs9GFnkU4ydw/opRXOB6pwnkpaFzikpen5k
M9MGRxkrpUDtz8RWFFBhQYyJJf/r1S/m9db4pzBaUID5avtIpR4DYIhrkhK+H1m4wyovYltOcdM4
SVoBAKiONpcABv8AN1Rkg7y4mhmYwP1eQD50J5AonRa65S09mYwU59jAH6KqqHDeAopPBDUkYGna
jXnElMvi5IS4oyquwZQmHaw3IsBRpFRhBkVeyLS3cYBXE+tArBDTKQWYvcuy6eZabEibtGP8i1T+
xyEcxOcq89Vs9dfVER78JH3U1z9YVWvKypkzyXBdtfNMlk0RgT2s45hvfw6OMSCLJb/i8QaR6bDQ
HgHGRbSG94qaCJgQLAJjOyiHSR7QNJ+AtkqFw1+WAYqCPylth50jcZfZuXm/TFM/KYlXHM4gdKmx
JFyWWBiCuFhsU+qgrYx4VUo2XPizH0UNRvxZjQB6qgkyQ5xbvzvD4W4CNJq7hiEwBiGjWTBJnq2T
GNI3vJ8Urw4AzTMrFFCjADD8IPQHIQ/XY/C/kam2CJZqt7g1Z4ksHn9vQz0U6oc3C91EvyJXxqZ4
mS5eUK7pojdT468wBYy/bTXNX0NZ82a18b7AnPqYmGzxkG8lMzgJt1s9ZRl7gsFto3cTXifvABhl
gW2fNe+EgRNmg1O9xV3aIiQOKDoEK5AXKG9TdBYjmxIrgw/1lQe/5TZXmpNFnZ8KY1SZ8xQ6ez3A
rhP57qHPvYrw1O9APZiguiLWSfjKX+WA2QTlbfzRKGJBsLfARNYJyrLupN29Oce9Kwg0LVVUGTes
VQBJESkZ2fdXpPMf716ILciH0/F2USU2unR2LUdooXYgu/m17vt7/F5yD2N0l3naSS5y4ALm9AJL
A4to9fRS4OqwT6QBnqS02mLnowGVxDfJgRJiqIXYyz7p/HJXInt6ZMCvV4Hev+WyoS9Zj/giQ9Nr
l52+8d9QlUW0sM5WOZouk7mKKX8yROAyiFzurRo+wFM8bz5GIne4Ph6uXOyu7jWu4VO7j1x7mkwR
pZD+ur1e+g8AjGeho5mmTP3HYyNlHwennVCo8wvHycYwenYXASsecHNrrtXOfvXLhYqI4T4M10F0
tZGMo15R1BwDPadaFP1FwRKpeixONHW7/HvblXdR/cqRVbWup3rX1Y/HMat3fQvGVRToypQqmQP7
mGQ+HSyxn0pzPPTjynahJfOvTJB4z4vJd4Act/2fAu63RR6VO1DuxqZqeOZVOLckbFIxHJ/nDefK
fyLhlnXYBwwTEGquWMEm4U+fQicBuepa3qcAmaUzB7UuljgYKFetWJW2Wwbs3on/TRQCZ0ORlndf
fLgV42F0RYbeKwtpF+LqYrd68EbqiLHP+MLI/TZLs4QioRUVGRdSUpmdxzeZiRiPFXCvM5d0TsT1
VCkTF2JD1OW1/s4lTA/i0KVfsbnOnNVOvRd0+llt3NlN9LNd4XTtnTqJyR6TNYjX29pw3uM35Ztu
q+bVVzYVj6XuEOqBkPpP3ESaF0y1yukxWneQPhn8C5GMj/3t/fCZccSw9iYBQl1gRIIgig1yXk+a
lhYyq8B/LVd5qj1L0rtKEKIMS2L8RJDhlAWyAnPNqul4/vF6/Nt067exhh6LCoDnesUfrdQkfAin
203kgm7EI5E0B5/RSS7OBK41DA4NyIFJww9fNRTy8MAe2USXnim5YdkYfhEpOKmVboY1mDA8636i
UYe6+p0CC+7m93cN5pm72ljGmQzHZxW5UVMrxnzQMAx75GuRZGP9poMZL7Pvv6u7fnKEAXttPaRb
O7cjHvWo75qqJNY/Ts7Hxiu7qBKniBgKA5ywF1OQP6TllMonF6zDUgTpNR0QuTvklrgUjJNsBsZ4
GpVLohFXIYA+SchkMAhPPWwqG93QQOdruCPMqKmeQQGEyL2JFz9BJUzSozGlMmfSoGQL+UcMF1MS
tnIbSHVmOeLlOmsYr5aBVgFwXpNpWGoKCNsPnuDTrpTY3lnZ7obk8EVZlXwju5JpcGgTW3WQjd6B
FP1EgVe/Oq76s5vw2YLjBScQfHREB9OrSbRo1dBOlW+D+pmdOG0WrxQ4d8ysoulM4cUTkQUARGfn
iyfQ3Y1XRwFuYFzgf9gKIzkaepkfXj1egScWSI3k2hWgv7U7NlMXPTPnc89xB9k+0GZfiiBPY7/8
H1ZuIfJDSBQx5Y2MbnPmmSqRIuWSYWOdFR9lhGQiJukfot6HyTrYruk5JJZOITRKvO2id74uBa59
Z2t3aHn9idUP756GegeYITy6bu0wlMf7UOdW/Hl4c9jK38B4A4GRPlDsoDHA06c6uwN6c48VD6Zr
x9ldfjm+OYLH3fX6WV6jRela/eoI+v9XZ032E2aZ646QdtnJvX9p2BGuYln8Qj8JQnO4eJTFUDBc
3EQoP3ZkT+a6zn8gHBXezi9DVNklTr2P1i/LtppwrXRK35PZtSN2PssVFrPINXPkLBYSUlKziak6
UvkUuKeIsAk00a42661DIh8Fa/TiCMK4hQSWlrzVzXeIjG4JmoXQ9uFiM3k8GCo4w5yBs4lMdvnL
yO0Wk87IdxrLjKZQ6Fa5woftgWXi3n+0C0TEyVoVisIc3Fo4BHGsytrzvTxe66OtS5UmbtdhOVO7
cdYMtrRS4dRpCwUA7WLFWhouPVeXNjNo/cRKVjWjnJGF5XbaI4brrEBcagKl7yyzlR73zqmuvIWE
vJtg9euo1L4ymRIfFOSS4jSYFBcCh2vdK5zInHje3Z/b57b8lc1zHAN0uilf6veBBtxHtVxnpUet
sAK6i5fvtw3sSt2fPfYaNwiJxOFZeAR3Lhq7hjTZ8BdLw79QTqlHlJZN9a/lJPmqkwtY1paGqiGp
nY5587IdW9dRmubjhW8UxREK8zvvblcRA5wy2jW9SZDRRo85U+np4qqZaJu9UQyK6ovdS5fXcy67
wOw6+l6t7DsnYxKlwvRGCSo9Ph3ryw6zF46+ibnUT5syfsVLOvK897B1KpqDT+8b79w+5zNJ7Pia
NjOY9GwFljcRzwW608RpibsOilHOVa3L1IrdT/dL2JMnkpeJcFEHsu+etiKcCYTkmnDYIz2Mpre9
OqKJOBkUblrDSlNiIXRNShCJG6dw+SYZIo+w9n2r9VSWQmAdzPxLZjWuqbgTthlgVLlAT+JJXeCS
GePImuOyW8FBFmyhqTv8iKnamsOsu6ycwlNdadGXbGCDM+++LxNIHM1weH1ai0zD4FIFYdzK4WBB
potwT4CNHnXjWKxovhy7Ktr3ilKvxP+FKwdqBKttWi/fYU9GHqi+z5gbYDwctdmkkyctik2/a3zr
cO9onoGWPUmDImd6bU6bvHSHUTvP35+H3K4fmY9sc/5QSCCvfI0+FK0MTLk6PjRaMTign9dw18yD
Ciu0X3yDUESy/JoIO0DCgVdriJR83lmbqTUh6ANVROrfBj4w3nQwsZ82Wmbb5wEXxLGKEaoNvmK2
FLVvifvNl86GT0Wcs1kNLHFZeZRiJYUaD+ZK5+Jtqy+FP707wRRN2Jno0DooDvG5KkAGmsywUdQx
DTg/LhnF/ta9bz6bCR7KwK2JioGucpcI5A0VfVsRr+1yFR2n+hUDRLUkddt7b3td3+8TkpaTeH/1
ySqaNn27O7yTvFo6tRdG1Ij2kfzZrTVvFQ2qJ05hTB9APTHrHhhbdoSq5SmbnNEBT+n740EWDc85
FntQM34WdQZprbdtEPxYUu4VczUkbOUYsKgdXAF1xJBSNKaeDxg8cDUlZ61hPOJWc6Ya8JynaUoH
RxcGO7+Old3RLsQGLmpfeW5As38pm8HNuhsmZh66Fsk0Es+I0lL9dMzC0p1SDaK8NY0JK9MElD88
NBpNAgg/NN7UbUUdpCjL7RmizbHYsrAWUx0UyrgwtmRX4RFC8Iyxm10/JrfdOiK1kmL12Y3MBvxD
wdHffrvpYcXoofSDy9c0c/H8FW+Swmo2Gt743CKMirwQdpaGgUHwusPC7jhOxUWRC7ia/Hp/p3oL
cq2FxrXuD5mWMyilxDeReA9DuiyTOZ4WeKuUpJIsJhXUiWE/cZwXeyd7lsZ5nPmKYZ3UFRbCqXBW
JFXCVKyQczsaW6yTgzN1U1nYVWIMBHF9Lrk2hPvGa9z25O4yfdXe/T3I5ZzdCX1GCQT6haLWZfl3
OqVJjsiLFq9B2Yqy14yO8o8NFhTdv01RqzQ8s+Vs+Uou37iFGoMfXxBDLb23fOyF3mENebpMtwQI
wLejJQ8F7PoJPNdJFHIq14+oPjLf29XDb38ThOJd5krveuKsPpt5vq7ncJ6xGtmF8YkjWNIwBfej
1+fpOAYm+A3jJuybIZquabRJ6ZQNNu97TFTRaTymDewnzizx1vJuqUzbQG8A/4rTKLQo5r2N2+nQ
4MAb5CRG/cykprlilXEjNtdq1NuRyo0UPXS+j231JfSj+6nkVEUlgRKahB9DCVVynGmM+KOHHdto
PIDmMCbrQsuJoXWKIsN5lSHIwk0TQtSmmlZw3ZkrXH/U0cjwE4532rATCRUL/bYQfwuLHIcJNEKl
n9LnyH+uqQJbiqAKnGd0tkL+97wxijEhB4evMy1X+yx9tjRg63l/D6ScCBIk2oprco5khcR7tFOF
kbKfBsLLHRPwmoDrhIRyQXYywFo2PQO1F+sCKiBlRrcmbr2URJAVVrBTNu9aLGvlddLF2geiFqf9
pf1wUsf/K07rIO1TWh0bKZ0uHAZ/p2X/uUcRV8K4F2cLaMIK1oDakheaDu2W9izvSdgQqgNKrnbh
XCC/afBiSLl3YVbbJa80z32kQmbrYNei8sY/ZxlgqPqz1p6+1LcpeK3P8W39qfLD2Xf7mEAxSuhX
xz1OwGoHKbEDtxb8/MMfOWjLhhaySL3RxKTOI62B2RTdx/gXwN9MwD8MQvuftfwVtKUZ59F7U7SK
P34t0PoezvYj13fnPvsi0tr52LVqwQsdezdbNc0Ahqc+qDoge7B/BLYG9wwsVW9lrCFiCIuyMheZ
lU6YgfLw+boYn29cOFyDyorGVdx9F/TsAIDmSMddeRUM+qKZpBakpV+jE6MKBRV7oUkaKAJAM415
y9jMEemOodtDyVXPZGuZSv5MvkDquxdcd/K1cUwu281VpcPxDhF3fJnyj0HQpSy2aWBZ6rc3+qeW
oxo3NO38JI1MV7cRCUBK9AcWywMtpUWKV23OGIyOQcscrk30S0LFASCNKHTaC7VK+qjOZZlpLwRr
pgcTsj/RP2nxGeCvWwCpi7P8ECz7KIAHtpCcjzWDvUBsGW9rTGqolXmcFn8BlhY1MMcnRvrlgVpJ
JeaKfxIhleYthiT4YEg36FVfyb32eVyDzKmDyHa1FxQA/sj4ObL7U3VsLt4zZT876KXcVExre1SF
bb3u0YAla98xZ3fci5597PciWcXQjSH2SOCyTQKw5ifp/sdQ4dFDZGhV6O9COFJmd7gnv5wmSf/P
50ZFHWWNET5CDhsbUKXsWjOjanQaAXgMFNBM2KH5CO5NWRgeOcxPnJ9F3nzGAzpl1rLJKPmsTJQL
xE5P4EZ8PyGWIg+XW8hGVGFdJ5R0+CFot619f6I+ICh9pBb6FgTUoeBAwFC0uK63UGhtIF37PoiL
kYle1aIw09P4rGXzu/HBkXUvMmWS5JpzQhzCHYkVeltboEwAEp12h0lkkdH7KichkRArSOcZrteF
SNEt+ri3grbYWNrbWPkm04LPJVBbEkUekPrRdBu9+gpuYJAuUmWEBPGsf3qPecXXFYZYjRLYQWet
moYi57TwEMx609Hd0M2BZvBlI4ted2d/qUORe7Ltg49UNYNU5+PPXHj2M68JHLbMVdbTXIsXDl2Y
sb5GwvTDVeHWcZc2b00U01hRSmMfaMeeNZtsFj9vyuIeS/3IoV61s0os35uaKcYTH0b8Ejp+9bjr
+qaEOHizubw1AJR8Uxi7ppeqnBBTQrLriaplLQl9ZKig0Ui4R4VI7B+PUXaEdJBH4uKkMtBlq5f7
5ZzMVeQAUtixLDsfS6QsyNnBlEYCbcUSGnwsTCXbeUcv28ZAZOOedlnQEQYYADHNhploU4guPL/v
bpyqh2FIUl+N6ZzCZXQPxuIDzdRvScdFNU8O/5quY6vKYIBOAu6VX0g579ar4hAXDvMZAO6l7Aqf
zmmv+8eNgYQbAywdMx8FWasXDdZ0Tuy1EaSh23bxAWe1IaHdkeOxMmLvyGKEdp56YkpbJrD03BFS
ZK8PBV01MY/I6vf+63VGpI+20n8EFiPo1mSLouUr6HGxuYRrsqvpi/69FA2RpiYr/umrFqMPaO84
yx6LxIj6tySDfC82Wv+ONRwbTbZ612hZv9X5DtG7B00Z4cfLO5MHhmj0dX3h6zpOqL2dL2ZstPfS
Tbw6BhFcpOS1noPYSNVGn69ZyHNOSk2O2G8Gzsiv1YJIb1Q21/PWD+ysjGo01Apyy9HoxYY60qwn
CxHTs8A785mLFVu1k+W6odJ0fc22WUoMRqzj9tZB9oMyy7taSteKKyrae1Gu/wrd8CV+XCDZZjDA
625AL9uXor5OtI8bi2nP6iaNwG5uumbGXV6lvUsIwa5rTfMFU7k9sXsv5fpsOdgnp05pSRO4Tk38
l7ovz3Q+M0op2L7VRWvUYWgODv9fOgSz0Uu/ocwQwtqGdFFFgXJXaVjDpydIr6u50VymQnDwrmZ5
nf0NYWoFRVBdN3KVeU03fyXosdKKzb4QBMr6QtHCZzQ3LmYzRWTSidlEbwLHunXeZUgKomOY2QkB
OHKw2GQe80eEEsL4JQs17hBRQaUr6KHyoDhYjrk7Z7ue3U5LHY5L2cWBQNZ163n2NRnYjQ4sF8ud
jAx2RSTRtLJEmIzKC0GkFoS6FxbhjUR4nhVgZ7AI0iVIsb+UBKsfZYhZDWVsjPLpd8xqTcJbxlOr
gKx2r4TzS43dK27RR5Ju3CtE7OrU48xu76fj1BT1uViZFDbxrzcPUTdlUxantetwNNrwr601FsdY
UwtoaCkmHX8YYp69ffAtlAlUYPxE3RVOkYs1stLjed6qlfyEr3hHV13QUkXNlYqCLC4b2rkiAhCu
PbAFcratc9oPgQO4zyOgouzl9FBikUJYuAksx4NBx92bsk6VUQ8rKtgpos5gIOEvYVIbzpcYrfvX
3dfOMLJ9MM8yAICwPBhyPlslJKF/6pu5RoTDENqZ+VgbshnvU3cqnkBoylXB4abCyK551QbyWAxT
YIEaccVmXTOdclpXTQl0+Z5WLi2lI4iriYJ9GmiZTxn8hCqZjbDE/604S9NaA2nd0LzCFJf2FZD5
vNQGY6oks1fbe+kPENPP4fPo8blRZlDspYB5MO2eI3nAo7UhzRAC77byzoGOsgCmU4T64nmcBmG1
l+tmUlJ/bnd4xpDVQ1kcTFSQ5jDAz+XI2uiIJLuwcO9ploVJzeOcubSq3yjCI87y1mOnaC3O9a7M
XtpcowDcGE92nTjnxjCrD/WJJXOX6lyth7TrH1UliAfOWYywk76Xuoh4FjIf8JrOnevWG4F5DM6a
5kbzf5V4/ub7Hl0y79y948CS704IajFtponQ74HEwgjjwRP/ge/tHBadeNeP2zjooROG7LUtrSxR
VYarCivhXJWweRhGRiD9V0yXF6QJrirtPn+rG0ekgysW1jld3KK5siBiHphghQ9yTHd+p4YN5Rxa
da88cq9SG/pXRxueKQin+vh/81wzhL5Gegvqd/l1r/WYE9A4IOpxbzw0eG5n+tz6oStor3ddYgzR
07Nb1u8sjHcysh4sMR30n3mP7JQ4soePagMokBy57iIDLb8oI1kRFDxVq2r3MssmqGyzHl+s+qu1
plWOvvps6rOx+njnz15qK84sd4t5oXCXf886rqxfsXGPQW3s/sDWn+AUuwxwkL6yXsX4503hVcXt
y3qL69476gxUDjNVmuSzaEvKByjRrb1gWimhUOkW1+ERhO7m8WTDnWqDDzUc8s+peinnj6QOTGzS
HT5NcbhGkgVOGiCq2hP6Tzf+zbJ2KZ4GbYG40MSs2MB/WIubLTs+QmGXrHKj5v1oKPZuLV+GAWCk
wcptKhwo1eZ9U7Se2s9KUYe/IBZ4wn4tVJhaEd1DL94078FOSdqxvoNM4KhnKUk+Frf7e7ssyc8U
UqWCGaOsIWG+Q8fmWzPzlxzhi8kOq1AXV7cm5k4VPYVIVrVoWGjbZfV2YT5QP8pvOcIFLezbkwpv
5mLa03RWCUG4omPWQQDtvV9GLDm4fC19b4mJynK6WdN/iH3iwaIsPhCC3NT7Jbt7s6dUx/EnEbnK
yW9AM968zRf2PBvpP10cdaBR35gQpCAytu64mWzgDzQvFobKQPP2cSpB7Vh8baGUlF0DFGjR2Jf0
UGxo4dbvLpbbgOaruF1J8g35eCoIv8szhf8dgzCg3ym0EzxQFLBxu8M6ITfxa8T3ZLQm5WReh3of
+KuAGFRFNCO3qHUQYPvtfXToHUa+312VW3/B5ocUCl6yMNMwjYSwhLM5t6ua73m7T2GW3CNBuczw
UOIVvocE5bFnfDwmc1V/m9X5sZyWBPtinPdwl06V+a3msnN+Uio119HmfM57upar2jbXO6ezKH64
CjwuO/k4LL2cFwdaSVaQv9SIzhbCvsAqSLqWV+eq3Zwo4FjObHLZaaBzKdZT0hAAFloI7MnEEZtz
BvUCKoFY5z+7d3NYE90SJ6w7Q480yyuiCCJQj+FsHvlmMyO2f8NnypNKHQWxZqkSpzTKBDH6hSfU
hAvpOzm2YRnYBsgWCX3wfMcE51ZH25caKVNJbYfOo7SK2Jf09fhlUwZ+cnerQtusrhquXE3MKwt/
b7X4UvpgXc+tRUbGRmlz8yCt9YJ7v0KZNJQXw8MrvksklopNWif0tquIt2iTR5w1FvZ/VUSt8HzY
se+gV3F3ZhTBYpcmIE60Bkt4gKobwjW5/EHcpGKKOvgpl7H/NHwuTQkQP7D3rgg+fTyPToQy1DPl
o6KS32afRxxr+bwoJrxC7P0RVs1soZbKb5/wYkg6Hgj9s692eYcuLJjIGpcrAQTyCZQHEem7ZxI3
wVF6aet5rQ52DFqYpx8H7YqnrgXzNPHbBco819/Nt6saqLqoPilT4cw94fPz29bf82coiwYmFxRh
o3x36pn9Vt+5OCuyqWGvLBscdE3s6rcoBapvMvdp1FKrlY+o3hT6W9VCY3PjL/p21fZ3MGcoNOpD
jmWfi7jXY6QsdbYQ5ZxoAh/ZRiftoqy4J1eJjYoWq1SnEjuch0IDhCFglgUFOXBpRL++zlL7i5sZ
2cWL5afPtE6dQMAMjpsjajfPdqejRgIkK2cFusYFo3Gc/VhwQLSj/DhDQS2AqFlRramWsy5VuW32
+kHsQ0vn9sArH9z9vUD/9Ue9qLagU9p/gHWLoAe98qt6uz2GP0KETgpiisvW1VKiA3QxGP1fMNTO
dUNyj3SZ2/x0QowiVo+sm95dErSqfpXOLtH+37Ud+9s3yMDi1UWwOdxJIi/fAmb3LzQiM4U8gsRD
RAAnWiOQnDwkuyGIb3u7jWfY6GNyZQVeO2ywCzbmsHpRJsaDGAfP9LRpTjyLfvEcG207Z4vOWeGX
c1Tbgu1OOu1PbGmUZtlpsCqAjKOgMW7++oShmxULY17EtkacXOusvJXU6rea8XOKAzDviEQ/YglR
6DJGAJzpwLGukyVJ9UKYNylc5eI67fnCW9iDLkP1z1oo1NX1yi1ZRrcBkmRx5N092RSr9rDpm4NI
pi/Awf0OdfjqPSV/abh6R+iDlESu/yP3NM1iVL2iV9+NHK2MFKiCRh1ccMWbvSQ+di4mC0hRN1TF
57gTuUHfDoLiK18KXhVXKbOFNjZwRCpmBgsRWCEef0LNmzzcasZOPwTyURSTiCWmS42Wbe/ex0q2
GW/bDAVh+XQ/hTtIuRuYeGC44tBgniLpRrLf/SUpc9+ysdAkBEXPY6ZoTqR8giAj8FL84iIPUqKs
vR3tTEqBiYtc5RHafD3MEhtgcvyumUMiPGlenweLbSoTFwnY7lBKuheqNhGjd1yKQuAri1aKZtoT
UAaSiPBrQb6+5NO/ZZfptpUG1oFa5AiJ15hALq0psu9n4dPhzJDMdkTvSN13WCJr/eFLB1Z28N4I
hHoubzCrGy5YlNIoJXhjpZYF4LnQ8T4NT/FyuXIeyKBi4SMMsAr1exFXNGVBvDzRdLo9/QJFFqcT
35SXcSRgFqfOoRT5g8GAvUSY8CRJetLisXOk/OZ8XZZrKobMmYMzC6uoqs3JGBoJcGS+vZ7BnkX2
mJuFuGQ4z2GQ74BXTsNqKidCrWTF+ugU1emD0XqxathI8F0/OdZaMidqNGcQfjOoH3U3cfGbykv+
fewYbmqFl30/H/2n6r6Z7KfbLTlbQymDCJRKTmP8VbPD7pGgAtYnpeSEm15uWvWcPQYuKyplxudm
6viR6aTrKZUGOZ0A61akDzyIDO7IJynkkmlCmYchQlf4E9IlQqZJh/ZIjtnzTZ+nCEKYynxEswLQ
b23DZFwRun38Ev2Kl04u8SbJj/wZ5aNKwoiM8HR5+OEnoLToTddcrmGw52f6WcjgbWxvewAVqiw1
0H+hFQGEGPxFRAzgCi5RQIriY2hp5kAFYxrnPpdzWgxIzHK6DDi7ZR/MykacX24o4X8w8yl2OuF7
Hl81A681jwqtlwlOMB75DhkMviV7DWpvaZGYmxCzLYOStQxEEWzTVC8c4mSVB5uTJXOM4QF/RZ7T
3FIIDYrqJsY/D40Dvnyj5mQikQOB0KmbHdhjxw1Kw7Q5nE768D53nE9960zjWXoAulIj5ehRusRt
jivwwx+4gJ2S319ZMFa7osBac5qmcLHaRrMtlCRkypaMnxzydmFSaVk/DwJ7ybiZMMgL1JBSlkTN
kIwlz4YoQ3HJEI+hbDd8p6aRhuSlGJkfElwM3QpMStSqU4hp+a9rqXeLGpJIPnsqlDWSG4zDJEta
AaiRxeR6BU0mWzx9gw2t3fVB9pifxYGnmWT0Yck7Sxx7XaSANqj9SeUyuAU61K8nwghXRIAO+m4Z
7NMB8OMBN77/j02h2wyRQY8GNfbXDWjANE+9aT1oUpqvoe20lK7TNWI9jHEgY/mhP5Jr7JheBdIe
5twp0RqXf6zmLwthRUoFNuJfGHCZvgjc0t4qzHewN5i0N5Sc0wi19vyWNxwiafpWk2pcm2v+bEFs
PzmHbI1vxANmD2W7ni0YjF0pWwQ0QcttxKzopopT5UAwgcLZAz9UhzpIAZ8WjigiGLjg3qnlEP6a
3iEezD0Tz/Vo/rn0IpzSDCJTIEmqVQw1ZbmyGc1zHfAHndWINeHI9x498V1EUrFE+wC0EQDlzmqI
pIV5N5qWI8vMcaZVSCohhlXYC/katTGtLYKmRMI4Q9Li16oHr8jZ8LIQj34srRSfVc51tqQjnWk+
2d6xMBQHUmnrZ3cQazi8/1DPmqcPuV+g3WG0q/slTeXCKyp4Je+E7Kk3eupfNnatKR/zOLw85MYE
WVAEF8IUX5vG14LmnHMnZt0PiAhMWpUeyRbWb7APp54qnmYqNIsbRzP1+tGj3kX6r2carzovokjA
x7SGTDB8LK3IXOSnigNbSjwZaNErHkaSTdXZgCGnmFhlIw8Uce7y4jpVaSFOTIAgDl6i54upHBwq
tPtV+xt65GEdNWn5xlaYw0aSV1UzFUiicxc/KO0gojPW84mFScYTKiYV05iTIMk4mp/RUSp+VJuG
1gt9qmpYHL/TyUqJbz1Xuj8YKO1xYL2xURKAK52W1YyRYrqjTFufX6++9j95b8wTdNKmtax3xU4+
nrbcFaHpM/pg0msRQ+0zyKPgZCVN4ZnOWpLtEIXQpIXRNCnzSCtfEuTfgQja2Kip1JJWDqto5iEh
REehWDUiT+SOQIDyxOdd1Q4WFl4mlLbXhLp6H4+4aBHwYXAUN5+8IoDk3EiOiH6aq1HOZiYCfo49
Yuag6QKVBWuagD830L9ShcATNGNXa6BYlo3mVUVZc92qVmwQ9fVYrLxR3Dg8tvfxKFTcMaBzeHUT
cYR7m3WEqfk6fOC8O+gaWiRsyqwozMxN+Kgq2GkS1eNZla1LXt5zRMHyJWcjBwmFiXMtNhpfSp2P
9As0aZpkRvL6bdcQ0TaAZcuFJc976342iwgmagZ8Ho31unKuPiTrGzOYN6F/ppVhT9cLPNEE/z7N
t+inq35CfuSRUat/JU7KubCQ6wCgZZhJPJBlw7O4mQmRCnMYJQpUP0BwjvjQq+loKvoUs3uecF1u
xHoqs383W+rL5T4qHyEINNogvvkHJGSVOptMEBo/m+THG0pG+bV12Gv4IkyZs+Lk71EClmriGR0W
nqOpQF6288M9jgm5m0hfM3klTumh0sd8sFGhoSZhDNt2p6QJ71Pw22Sbw/useW6zpzrEEckzo2Dc
+uop3rU3uD6fNTJ9ktC1oUE5ESyQqZX/C3rWIumtcxisOyYBmCDsEb8TpmvOMdwoKY50JNFsQpAR
1S/v39WcJeVj6N0aYd7BKrMXTQWRgfkY+Gceb+3w6JYhxUBDLJFe/TB35SVbGGVbAhSZBl05uNmP
8N3GE57IQBM67zsgH9KrF1izERgDwxXEfh1HkDUL9+5ecg91dBlnU2MIS/xjzBYnrWU9Idh8JjDo
E0pxh7DZdeXVgsWnMbFZTzRPP3Xtc4GctGcfVV+o4j61H9xC3/lntJYw9AW9kXZQJx73xn9lrmRm
Em8BIY8NFGv4eGEYWa0IM38Mp14FtRGBQhASbZukb1StLPY6WLCwopaYK3kcYb/c7lQqUVD3zt3k
edNpgTYeR8su13gyASgUAXASVYYKpg7/ThklrqYmxGc6H3Vo+jMlv2nkt8lZIzwiGsNBdmkaEp6K
OgAqiuG1r1ablp14sZv2kR5qRKwre5VwqNZN4xmbQHDbWVlX5GI0OmX6JrnKZ7RFTvtE2dL5PDbv
hYmMU/Kr74gWTK1C1eUMs9qzOIcA4HibJLDL9vUBxTT3rGtElfifgBTiS1ktKWzGgmQ+C0pIqWFx
o+Ru8a1tL65QGGQoDSBOqLtHvB+SxD3d6484nUNd7/swpo5kYggSqJMghlkTMtWWhcAWY6YYcg1Q
S7EPfd9D33jqdgE9gdPCGWXOqpv+gmvQlVgt4+K7R9aYq5lWzZGHJg8+GQg8RAoe0CKB7OI7c8Li
vKV06XmodncqoDJU3LiKaLUvaivseliP2Xwc4HF+Jv0bvFUHiDPcTDpBpAQWdpD5kQVTiXItHTNf
RW6nGAHx8jBGceA3zfaWWN8C/0KVmBBuSEuTNXuDTPKlyAWsfUWx+5QnXGmgkW4G4mDpCL9XUpIf
wdPELXpIY16YF3DK1Qs+fAZ3ChkSzfzB/1TZZripLe7dA7l00eyryyiLjFF5pVbIB2Wp1MQD2cRM
tu1vxDaBI+zsHVw8ocVhIkIgj8AiTLinFqvDF0StlbEFhR47c6kH0cjv8JBUhQFEgMjLX0sHcxXT
1+mgW+NcvVPtA6X7SZ91RODtAa4SyOz8rg4jKcF70HfNLuBFRFhSoZANPZgawHgG5F4lDb+Aw5SJ
EZxl3BgbVdOtGjx/rm/DYy4Y8P+YUWlilVC6uIS1xcEQLD5HkYgkxvK1D8iLKqp6t9/l/TXvUnvU
hemXS7Mam+vQgXMUT0J1OZwI4P5cnr3mTYqzf65BrH9asK99hhQEnPFNbd/2FLmmEkoA6PG9Ejce
fME6m2tSm59pIrpYlGQGotACiwg9k2Wntl5lF1wS0zqwVNZ05o3WHdt/C/6NcBdCayjnpBvKkqZd
f4lPkIEaMqTKEUhvAimdkbJA0ioj1C88dwU+GIv3pJ7NUp1LvHXlWZSFMK9XhkLt1c+OxLRHkyms
KLnr1ZnnBr16NbNmGUPlSQUs3gVgPVTZQGOfCvZ/9IVK9ZHqfdCBmczvyZge1GcfH5Os4r0t1Bvh
wHX06TOUX0UijEsQn3GEgCipeL4pQR4x9vvDry4hed/9fM11xQAxiim1UFjCMzz+FaPb1Zmt1LbK
dLPJMnfZPHwKTmzIsWpLTIB5NcHjgV4bPlD7LGbQE8bWqMO+oFimWNIUI8uhuEcT3xeLnRhCdy8t
uxIHL8LhdlJgqwXN4CwW5EK9YfRm35jpXK5ZA6AFRnJ8QpgoMwZVQdm/TwWPKHrVPrBfZqjbpllz
fYc15vvaGXdnKs8wW9xSePsCF8OG+aNvZJXGBabfQvx7jyIc/wCHn3uEuVQ2AqyQ/ckmV4WKzkxJ
9CFJ//Vrk9V/xZeci5Qx+4pNhTryUjvu4InHvFhHyg2++JcrZo2YU23wN6Jc5P3gwzmIZZBNaJrg
65g2m8J9rZdOCd77QLaqm+sWi4gSKiDJr+RYkgvg1RQCPEVTHyhR9q0e9kG2WDXtalbSk54gWYtD
YC34gQpEFtcNYonbuTs7tOUPmd/IzVcFoxmCKMVpIsjZ5ByhYsHymZl5rLWFx46UrwfXMlY59jcv
rmbZcs0MZgevOkgwtcZ5mK0SUO17c5WDv9c0pGw9IpFUkmMGVZF4R2cEzHxmLtalvw95T5Zwi2NI
c4MKX8tXAUy1ChQ5i0j0Nu61uKuBW8ShOnmYP6SlRbVDVDG3aqIVwSm/rvhVQJ7KVV+YCOrdNkwe
zDlD1G5yTV47ZNXlcx5d80aTPdefVzuIAStcw3CrUs6vgKFmbCBPUi6ALaY12IjEb07YcobgogIz
SBRv/+3u9m8i+C+zlQcaFo2sT5khDsPCGs8jEinB8IpOUQJAYe0aQEJJ13stHZzx7SPIC2VjMGMA
iFw0kh20muNfN6pZxx9E2o6aOm58zc+/9smwwIZPpjlXsA1vmxMrzEkqvd9VxxTmpzgnizCS5+Yg
MKYrUqb6la7Y8i7uH9RSK1r6trjp8w1teza+Wf0RXLTSXhOY6kgVfNa5ds2fwqW6jN9I4OefmLr2
66duFEKW0njC+wA9wudlNBDTUaI5nusEei/k+gjeAyYA6dOA2W5EPmEyf/9Z5iW6UmP4GU/Hd2eI
82hZx7BeBeSvbvNFgfpFeqDRgwRNT55fnxsOYj7Dsiux6pqG0oocGxa9gu/dRJcm/owkS6A4+g5T
s5st5Pc80z6u3w5eREfXRpYYPUy3FaLUVxE8SNmah76uPfkxX/ldqRgkTna48oPftezXv0DJegxV
voVoUHrYGEt2pPXsc52mC9KQ5iav+Q5I0SglijdYKVXJg+5htMQf+jbDCNVqhRdht8XPfi/u7oip
g46kflJayqgH/NeNAAKWAU0D/IGCgX7outYlLB+oyp8QjMv1eArSSTP+QD5b7df6PZjQvnmPez3L
lBab0yMAaD3RBDu7YKy/1nud7GIRPfTkXXKWYvQQpGwFg9gD9FOge80TbvvT6ebh+cGmzcgO7P11
1n0+Zn2f8FWLSooOU2JJaCC/yHreut4a3C6/1ENCVmhSA0N32gnGR6BfFyHp6+Dcvs3VpnQCPzaL
ZCeJtpLp34qw0yP2qO/9RD+wPrnFzTyvX8b+z0KXzmmPCqsCf2OwHto5f0ZyyUxZGqRBBt5E6u+G
4nL7Cywl04T7lJFa8p0tT+GFk7c/0XkSgWV32K51rXbDlK6aodbsIAe5Oy6lg1rBob74on9hWj0j
UJrVl4nPtIod7yyA04M8mio81D1ohasVXd8tWZvObBhMS6085k+bV6297bPRABEf0qzbuNTL/oXl
piRDebBAssN1V2+AaiUg3r2EWvo6oMVteFcPsC4gnOCoOTkSJWf58h5EF7dM3Iz5PMWfOLOYRXZ3
6HrREITjYPMo6Nzp3O/PA5FixJ477zsreUeCuQzO11do5kiI6YouhngIfHsCVGi/8BMUMQ0O59z4
FYQmM0vb/p9jyDVWLnRSwzHF3oQgz7Nk7yOy70aQj+AXWjS1sIUBjD3wNmwOr3fjVkd5LNXDohax
LOelXaqd1gkxlXacLmG+GUe0JAv2JuLdhPonZ+X7a6Rkl2EZOZeAYt6YmL/X9HCv3u50NOTDKkxP
iACr1i8RqX8aZKQSYoV4VLa2liUcfSDZTIGBq1G4WfQGHSAXJFasNH5vZB5Q9ae9FtFh/E76iZAM
21iPOoqc41Hc8N/siKWPeayLLfoZ9NY3mFmZ+MuInl1KLAEEBOHDYb6DmBGtyCzpZJ3r8u4UvnZx
cWendeVEjJJ9ypxH8oReSXuISZzwnsJhZHJg9uCLDmjd63NgdnKarqGj+Ml6gET7oQ34Yib1p0PP
Za6q904SGNPSPAetUIlaPzcbd1hHmaoG1rAkNukQPejT+CsEoKBA8Mp7a53RUmXUnhz7fwLOrEN7
RLUIYb5jw0+W8zPBj7odSwov2XzU+EWRgl3L18S4GvtjoBilrPkT0Y+eunW1f62vH2eN4c1ijY5U
rdnmNc9q1T5tn6Wgn7bafo1VW8RTtvx953ijUsrkbq0ybV1LW5cHQSJZVTLKJ5vFijprWUd/gv0N
0Q45LPER2QX5WwQGPgekA+ce7Gc1VMcB7WQzJ1lHEiixTmNxwF0iyYP/6+UyGK/r6CZ/tbmaQv5j
3TKJwK0mbdlJl4QDZXMGhzIN8w+Kv5wTQoGo7g/dmNMeyLCqIoNRZ59IpD+vhZJUeVSGTiDHtICV
MNmTsb7Mh1b1g2lwxG4W7Pac0g64bL23Nqrsze0BP6ilA3oi6xlKxxt0riAgbUg9jmkfaD0S1t9x
rdujhjiNEb7japEGwcrjvsSP9OifgLIMygnpMXGta59F7KhAy9ktQffJhDzJBEbVnaAZliVQfeyE
MazYWBcdJVaEHz9C+0Y2de1L2466t5nL8r/bMscSpDlapjaHQ3E8vy384XglJDxGWn5eEtuImaU5
MdHI4rpeKHo4F0otwkiDraYf9mR1RlWrxHbvrnhzf35Xkpp+QKw9Kt6FiDy7wNEO/lW4Khu1ukFU
HZmqC5ZQ6FsYrQLtdK80pAQSul3RAzsCGEac1ChNdy91LvAWDqYzDi4YY5Iyufg6VntS75vyvkfK
04wTUQHCIuKuzDg3ILk0fCLGjZeBHJjV3Lt+A2YTBSOMuLgBi1NZrWLOGtDLvbnQi7csitUi4SRn
wZelLIfghp74GnuWVy1rbdDyLnwnuenUG4FvMum9xG7F7Wi1+G5vbL6Bm1JEok8YxfDTeGwj1UNi
f9PSW3jxlG+0mfDQQzo4J0bCIk38ivJiyjx935ASMF0gnv8AjzYDnMYjpomqdLqh9dprEKOiN829
c6glaJBAFK742xSaL3UYTF2bllB9uKJ08seI7HaUQcddwnvi7zWjcTMTLlfzUWlpDjxLnOgDtZ+m
YRQyuCq9XRl8f57QyJzFfnTIYcXnS7nJGJO6AIWwOXWKYXUbf7rjgJ0kiBchxjgESnN0573usoMa
fuecV20ct/HZshxQGGpqQhbHuQHjBLccV1AgYujuY567XWXeIzoQJPnzZeqvdegDWvLK5n7Owb0g
rL56EH+CF930WbxaeErrEnmXaYjmJFWSK4HjuvhRM/twlR98WLxBE7d9V0MMC9tkKe8jQvbBovJL
c+9n3/jZ1+DQpjtAG2loQfMFB2gIOUvrsMJkRIm+rPy7Wx/ul4CaX+nFx5nqhtk5D7irMB5k1Cye
s7JSmjcgdvTpiK/ScuDmTFvkwJt8v7/e2Mi3srsAwlQlQ8bTZuZciiaheljYGG3JzBMDqNXBQesg
eDunQjR0iwhkhQIpZTfmF6Xihq7NiNGkF4TolrzXjnkjbO40dbFFUZ03XhbpEMUGYjAofNHU88RY
q2avtXJrVrwtcnIdkfYhn7cQiX43B5Jutu0eeBzMZKh0c5nIbxEBBgJnNnnTv/PPibLmxrmT7otl
9dLQqraN+yU4Co+pPd94cIQFQdVa5cSa9wQiegYQSZ14JzXxorsNMG87JCHooHaTZ4J3+KYwcq7+
ib/wQitIymgIF9Kv3PqQlfQOo/gAqKWcyoFMoIjkj4NQ2SRSp/wabvU5cBdSxfbwNT+e3vYH6WgX
5U8RlFBkwhhf8k+80Is4WKfmx1XZdad1IfMNP8esOgfY1uzgC12ffn/BNUKFGOrc/fdPT9PNFoj0
ZfkcrGhhcjGPxye6B7YD5sKJOdvk12mzpfQSFp/kTydK7usc2m4ronCUSqfGa9+lMjcUvweRCTHb
Gk3DBim1dt9w0pJXzBlId2yNlCqDG/zKDlJsnZNr3juS/pneOtOhiyt7pPI5HIYacJN47tiSbFWm
/3yY7P7rHmH/X79dEu22Qj0W/kWFH473zeheOzs/MkxHYZc0sM9Pe2+/odniuzsd6QonH9vhr1O9
FyCILAk53z7awzB1NSuKOLFENqFdtEogUF4UaV3CF4F4B7QYF2gCiCtSWAuOILiJ6an/Lx04CgFe
4C8i+xlAzNVlGq7HJkJOn/tPwa9q7juv95XJsKiIHCtiU2W8vI74BeKcOP8vJkNBzkY7YzxvnKDd
Cql116l0FoO2PqtAF2AzBJK/6s5QjCBBkcoWIXzPMbiVte4CKE0LuFJQBNqW7O8Gn3pCb8YWBSIh
db9XTGH9eP4R4LVzm37SJlRxndLSI6UOFV6uasD33CmuI6S70f3DbdoL3OLEGYQARMGTk0Uk4c4+
U1uwgat+em4/p9sGKieDCvtycf3hg5bbcD493iKU40x2y3VKtdnZ3SxjEVyde+FqhEfKaCVlmQun
UW5XVFzBf+1XjtcEzM40g2uq+3+SRGTDhfSDbGQ90Hdfp5AcYMFqtPfdl8QhGnSo+xxWSzhlARvV
At4E8uw51S5OSrYRKAWU9MtqgDLRE34aj9oQPZNN5/j3/BSGRhhIG41a0iqsormv7p4Lod47zG8h
Ysai8/IJyU9vtDIJ2n+Pn5SKW1DqtMpvUqdc183wk0NhRAz5lCJum5bAdGUd59qmSmiwDClnSuwN
M5oTSjMeQqXATo4FBdteqEWTLx3DSpQIL1LEKqQ+9GdSsEOnj5i4qmLnNl2ANaZKhxxGbEj1tdTO
ix6w49hmbDDLexHPCSgh+UOXnKqgzBUtXveTgJLWl/R65lm4YnDPuwM6Jha9TaI6FKUBCVkBZsf6
OSlq1q+abRLd06itWcazp6L6Q9H+ve86PFIgI6aPDEAXvVbaelVb8S3Ol/qeuLY+irXHLKpoBTPo
nbmoLSSEbjtSkpsedzmHgZKQz/OL4UNEB8kcI35KR22m7yLIHhJAnH1hFz1Gr7e7AUscxRuSDZUh
tBRAK03v0QwNTfYfeOnBq99zrsSyZtXFaatczesyxp966bFqezglLIfIo4WVW9O9HhEV8VUCuzCa
6Y5ykO6subd8V171mDS9hWZ6VyxtJpUpPAOs+IdTdebNAxs/vWMa+uv6lp1CCXcQ3dWh1tcjxBO8
5cXlecUxSoztHxXitbOEab8ZNu59BSraTwj1Xz27qAxPu8oamGKTDQHK8KNHsb1dVRoLZ1FKZnkz
ggLTIKvk7HaULpd88pc47c+57ukmUFejFaH4Ica2KrLE/yhlhDuJS6FEIWIfLc6yrrqaUBDJiSwS
mf5yLBZJQvU/5GebJ3d+ncebRldYarYBckIdUKDeIC5e79BBJHfSnxMpmsDodo4v72N5gQkJH2zN
7OV3glcq9XUj16BF23+WapYj/82plmcFGD+ZT9PzoRxhO/z5y/jvcgivVgJlDlDujXlAk/TNJeQE
xHK1XGsKTqCBX76g2Jc679GcOzrzLxvcDUr24/aPZU6hjBXURol3m9XC6FQgbKkQEg4tI4+n349f
mwenoVka6FmiGI1QKuTzD8fC0+Lb52mOZn+on6XveOrCcLz7/pI5HVLc2NfVAcnQwLO8pqGOJpWD
khSNBRtsFISJMJXu97iXwz8mZrs34d6RB7FxBQ7MY1bl+pjtbUtK6R3t838UEYOueSFd+VU8MRrL
XLKDg9YTXqm97VT6f6/vWxwPjLPs0zBYL5yferCMaElzOmCtxCzPQr1bhEfYVJJzgveQ36FGl4qG
VCI416QYEyaGsGlUGJYSmjnYDTiKm8XaIggrb6rRqkYx4Ka6NgIYm3c8fCRg5/mgRCEN/vT6+nsY
1esAd6gZFwRlC0B2YTHG9wKOZE3a45Zy+fMbcScziPjdXh/LNw8fG/EOLXWIZWoTNTpqtISkLJsb
4rZIZnpimsNWQcV9nWAaylEsalB+6wjy4Vb1MT/AeDC38pyfyC9wsr6+kdvinGyyMOt4biY77zEk
hJm9mGJnKaLAi280xTiu0CWfRLw0eRUxCo5YenfMmRoAzZliM2mJBDvLZIDltgZw1VzOSfRShUB5
XXJeTn+K5r2JZcqsEqUPY44DZUwhHcxtAr82bj3O9xH+gujk4+B9coNiCcyNb4X2nYfSnjPyvy9X
OUmYdL4YzSW6CfRFPjmbyokLSNL2xbtpb1RaZ0/CK6AlAmEsqLpB2VSvCIbaYan2AmJjyx74D6Jd
xC6B42wG84jMiG9G9LNdXAtUzy662xk9BY1FfLsbR9a8JW6Na6zikUIj/nFgHwt1zXyGBi+6Isp8
fLOdU52V2+1+B5rNPrvaNIIOBxEM1977QoPmbyODHDCf5Llm2cL6V62PtGhzbKnsH4G65WNVBUCV
Dj+cZU/eGeNpWW5PvvCvtHFrsODGCZCO6EwvXy+eRA8qwue2KnbfpCwIfRgxtRyl1hyf3+HTniS9
H7K5Vmyd0n9I7+oZ7K0I7hOyEWcvOgrURswbt+syX0qff3oDWXN4MfovknJh2Hf/lGVnQJgarQly
VJbVp5w+u+B+YV64LtUrxwtgpBO85XknWdB/nI0iBZaOmU1oyGEOaxGlaz262LuJczu2ACdnnbmY
t9kavck6QVp98ekCiXCi4SM3/q9lEzhxHMiNKdeGvtFHvnLvApoiZttMNpYWqjhDNYsLQQDwRRC7
K0fGHmolVoDGQqRaVqiicSl1bSnqaiiMsnJuujUOzbMnk/RJqdVQhqDWNvNjUReMl7K71X680oCv
37HBIHRblTTdomPYxbbKDGiWOHW5beAVpKC2LKEK8CKRKqzAEGZ0VLvln3JmURmG7PFCJmezQ3FA
EQ5GaM4ePtTLaiBmP6pcOsKZxqLBufp0b+gcV3SWcxQlADjZOlHQGmx8CXiyvOTm7mDQqOuPa0T/
GU7n2aK+lHd9RO1ibjBE5vaCH/yzyd5LjTDScelhqcB7yV7pA4rmr4QqY+3S/KR0qu0wR5/mqwxP
GKt7lhrI8yaSlDx26l1NOy7V7pxzdn6shv5QZeSSVhZQ0vexRuTwjzu5q5qUv4ofZbrHuJljJ892
bYQMAus9VOzmq01WBIP5z0k/SwtHjHXg5CBf6dRZnPSDuV92NjJsUYD7ArSsih9UxDGMFA/qoTEj
wD/DjNSW6IKoQHz9pgcRB+F4ngXnTi/OGDr62ZycI/3zTMgs2YYWxOP1Hxz6ttXmRQZ7QToWeHdT
J7jD4wUUPuv35nF98rsDOBxsT/1mh6WA1p3fw+r0QuwXUci1RSDQOifenfpuwl9B6Qlz1EyzDyyJ
9R4ZzYcfsD9RgDUNCo25ho1ea2Jq0Lv+3oYTnrEg57iwMrUswuIW/1CFAY+80t+mLvICq4z+t6yF
HhQkbgKJoMk++YDennbrsjt+cBl3FkuNULucqQuyD/RTXnWc8MRey/BNeCK1Ja8RBzVVU4NAomFq
MNshUMa5J6+JeD15VTtS01xHb3QXqf/x0JZBpJ4VUySwRzCTbQZx58uQ0/LMyp0JiQsTc3kMGfd2
ArCUO7a/e6QZ00K77LDbFYWQW0cI1+L3271DqYEximGs1Ap/qCIq8IWD5GwjeAHQYaYvBzm/Yzbe
MrmTonrBIl4hwLeXIIo9x/mBdS8ySsLt1NvKD4K3LB5+45Tztx9H58vNAcQjqNMlrvG82mvI/NUQ
AaXUy7P8JoHo1nMy8Bfgc3xkL4JvFEeAyrpt4WLEX6sGrBGsUxGLoGnKbMhZies5Wq/w7k6hHLO6
irHuC8BRBNSLyZ6P6uWXkVJEELw4kXzEEzRMZo1BtcrCNLm3AyCBDmQfIqAyzzY5Ah/k3F6lWe+C
L/1+I95hwZgoqlChpUMCSm/GHEHN1GX2jh7Y+NrbUA8ZOs0h6vbburw5ff71Xt0orTssNSNKsp5r
qETRHRE7SKQOztgN6OF6zoVfwPzelbyeCuEIgmx+FAW4AplqBMsJPCHqtqErC8dMVksYPL5oG2Df
jaolhYelb6h2zX/eH8H0rKj/je8VJpkzC4wc6k7dXgtG7QDHwCqUDuYIUroXPsFtxoVtycXiAWbA
BSzGt6RBxvZS93B1m5VqzxfIFFmFE+cGTO/I9IyuHRaksNCWnx86qT8sexPrzOhhjba7IxR6k6R9
5HStzpT1lxp+w4ESvZh++xHjDXg87dcm5ko1pWNX3zMJCtMshEHUxdVbVESDrJV34aie7ktyI+r2
L4Yc9+/fvifVUvSs7/x+w2LmZ8fAWrkaJ97ajATmUG+QUidR5mBQElVIvrH+xMVy2gQrHdRUrKTN
DMCJD5u0f9/2aHeF+jF43o4VC3oIzdmthAGa425+NXzCQxX9xVoToatuH3aJr0+FrCtgFkfGw56c
uQTvtykZFwZT9lutHT3yAzJlSsqCEWqzuU23celhv22oBsX8Xt8wJ6i94Lz5fK6rreKjTiYA5qxc
tIyREPeeD7eLaKMwade2Ha0EhWh4aOReb2wtgxZNQ6yjRFDS4dPrm4xIC1pS/RelBkVJT4PpZad4
qcsSE5Ar5gpk+6PzxR8CfG2HLAMVVkSwIAATRMr1RN/wki8AjjjCur6P2hB4E6yavnfMYbIHaWTV
TRHe/p0gbnlRPdpHh2ddxM9Wpb3aZYsCMHIu3z79Hz3QaGxnATdM0D55rJGocfz25qnSgHV7fliM
hgTcVZ2eEx2uzDdqpswkAT+EWBo4W5oTpr7M48v9e7vmAP11hxPmfk8jWsQvK2ZlGF6XFQLeT/Xa
FS0gJWpqax5Qs3VlqKKreAHvfUgZSMuvZohJu5S4i3z1kCth42GF7g9L/NeGZ/KXKB94zY9+5H6p
+BmA+U2XOuQ5VTAWn51hos+tjzTcLVeDs/JIXcEc+5+hCAD4fR/RBI0yjPD0cabs8GnRtJ5XDmjh
eEEO0c/b478BsCy1cRuPqTx/HjsiO/X//MTDrGnbsZpsvl0aHafmIis3Kb9yK7uyZ7plw5qZML8h
M9/FhxYhqsBa2b+lkKDwdBGNwtbZ8p6tT7dL+8Zyj3bwpRBm5zcOKFvnFU/9ZLp+7MUGszKQ21p7
FTcHAKdtRppjWx2C3N/Bhg2NUMZEdTFcGbxqJIbX6emyiOnfeaT7z+pUp3IDUc75wW0GTduOzRgk
3JR6LRAeT7IqoqCyhSIUs2dmHhNcXWd03OH/MhYfhnXuU4ZpHnMAv9jPBh+KTXcSWcSOUcY+bKuu
REs5ysqN/HtV4YAkEkoq/vGTu5u3QcCTooCxz6kUvvorBeEh8tjWm6l4BWKiTJlKKARrwGA3fpNG
PQptRcUz6FVqkDPt3tkxUff7cOQwt8czoEzr0ULZGklY+OSrnc/mxecxVE9VnRrY9S7V4kGJ98Kh
K4RbbZjlO48Frfe09K/4rWZzGvw4jNrcKruIyKfv9neaP/lV90XxBmi1YSw0VmFMZX/BZ73CQUxR
dNYCB7EWFlMwbdORNqtLy3JLFPBpFbV9z0/KyQMrtJSlWRB5FDHGUyXM1spcMR9CvscK1seLo1UJ
/suU6TIOJMi9urw0DHGF6AMQDXeIBNvrEOMLci6xL3AtHhj3kAz60NbjqQ6Z1gCh6r5WpQPDo0gH
3h5Nr7lrXAc3fRNgrYLXUFi1a2fYB/MNydzQ3hETHhpK0E0KX5wSjp6hCzrDZXOt7UcWgr38vMPe
gILL0AehDCHJh/PBYjJ/XceuVzTkPZrZ0lk8mvrvDmQb+MndO2eDrRFstkLx8kPLBB6CB7WpV/Jg
vtV4MP5Zsac0w2Lhi3pKEzF7B23Wk8Kk4QDTG+BMNV1px8j3d43G1qUsCks9kWh+Bj+eAhE4Fe9Y
5ceoaOGV5rldu9b+JKlsoDTSEFi3YZByOUYgLT1M3fXrP9MPTstTTizQWqNeyPbrVR0jRVoPuBFK
o6IbqOa5Zd+HZx1sXUqi7/udlBuN5z1KSDxjxm7nj/1YIBDFtL8xTVkRXdQcYnFGIr45IhJx+kym
iKKuHxAoGgIUcVH67Q5Np5Wlom1xMKo19EnucpoZ/7ECsHl2jgW/oKd8HOfKXs5B1sObwm5+BhSw
Tk6068/CzMSZPo6NvptAb6VMj23vglNgEuBgLH1m1tnmxMvXxXmBz971QIGJGgDyvNB6ri+/tiAw
2iVayoxm0ezg4sDR2fdQ2uldVs36qfm8If1VDdU6spTn9bXjEfsZtEvNZC27L6Iu6EFtYjV5klNo
yG2IsJO3W4WWXADP/UmDAEzB4pWmBdpmu7ZDufsdwwjWgaAlGNrSkQiPmMclnRPQTWZceHepEi3O
tFbtMdAiDNWUT6BHbGzrSsMuSBhDjffW6Q/KU9cgdPuylMRIWI1F7hIS7G1tSAoSA8+1g6+Gb8FS
ja/hmOVX6m+hj4RDpq6ePg6Arzr9E3CuVFRbvENOUsiq8me/rtruC7uqeRSaVXaLfbXBXRa2taT7
53lnPbaNmbCkP813rqKsX1Mu4pvm6bXFM0KOs3IlgpU92aNDvijPEFm5bM26ocXI96d/i/R+Tdmr
RKef1F6W/rhr4WB0IQK8a991e/D638yMYEKYaZJwlJvLGtZKyIDe4ZjopLKTxNZerBCkpE0fxX9o
fMRtLgoJhXUdsunRVfiDV4+YpnLaAAOZ0PbRajJCegXaYkFqSETRnnlFsBlZGvm/ljRo5Qr0Grqj
qMKFXlIaMOgft86N3OdX6r+hEOK/LMbKI0SrNQXJ1I8cRaegFJMGRwudL8J9U0yMZ5+r3olwkQUK
IxPZdjhnVG0kLCtiBWuygsRXickEJbMCf8PDf0hMqyY+2+MJjiAYtNA88S32ktwu3duLG6hpiZnp
SrJZgcjREtSDGlIAzBQhm7Giyv5NCoUdJOTdjUR8UWhONagOvZKPGIh+ATKoI8ESyhwsYb/wXpad
kfDBcJbJG9925nFInrQtemkDZl05TbjdFZj8qLvx0CPKS2w9lGp6LTh0OWvR/aTdEZCetaVB7XzU
0beg0VisTePAvAa8TujG7vQqCj8srGaYlJSAJmSHGQhTl0ame2yerWFkNjVNYeYEd191JNrshkyY
neYNGOC8eKTsDz0DK+CBiawa1KoIbCNHDy1caQ+A00Rog2GcwhCooO7HMOTBZucoZ49JbCXZBh9S
6HCGLEOs9GTTG7o1an9PhpDb1aTGHa90OF9WwRrNzlXJuzFcOBxNZWPok/egTaqyAnsJukNrN1CW
BOqpbYUm9BjpqV5ycIBofxl+UPJLt/b3BxXUKPJfSl2bqpV/bthTtEn6OGCN7hLrRFxCES4/evDF
t7ZYGUIuRfajFKos3Agk1MW6Tg8b5QccFtEcfXDlkk+YREo4Sm2A1rODhW5wZe2wSlyhhkLODSy/
xpzfKDlSolIG6Eq4Lt5QLdQMx8C01E5NnpjwvbhePNPqqQqkpnRtUI2QPw0tUSc6DTZLNVET2NOx
aK/RGdDmq5yZQuqPVrJLUvbh/+yp1DiRm3q5vwr8ehnZLup3wsCgumDWRX5XJvVT2zrzp9iI4rDj
MvEWOY5+LUW6b+YqNxA+XR1k8CayOAhkndDEGVcvl3oCTBgWv3x6IHCeEl7PvLaN/e8QJH85M5uK
79em0I5CIl/I7r6Id36LKpGZstFD0pntlzjtxD5cQj4IlMJJHt+WElm2Mcf7CikS8Y6IhSdJ7duQ
gNgpN/avPXjZbyu0NMJonD6dGG+1EFbfn7u95bULcXaS8szLehmGzk22nyqTcjQK3YyIW//Q58lI
g9rBXm86KrhyDTo5BjPHvuOIaWMh72XmeNDpBZocNVdoBAmhSnMUkjfMRjfPpPXcqqn7Cl2vzcNN
hArRlq2eUXvLiatPYauSYR4i8HXplDh8hMMQmyhZ/zsYCpEF253rX1AHXzX79jXBi+3gS5SJ7oRw
VKz3TnTxnnh+coXcNHgKTB5qP6K0lfpjJ6EfHGrKbD27bfQroGeFyMfiBbUys+MKG6d9rB5C5qv1
llVIhye7GcVwIgdgUoSlOLXEqRL/cSxSxvvKrRnim7S7vKQVekRZAtsJWMDTNZx+xd3YTkJVrrJh
glHsvi9U8nvfwbEl3/Qp9dJJEosfdJb8a9h1osKhAbE6HBg4EuQiyV+ewqE6CLzsKuRFDyayopI+
Bi8AEJyVpvCC4JX8AoZZLqQxhmmZlv4TYhYagAVJWG341ryncteNa0cdclG4/s1s2XK3rcUx2vz7
ZbPsq1BTwxWZZDxznNOxD51SYL43Mq9KQKBTO45L4n3bk5xI5ghD2BHYUrrHPqC4THF/3NkUnPXs
9SarrX6TvH+EFVmNYTvyYnrtjD7wblq42qbl2r/HnVRBYnxs4fylVbgYrukXhj56HWyf/fhtJUUs
devCs3vLyQiM68DZWhVPf3OwFchy8ntMiFa9XqMnxj1tUCXxWZ+FXmL1CNFwtUPqJjMt8aXDjBWM
yQbI0YBC+0a46ohRinGsDung9mFFnazEhfnYl6kB56U2GklQcADJwK1w66d2JCz4anuqziiBH9Ue
HKZF2C0UIODgWEZHR7Vaq0o/UkY+La3JykXwR/MUOV8+p7iwhUY3LdBMckbfVXJrLYjUKcyNinSP
9EPPq+KNRtz6OK5P8y7qihtzKjTZuCLKsvEHXT2V/R8jE9WqneQRFrw6hvQfFcyqiFyFpxPfS08X
rUxMli1vx2YfxWTMi3z1JyVVEb+x341CxQugCDZ/HWyBcFIYH3QECWTpa2EfPk9AAx8ewmiflhnI
Lzu9Zhuogfz22djhjiZUTSab+LAWLsWiKIApguHMA4mkm+t5Z4qcV0g4aMfGyTeyucltAJNiorGM
Aioc9JQ9R6CCOmmmbZRM+55gPTGpg4H1hNZnHLU6Anczl3BxXqwPBoFLkORkc2gQ61Y8Dcld+y8K
/qGUw4KavRJHXrYM3N+KAy0OsxC6LEHloWhCMEs9bOIIB9kv/X/hf+AQ2xBVdKpWifIk6xCMtkxv
nDLDY5NJ1qszVzx4rUH7M9AK7mv77n076Zdxo1+kMmtAsARK7dJdc6EMgMA9Eu02ihuOY52igGw7
1/NBaPY40BPckORjPuv00jUmQ/vpbywH6oxTS7MK6PJxu9og6h4iNTP8ssJeHHpk/IIidPlF2Ggf
mgtv2ilVv2Ye0XxBvKMW0Fbyu23nzDMupZ1Dr+FmuZDXmh0pRj3m7sdxe6KK2qLy97qJzrLpOPry
wEu0MJV4Ip6VBm0PS9yvSMZssAWytkFscw6ZHuGDbozXGI1dyTuD0wIhkX11SaKBkqSuQdzzVTYT
SFT1e5Za0+Ez12UHnWOoZwsRQSLRrwUFI13SHza3sDN4I1kk2NaAzCoLgfUXyZYYvevjKpB7TEZ9
DG7Xldz1ISpGsTxDSt8wg/6cZXKBp2LN2IT0Bm32ihaU+MRnHF+cr183yrBf/6cYcc7YvGCI+cYM
d7xUgzN6pfEM+SQiyuqWMJqA0hJ0glKo/MxAtQag6RbW2djrEcqR/pLgJjZu/7xkv/aafJZYnp0M
oOUxyXwUypuH/pd7ey+T9fCBX4sh2y0yUzPyemTW43jiAtOASeIuAqio/o+U5nI5+rHKZdTBMDRu
EY6L33CuP0YSbOuPvvfGQFoeQnkUULk/pABmyxEKJ7wAOHlit8TnNmXs7cPbERCjAcaWA+mwfR44
0jH9CgWjPHSZU23k99SwrZdQSJDw2IdujCUgES9mA7WS/uxERHCDa4pNkSrHkEdQyKr+06AZND1+
5UKThkBBBS+4cxtpzQmF4YiIc0fB5uNpawhgF97DqhZkXYoIksfjpokPoF243sfKzTcFsZXar/4r
M2knxnZIDHKPT+A4WEFDM8g3xYNQPEEhF0aX/QFlfQ0e9JxAUG4vfm+5p18Yfo4Zvj6QNHylZ0Lg
z1BimPSdBzfTmBfCqBfjOr1NgPLt+/rDKPzEuB7maqqA3DBZss4ISOU0jFe29UGQoA9zKYudeLdJ
x/16d/rIuLAH9hKyvutakk2B3shFfEwpmbyi9I4jgh2xYsCSzL4xuGX3DK933iL+Y8dfx03D70xa
VSpKJYR7J5Vfl/xQkTfZVTpS/bEIF965735pOo2iz8jUBGHZevy0gSajLli9WX2apuyFWk42aMm5
740lpAbXN7ut726jxKSzMCblBPdXmIJE1TWOtIbYTrpbzfnqdAyOfhoqiMfv3DuaEzPKHTPuxt6r
n82RIYbUqSJXRFN4u7vlbuVvn8LNw+7BfcW3zGw0htqYxM2iO/2hT3kcsoKIFEHBqE0+fdEqfryb
oq8lcJI2sYX5sIH8yNBDpluMfvp+yFK0Ce1PzNJTy6YqkQzc5wM4RriALjJcqy7H1UuvBL8Ivhre
SbR5OhUAkfiRbX9SsfYqgOu/JVW7/oQe4mfStxlWmqGwNpt2Q5AuQGuCZQ9wHfSYagN2lFpB4dz7
WBs4weh/RldUpGKnzRWG0+HfbEOwClQkVNGSMLDLwmM9YyKT8ZLYcZ+f1vMU6uqdv3dE7GHM5Tlh
SJW2lMej058DhTNW2IJi5RNIF8jrmhlIUm0289F0UyP7Bc0XUmqJNA+5klbAZL7x0csAfzDL1Ara
FmH0dg3su6+EpBMSW2vqDE86Lh7qxcdkKSCPvfXqpjPvceleWSH1NwVKIcBkpgWR2MYOoFcEn5yD
gMtWuc+fj7nU+DPfrqZ1oiUVb5Unz8RaAMx9SV/Zr42WHakZzqMF9VZv/CjY3PAxWl1vESIAUSV4
oPwWOHFKox2M+8uJY1jUsckURKV0YUDdRPNnXMsZmvn/W8oFx8WOGMOitSeJl8rjAwq/75pq6IwT
RU5Z9Rt4tfj8fgtymm7Zmm6hnaFdctxX6apcgr+tYmMUBoGeVLZhVZJSiwJowklk7DtDcUaMlW3C
QkCy4UZaGGPngmyGH7kcW6uggFmWekPlBZAA7K84JYJUsUrZYEd0A6xdMxQq7h5y9lrGRwdzeUIT
A734fBQIOaZHHosb3GOWH3H3hKMuxe1unXe9DdmheUvDqKRfyQ5491hG5BYF9gR/LyzxzM+tF3Yh
kceqHnSXphojoIr74R9Qgmm0Zkw5QbhGUpj0TFe8jvxuxRJdQNv+1tY4uqNO08k/0i7OODXnkVsB
xccAJNGRZVnDRXr4/kudPcQW4zj1pyjjTiBB9hGe1C8P0T/CuylkM1OXhnDq12zt2J7Lhfdyj0HB
bYLO/q7iMfoWtO8KstOtOoV2YIAy/OHyaPKY1kvlg6VtOMyth9mmcntgpEpJ0FDDhgOCkZ5MAwn3
jmb8wp/iEGAHwiXsffKnO3GaMRwz62cKtB37phgxDBvx2Y5A4+sB/A0rwkehMxqAzlxK/lHY1sFA
4zedgU5z/VkSTBUraEvf1zOE4Qanvw80JgAH4bRfRLTjHcwp8az8iCdYHyOvZeOcBf44Ap7ub9aJ
dN3Kk2wh7k6ig35tudg/AAUo/YHpN0xim5MuIOaWdmNNwV3P3Pm6iJgHl52+oOt1qO731XJ1QwZ5
tSXmI/R6bdykIhz2zTBm5gB77x5twc7b62VjQDQkZv/bRqu929aDUghUNvOj5za5IjkUpWdWj58e
C5oo9lO7big5IYNHTfsbIfIgCiYcKafIC6jWOzdRoBPVRuQ5lWPoOFsMfYiBLdpZUoxBN4cDVxMD
lkGEO2c1YdOUfI6HwYJPUE1gBdOJKsK1kbhA3vY8Py51tvVOewpi0/jE26u1OmEK3IonmBwXVjCF
HAs5GATXNB64wgTfY8ViWV/ebgWNzynv2Wu8hD+RaZxxQr0QA0QjWqo1jlbIGb99UfAQqUcoZDRz
AQgIIRN7vq4drPcyK0Wumwywfh1TrIINsuhLMIPt8indSG0zeIWxBCLMchBicQzXoXoEhd19I0Ha
/FcHNdAQYXjoCM9XCgFVUH9+EKJNUaPVCs9z/VZGysMH2AsS0jvJpoTlWMcwMsWHpagzbfsiS2G0
QLUCC53BtJGNkiyjoRg2kxPLV3CHvlcqUekgGs6tr+1wmvGeJeDnKbFtQ91gFvH6txxPbLQRQVwz
YXhNq/encOzhmDTuNUxyueNdHRVkx8WUxL1KQZxj/4dO8NSV9V2SstDBLrA7BpjlOQIhFGyfxALb
9voFZFpBe8blpgqy2VXC8B5A0vnSV65A8wn96GTN2QMzOtCVS3NzkfhaK2V1RqUQUGELpZ48emLe
HlmNDSQmNk1pcWRNJZeFA5O0nEop97CltxwTeyQ4qZQUuIZWtGezrCOlfEu1r0TtX3AfipIC/Zn2
Kj0dmSe3RBrJUIqH4/YWf8b5ZFdzYNZfSR0KHKsfeMRl9dpz0DWR8zWuIFdBw+bAldGDgvXpd8yy
/A/FtVzvPE15yNg5LqUEn1XrT9PP1R5/qhck2zP49kLikRmf6Oqm6wjrEUfHOFjCLAYJFFNG/y12
2tIXGc7xkw1+GcCyK/XeuQyFVFwLQzjOsQD89gWfp8MKmYU/Wg8JwSMgKygQnzauDHxzqUri0LmN
cCRekRdBgdFiBI1V4mScfXk8LWCosZKx7PlJiPLytJ/Rd2uvlPgNWWCG1NBU7bQ4cLuUaH3/plHQ
LO5OYe7Iqx+5LTn0x5O80H4ek2kUNkz+lCUM85w2MN7cWjNDpUrCoDBpQqQIj1nZnBfXtjv1/+Ym
LXaGz/ezDmP9lpBaT935XPpfSPxxtXuFRiFIm3m7iqp1GLhzeqiCeZogMWO2dXr3u7OtAqSE3Ket
h/xxMa9Sw/R/EkGH38+UccWnMydOSJrGp0gwBuIMVqiMX1GowbwvaVqClwPBnROwiSp2zR0upppO
uoLDAYV+c0GxwLUoi97aOKPHGPmZpvCDcjIViNNcr4VWPEgwfmofp29P2S0OXUbrGmzHlqBEQvYR
q24N2YHvLs/CiO8I+NFmmZbrEbccs0C4quyKbTBnv+sHv2ydOGVCVohxw1fF1LWCxUr6JvMSTAet
swu67QLjQ5/ZDHQJH7ga/HLYTTUIPMsPnVZ0biUWs0SkTbazpcjWmnp0LB5cCqpw8REZCgDZiMwh
rJT5HU1qLunknkR93mfJuDW2blWuQOd3cgctjvjxInxQt6u4/p0+HzjDruzKEGn9TMjlSjh+FE9L
55a2adZt8jjALq+4MY0wJZHbNsOS+jEWRHG1txxSxxwWuCH+Vi6rwHPjxoQFjjiXJ/4VraixCkMF
/ktR1PGiHepZzRJwrwDXjQlv6xK9yPERIngk6BeAJD0uydDl7lVmz19yxhMFsdijRxklLo2nRXnF
fB/gwNtP57ykKqi9RfUx7NAZ8PgsWNXbf7UPH0B0epBSDl2OMdz12BM5R8gMKzUPpZp/d0O36EDw
APXXvoynX1H2ZKmSaVn37zYJI6Kax/jNcoqvAYRxB1usSNHU+/gZHviwfJhxrkOD2XG4L2ycf4B9
ggotsXYlMW5MFwf2eVKi+JYu0Md0q/cAAyH8TRGkzuXV6jVGHKSoIsAopr/d0oCoEobdEIc/xDlx
HqApyaqf/xTyq+4DRGjPS3AE1vFKPOginDVlPvEykszdjOF2kuKMPeSnopp+FxgU+y4lYEAHVobw
VIlvG80a6axIPTmne1m3KXahZLUSKvFMvIcwHuPxBAvbGlBtuK+QcxlP59bkwnJdCu9EF1h/V4vE
j553sOQcI95+ByA3Afj3dp6Q4Ox5POHFvW/2uEDVHKbOE/hq0Qlf3Jl6yJYET7KLT/IcSf2jv70n
aSPiGeSqxDW2MTvyZ4CHCfgMnZeJ4IBHMB8MRsigdb8BBc7Z9ziccKM94sBkH/b+qE28Sfi+2fbp
4XfwLLLJEc2RMeZsQSRQ9zvPqVg7TtXEVFvHxDthC+yIj/Q7DKOT/b1aUcJ348irYrBWd4yyRctw
bxFfQX2FvwTy0P6Hcl5Swa36OB5X1+jMJkF2oAnEqdHHkZoJ3phbh67/orXT7Dzwehgz8QsH5rPJ
aAuA55GsJ7e6N+R3NecxpPxASjovuQbpteYjAqb+62pKMMI7MU7M16hMcG54JzOVoIuDfyGSbei8
nnm0dYSpW6JZ+x9Z34G94u20wPyTCQL7/sB2iOHZoj/I8xORWIKCVPEFi4WpZZPPQRNgSL5Aseel
bD9Mgc1ThEcPlE1csMFlkktiN4dUiW5ZfA3OKMcYi0CkTz7QZAfrnlaGkBQa7wCGI5SGW4tFifKS
6TQSt4vrSto7icLEJUibFsx06bBuZucRPKsvQIEo2vZVpwq7TyFhyfn8jKUrqJ8dgMMLE08iS7Bq
KbNdGSJV4gcbCDdbcvNYEqh2opzjmQ3Cju4HSO8Ckdd2sQE5+0x/bWHA1ySchdvp+2ycci6DYOl6
cA7aUuDgtF6VGNDhD/rhGpfFwigZRgxHUKBlGHNn7SL4hjkIJSLG0tupjUYo3ev/pfsN0BKrUh6v
8H0M+YS1fpTtnPjO7CY8KeWKczHkeBhSIKzmGcbKB4GPoNNWSLP4KNnRG7T2p0hLlYZcxCvtkeyB
aMlAe828q8QLOk5VKNg8wbFSSxe0I4S0OdkBO41DraMYoir6EThun12XJttd0i1Eyh2y9ErpEqzZ
4heNDUUdb24HxVuVq27OCVUbfnr4QpKJFjyJFsEnT+1dUjAtKmlYNe+LBr+zNSpI9oJV6hVAe49q
dH/uXAYsQgadiFXRySJYCrjIQXceRKJE1dFbH5Fxene/17W0T5hfvWp6Uk7DkJqRSHhs6NH7gDjJ
12QpNpeF94ZfDyEhzW2avvTHyGA0eLlA4FagACeXOyKIaQfuXk93z+2gsVq51194bGPPFVk5X6xm
mFumZ88zLuaC81xdlKCa5FPXC4Vkugbv2cQZi+nIRl43vFV348jVvjHBvrgIfgj2MLTPtl/j8XYc
HH2DlPrn85eE6JqkOZ0yGuCVdvvlR030Cn9qktSRcYz790f9i2pe14WeocanvK8UWWcsyD5kYFD+
E1l9m8EgJdpON3vKJGMF+UOqqqzvm8JtBu8i6L/CB5R147ct44rRUoiTYT+yesmWRiURCs6VVJUW
OcBIXcyoA2c/JXo13ppRvYLvkzwNyyEgXOofGv9sSmabUW+1SVoH8iC/Yc7mybi8eAYNIeliVW5J
tQn8TLwq9jVz9d1wAz2i86QRQJ/dtzg17LMmXJSlWbzimnBs+8k/lSt+5zozKmg5946s+3hJu9WS
IHBK4bJ7ZHmkk2tAx86iCXZY22oJiC2LQT+CPWsROw+LVJOLcDNTS0Y2fepAZPshksUPxtb9IoAp
nnrKqa1/pTv/4HOTevkZ5JzSiQdg76igLcW7DNKt/IeqOdsv3nnlRtaCExGZeElDy3iWO7d1fKWL
RCKNyZOJC1jzl9+E1Q2sD2Wi+rjaVvZbRgKL9TfNmmIVJTuOhTJ9DZypzrsrNlIjH7Cy+2J8P7ch
IEHS9fD/tnK2G+8V4pRbXOZ1QF5Akay6smsS0wf+rBTceTw0LjZ90d47oz/WAuQk/kLeK3lLE0U0
u5Hazb+zG1N3KPWJlA0s/KeyzqeGnUJ/4m77nWrG09z7Z1fTt71JkaF5g+4cKhhPowpkv4tQ//ow
TOWmzxgNc5tHLApIChDtmV2BGNKFVuxxGM6IFVUI68prp3uMViE9TvXDi2ke+Z71bYY87Bcdr+nO
pQC3ov8d59STH8FQNeZOA+XAEgSjzs1n10VcZc7PDyZjgH6m5bK44w95jHKZvI5LetdtW0QdTjyF
j1O+sayP88pTaUQOvZR5kbi/bB1h7mnDq7lmTwOvthzSw8ZanGywHyqm7nDjQmTLlja797RHEhB/
ZN5uuX4oNxwtv1Rd3R0diP4wOfUWNxi/TcnR6aS0lF49khGKmr8kooDSo3ayRKwIz60UDIMI4E/u
P9pttLA4PaDxYNzOvzUl+t5wUaSBPYfiFjgtm+npLSqaLxfKOLUy/QPhYEM1BkpB5sjNOS6OIlD1
udpiGaFCHwthvupAe8jzTLzZBQSkYDVGErhr+QFAcYjkh7dD8sTHGSEPy6A3cP7LV9E1XLObClhK
QnZnVXlfRmjEUt8WqabbN4CZZrILcrtsnS1SkpNzBJcQBEhjVzArpwZMpa7twlP+R/F9Ig84+6nL
7+KF895X7wqnuuyniVZwlNxu9EtHC15YnBTmZPXqq/TLeiPSc4e/K1PTFIvU6kjDER40OYYIiiKy
elODMGr6/XnSJRQp9heag/nRPhjnjIj6gf+s84pa7Hqjxwz/yjtYLMzLcTEtHKhki41g/dMDhjW5
oqlqoPT2yNL63Z75o+UWndS2KnY6pKLcHPQxRsPUY4cRGqC1CItlUnfhftHkq2Kkctkfy16yNXeB
NnHQKzaGuWQfN4TjLKQkzgk8qxPwj7LRpgRGLbPJ2DsJ7xlmEDJLpn+F+75H4k+uluZrjC1N1eFM
/S08NQicVMqYh0NVK0iDzHxl1p69Nsr6V3EHYGXIFpG9y32GtZetCm7XYWVnfv9fKbhiEOQVQOAr
9mJIL3SxHnCYbgf3l8piArpKnVU7aFc4D00qjltsMJ9ueqAypEBaRLMY/WjHuzMkVcgPbNgU158D
VoHkih03XF8kV/7IYKp2KgxzFxBWAUziYpdrp+tEOiVY9jXuZZ4Etsp5fplGpSMOJkVESnrBI/jx
1llT2FAk7G+dcYF9YZUA+BpAeccrSjklDl/hY9xtI12dNr6ceN2/TgsZ3ngB9ekn7leog6DJd3Hm
Sp5eFxk0X8/RLNqAWZa9ipH3QeqSvanxJreFkPVbNG8Nz5/VOFhlrSje1okrb1b6rF9JKGFx1S2J
T6UUkVuurYKZ3aPZnlu1V/6Jg9oFWeMpnP9v/XgCrfET59rHRLwUdTtnqKE3ztD3aogY572i3VTR
Sip1Hk14taLXloNRbc/nWcPw8CMFJqc0jpI1CMzVvUlvS1r6Q251MYtlFrgJmQ3go7mn+WMMfd7U
qENNXCqoOSncfHzkATL8dUSLeKMBGJUSuioBP643ddHyWiQuHHi8uLDGQpzSMTJ8py1ViCOEfbjS
HgYZWA9t/BaSx3IaSt/e5AXtNTC9NGdK/0OFEK6shXtkpcXDzKfYbrXRj4lXKgaQsnVulybIqdvY
GbU1BF/DADntipKBYXhWoS3ibu43TnLw4xRrOFKA1P166j+3Ez+ddctDK3o8g1ry05VANPVnplNa
IhL1+J9bwbfYm18FzEbHcNCbI1DepJNI8EprRDAbVcequZq5xYVyotqFde81DMeTQGWIneve36jY
ROm9agQrWQZ6LrWD1v0we0K0ppuOTIsz5sWBbBlzuWgvINJ7QntlibRRk5eC5ZKUuqf8hBgTbdxH
t2DG651IJFjft+PksXPXeoqWtBSROpk7UkbleJXD2ZsvddaQ84qy7iB6QVL8UjKHxG4GqanIeAgV
F4+1u1ozVoWIShfVSMl85jzqdjlvleXdzf6XyomMRy8Tly27DvrpdDqTJeUAw12lvlwOt4Pcr4N9
n4QfOdOKMsnLutBtZDIkX4B5jSSnO3+1sh1P/qtcl3rqWIsvl3nvf0cb9DUpJjePY0QRoh3eGlhB
4rPwZl3C2Wzcn1TZ4kKVwtixZe6SYHLNpksq9crHNQhWEm1i7x/tY5YvSXgVX92DQPkCf8wkEiD1
PYYuPuWJEPmX5Zx/9RmmXLmqrmi0JoMa6eZqh5ndkIEGmTJvDxV7xrTC09OszSNCb1lGaxfiLN2x
w4UqK4jKbo9okt7vqPFWKcKS2b3uIMKZqYJjgezRaT4yor9WI3u3H22BXOEB6CQtVNWcKlWjc3W8
jZToK2ukaKEp4p2nhOJJga5FOLRr0OuuVBAy7/ULtgL2wfXOWYmWt/wbyc4Zm/7dz5mQI4hABwyk
X+fXKFL25wzqR0IBtNSgFxDzbvzlr9E7Fqp3og4h3xjLQHs98oRZfnP1NJSQCvHfwdkls0RQTBZ1
DK4AH2HQHylt3kOPJeg4HDCdfpYqFEkDSR9PYQwSpWe0vp25QMgwM7mPhCor1RAGL7KNytkWxARZ
rXGygJet1v/NDKZ4M7TKMD4AV2pvAXNBwg/Su0dWWIZCh+AIgeUDea3Qebf4p6l0RYBMcScmXxPx
yPLn6i+5xaU+3wUVpJuYPnm0VNX3Abj4atIYCo05guoNCu09gqeutg5QHIGbI0FcVqmt0YDHgeik
V1T4GAkBDhWHuFFO0KOLknMjNfNG4vAZs+GZh1b11sjYdm6H/mX+drkGBEMGmVlWT+tGqlh+cQIp
vM8l+1/e7yWZS+dLopbLGlojP7OI0eFY5dAioeBaENHoLoppRNnqbPsSWZASBBYL0Q2mFTnsuWBX
Hj8Q1q93s0ahOPkEpV+N+5yLcdEZTpu9kBSSkdKrusyElwbu4iUgeCU8HpHLG0MQgSv5DxgA0Ght
/yPVJI1fFtXt8ppJkOtcG6FK1t4CzhrUFRZVnqyB9nj3P/HM3KoERFKR3zUD2FeHhxAq8dNn4zW9
iu9v/5+KOL7E0kq5r/tvb3XCSAu0uEtTL1vXXMtyNIDxXSirY7A3R/J0BcWU2wrSuCZbfCsaDYvv
j6G7HYAa1xvW783p84kQX5v+oaK5JLElyvd+kYeukFsTYxD8rxa6c7HPIN4XZO6QEXWm4yRDG0Xh
ghBoMu7OOJ9alpna0yz9NgEwYSdSPVg03XS+v3kBtXqMI4pZtWxysOo/IGKQNUDqh3hbl2VEAoql
7HypxvftjhkSuFryaown980FHfeHFeK4XK6yaD6AK4+d5gMmEP5kygbdUy6H+wMtnuZO5DPQr9fH
sOWuhU09Ff9Z+WQwjkOLvKMV8N4HDU6yumNGKHw7NLalxAggoaIBKtdNhvkQUFM4nWJPVGG56/EJ
E3i0dKxWbn2CZMqRHJh1rdg//CPKOItMm6sKYfxAxe/kOkQ6Ic8I0SU/YpHNnbrhhQolJjgIm0fy
zcCLzmdJycxEvDjgh97u0sHzvh6+ReGpMhXHaLOp4yo7aNsYOXd83Ok8cK6LJfOTVRG9fatLaEWH
P6zTYYVVSah6tbpw71HrApDNpciaW0OrC94wSTcbIzrYj1jYhctRo+PZ6sTwSzcqISIlcstAUrwd
raAT3HRDmP+GjXnvVxV04/TqgQ9znKVaKVsAzS/Xfs3S0lE+oA/QI9QcWVo6o5Wo7LmSe1baLxTX
9PuchhL3HrY27R1dXp4f8Od9gQdnDweYIvXjsY6Kl+0vkCJuFJmnmM7dOdOlORwEkLC8/KOUeuSF
nOQBgdzEnqML59vy9w/x67v1iI3GQTmNlUJjUptAPfq0NRxKpCC4buKY1/Wiv2x+wbJA3m3bzpxO
gvscON5TrAmv5ZAsKaYSVbkrjbOk8WqMTLX0T5exClnAg9rJUNdu0mFnDn7RJu1wHau2nWmacO5y
chQgl/sCnwHUsuvAPyqa+ISPmrajqOUHwx7FUvZXHBPyhCp0Z4eJ6DjE68ARY6QOcjWHMk2jzp48
5Ij7lPGwcTJNb2ZQtDtC2nUdutP1XdJbyLSoxlDQaUbggxuzJXqMsGw3F3HgkCLlJfLy6YIxh7fJ
GJk6qg4j6oFgeyqKsx/6pfJPlDEzA0Y4p4PcLLEQQRH0FMiwMsi4AjJI/OvL8f1zEz5u9Hr5s/vf
0pImmu9UMdvty/RQJJzGEG1dU8hoTBfp/EwczJEDUg6f7ZxW1gC64qvPL2CPNjVe+1VAR6qaMt1q
4sOnCmxcNoV/4IR//Ej/83XSBiQ9YG+PpYNY0cc4R+cx+YJg6PTt4yhfk6hSNzSev24Kx3PzKNTb
tlA7J8PFYQ34eyKUXe535NxRn/wS18H52Z0viafdFnZTI04qqbxSgiWpg5gE/3PCCt/DpG9usIQI
CsrRfCWhnsF3FIKtlJnJYyKpEGhIJG8jwfDDN8etiNU0srTHFPTrhmG6aOSEyaEN2pu7KzVehyqG
LHE5cfoGDFpCdW0QSJntoJ2deBH2wR5+EEuqOwmRZkNWTrxn7t9HByfOUQ6nvwNMKwWTC0xjjUeS
t75prA3IRRhP5aJBaDTo8QKdrVEw91ZCOLcAURqJjUvxmXVYt/pVB9nmi+jn/aX5Ds9s1/61R+jF
LZE/VWCZ7DcCMsnkDYT96I6r7YQ27AZgSgmzFZZSYLwmUlUDM2mNs1TmaGabNcnPkQivsNtKcKFU
El0K2nmYKM131+XJg7U2vxL/TW6R9vhIRgLeIuTsxguDfFmO6bi2NV2QKeIQ5bNCeoacFEwKzCc+
6HkP8zhak0Mn1rDnoJ/Lg/Q2O84wKUC1aVElILBNZFQO/ygbP2lj4ZABe0Hi2+oOmE4D4QqdviAB
D5UCQE/mrSmvSq1wr41Hs6Ie2i/qVn3KTSq4VMxg68TIHMw5CabfyoJ+nfYWW/+rqC97x/CLNkM3
jlzt7HQPhXaaDSLzpnGhrO/fqPkbXSjDJ8viVszuhnBH8XtxLZb3kcrEubyesauGqV6gix0Q7Avo
w0Pcg8lT7OPZyXLzvnTAF5Fs+NHJtqbWyLrBk5hLgp16GFh24D+C8mcn4qFI61inOVIqTwv5nGmj
558fo3J4gvE1ftuRLYDg5P8ZBs3Mhz7eZWKha9RqsE12uRXb0mJx61udb7DPWC6bKCpGD8uLLPWM
aLAEhS/6GNRSa5ZlUg5O8TrYiezu8PeKLQgMGwmnIC84UtPI3b3Xkvd0fzWRAfVkHnoI7OUtZLNK
tGKurj4TW3DN/LIW0s3e/8074Kvh8ksQh/X8F8o3E1RSYlfSeAd4QSBj6DoXNH22KymOyDoERd6U
V1kCheuH+3ZhCoYSo361BdULsjbV1JVxkO98sh0aisgqhZZDtDQyPP5POQnmQP970BKWVT0D/w3u
HyeHeWIHGiXjtJRWwPvkqiJh/G0bn2OXTYjd03xHkEIuC/GXZv2K5zDljjSaL27anf9rjAalSUPS
brmqBRta/5Kz4//wVKzOsYKk1ayX0sbCM3MQZcnyql1B9dsSS2UDcyHuq3Tch8ViPfzudwhlMVO2
oKuUBb6L77ZMcrbI0RUdn4MLIDAuQKvMfdY+PuX7vrBmVjZ+M42MP/AW37fd+/EYzJHDB6uNfoOw
Ob2Vob93zihhJhFKiZhVxN2dcZRxCv1gNzzzn+QswoCKxtkgSqumrf8fYQZy7OaoUNmvspthwWiW
Rn4CvQcVGVJydctgnCRqnuGwXQhpXW59npmwc6V+rgfMbHGCZ5CJ0+HDU8mW3f8RiUmJNIIu47RA
BE+qoTGVDbDuc6Z8VKXWDLjh8Dbc4xbrKDp3L+X1SoZXZLd+uHDRYWYpKxWXOLznKUHJfelpulQY
80xI3l+4bJKWmmEbpaROnzoDzGFWyOE/4uT+p0G/W1DImXQNZPXTTEyUkvcp0mj0mQipwTo3rCsd
OFy5kHaZarHIvA1K79OieFp0LflnO983jdm+9GoDQH/ZfGx8tNErqJdb5XcMZom1VUkL/N0CMy+3
hWTHLF32BC5eKLlIX7JRNRnZuV4v4h1uEAZ8OG5T47VWWl7Ucq8IBa4/R8YPrQ77clBUK6eNMPSd
EPi6GMYHyVjMBoSo7JAlj69H4eGB7csJtKk9twjI5dgLkfv33zNN7ySmHs1Y/eQ91jS9zpLuOV/J
Zjt6kOxFHOqbP2CnI9B7n0ZaG3J34b+yHgsIygzRYf2qEtB+ClFzx4sKk6tQif+FSXmqQ5uXhwhD
4AGWNIvZ3qyFmTWjIrlD8ChxL56JAXln1Z+qzVIjVRDvvQXicOH8zQW8IIMefv9qfo08o5JeBJDB
xUA/tJWCi02u1+BkAMoESswyyirxpi/oklVdf5iAjNReEMWLKz9palN0TuBcG2M9tCC8od5Solr2
dH2Inif6/I1M/aodVVSOefMayXaJ1so3Dn4LpjmRjwh8T/NNBNS/JFJKcfUkcPEEhQaKVr8pJZ+Z
MQIyPg9Frk3KKunlfroZFiXKG9PMYQnUmrvIMrgEKJMN5eS5S9cOiWC6dJzHX1qvQK00GH5UXlkh
R+ibxEmHSLITJd0ZuyPDCYo9XyhJ3Qu94vei0tBot1yLrAQ5DHFWqO9eK1yMdqNiu9m54CLZFupJ
ZF0iT0ujQkgl6WpohtUDsQ2Ct37NUr+3LJbU1PuFrM6W6gBFL2EP12/SIT/ek6aQ1rXnoFU35n4v
UdGqy9b97dURbpN2rhpCCdUW3+wfkLT7fvY1dkL34uPwSQjM2ynLdejOHqXti5vz0xaUcRioEfyq
VnNVpIM+wecR9BLWyFGe3z+1HJZ+AxHKXtvMksEdVSio5lQOse8UAqiweqhbqC09gPSW0Ak7lFiI
qJQToEPtx5WkhpOA2ZWSXCTGgTj/RDUbVYKzbn8a3bUwahVUgujf5m/JHauAXuQZQVi2HQbZv9NM
bSb7025A2zC7AqU7OE/ibfESiSJxKQ8FFr9StowVW0/aBq3ylsXpzvblCQGE9bebXPMgrMV5KOOO
kslEQZumIpu0PSmFxClvr8MFAJ7BszVMzJMLd6CZDEijIYIgbdpbHL6wP6LhiaESOjsF5zdN6O70
BlegbSlP65/GGbvLglUMGc5muNhCGLsaVGR9hZHAbdVw1Jh9a5vNWr9h99Wc91Qqfp+UV/p/KvtU
twz9Tx7xN/aynPXlD8wyUpoeOkVxJqs66O4ts6lp7R8vZ5TJo6OyvEpDC1bnja70sbyc2/5qRABd
zLj1L4T7O/IpLd21apycKUPo8qwvrjGgDfIzSgiz6lWp8nm11BpCqEpu/OsMc9+6icW1qbOZQuwa
LL2qGqfBwRDUbvjGCnXdlY5ishpPdDnV/iKP/MD3rNBVI4J7rrqZ+6JH2O9jKHZE2BkNDKHXos5Y
QMdBIb35wcxaZ9yJDjAIyiTNXuNLV+LqWpClWkM6FdrkD0ECL6iaUdxFKhYMfrb5sOpuMSIsFv/q
zWAE7Jtnv9pMhrESupoQJjeAZ8NNwceQLFqENbjSJysnjmir7MhaIWHoxLTYd/RJQ7Zwcm90aEIo
bSPTHvO4KOZrc4GCDXe9v11JqADl/929xrf0RqUgFTx4LZuoGwcxdUFfpxnhypDROY8Q4Aa2wHyv
rFePZp2CtYfb9Vurq95gLda1SMHZ7/D+t8e9yLrOrJsglKvpsFbMi8zWS12wotITUlxvJ60XSe+P
e/Bb2JvXwFq2W+7jXy9q2oAFItbdJ9zaA5mSOSRJ0Daf00Ed4sezMa6SMZcJsL5Jgtz6Se7A2R8L
T5Ah7WKALQ3LzYbdZSWP3C01Q946VjGzYguVoPZyOUfK7XYo/rSYfmY2sMsisblPH9TNpj9rwVke
0SG0lwzlxVmFUOv2OyJPq4MzYeRahCNLfL5B1CGZ+o7YB7F1xfCBP1b7GEpqN8KV0pFAMJJ8gESU
hp87OGjW5B2HzuyaKj0nhxQ7m1kDjxd8TClc/vnUJfnQTPcRJBbezy/poJWYorB3rzBn/hHfURhx
OXBqk9MJOtBJPuKcvQFKo+paDNTMshZ5kktopQWCTku+/QReSRU/c9GCemoypt6S/SWn/UYinNI5
tVXTH9Mb3Ty1X8mtj9ZYHhlXAfDBuO+ndSgko9s95yFLf/hBcjckpumjIKSkhcBhmuy8hG2WFDOh
On5VAod4kUm/PHfm5ChJDjsmULhGgJ8o7VNiSuvw8alDPf+HMVPQNqLq/MjjZxANYhcCg4F6Xxy9
jgVLk9pZ6r6uu944c2nF705GFAyWtqs+OaPYQx1S22lZ0uZlepxmZIFePxzJhM3VogmvC4oAfDKS
hOpSiF0OmzTVTyMMMZoji3X9EtK+c58PBF29P+FM8eot2CxWJV0sfhesi1mRRtqvhDNzngFWw2lN
GpbnuqD+Ox9deAW0hIt7PdgxMOQaXnmozcwX88AtheUA+MnC7m69m10bTYvdEuKchPII2ScugA/+
TC9V9FlGnuAyxwz7SMVUL6SwdH/2A2EDQycE8GsXIjnRutV6HCHgbWp0M4/oFgRZ9Tj7Zkyf9wgJ
89TkHURRRSYAK3Rh1mlNE4XkJ5W+OCWQ9CvXB6ABUrOIM6aKnEpTyMlRwcV3ZZQhjjvDzrxjJOKt
JGCZge+rGZd7FwRGnihsk0T+veo+f6OsrijBkyRjKxYxTdSGQ2sdNerNRyYVDxih1wcqOk9H7qMQ
iDMrmBAhkKSuvz7YLA79gKldjNZ/N4AOzimDzqwRrpi9egbIb2A/If0jXt0CByJ9/82T7Dq95NHm
J6n75hJ8sli1ciKQVFP4nz8qSTkRD2SfmrwE09N7VoJVPoIa6Ri/TagfoYAz924rlRtQveyTMmo2
F4DfM0ZxU6BmGdw4eZq9u6JRtWhR31cnrbFCd1zpzZ412/waoveMspXbAITvse03AglIYnQUFuSM
YO/sLAj8vZ5dXYlaZoRcr79VRQX9XTA7FJKCeIyyUryVLSyD/T8Vj2rZD9pZynGk4CjXy8qHHxLf
A3mbi8Ae5OFCAcuAcE15GB3ILvHMCtBuuGGodvDqQjn+tukP6FvVomoM9c8JpPB3khmBJTOSKpjP
vI3yLi7fl+bEozc2Zflmxkaham86T+ozCcIiXypt6yL0l5BJ9V5OKtT+Ij740V5FeWJJ3qc8fkvf
crgXtcFiXrXkTvQnuVsuJRHtQ/VXf92o9GjiYD9VKIeoFBcDEPDrAqp57Z/5JGjp47deGqIcHNwG
LVFl0564TEu2uChwWESI+M+iZw+2IYGjUCPjvoXlW7N9PgQI7xGuV2jwJq+8DbqLbcY9+01BWxGO
ruXrx27X4Cv2aTCfIeqIbAhTxM0j4s3XsM2x/x5S3bGSiDNcL/MkRgyRzBuITLXcEyjKKmGT1vgu
SdNd7L6FgZgQ9NOL7LhMKRVF3Ack0nI/uFQpq/PncOT0EXTIqrVLqu0VihCbp7F1Zcl1xnpR/BE8
wAzAKjQNXe2tHKQNLyAHcuncXsjKX6yBJQsqZRd5JI0VQXbIu08w5xNtFrGH9gH5ZAieJ+DLu51U
ygqHCNmMw7VrAbmJIUqR5s6IzJtdRDLuCX+CL8bmsqKZYj/84kRnb2aV0IC4wY7pHLU+DLsDKt2Q
T5ww7PQPL87D74pY/2ZLK2Rt9aghjNlhhm+v/RCSOgNPmj/IBDKs2w2NkQk8sZE7q9BkGOJMxuyM
Yoa2MwQsvwdR2LRKcsL0mCm4E5suHBVbHFiNo+NZsRszMvhvaEM2bWr6Bp4l+XNK4nw9TZfj/3PD
vqab0GIR+o+BuCzqKJTBDxKr3+t8ep1QlBt+wIWkzu6aaOajOCxrQpQaKP/zMNFjoLwAILhnaw/3
og8zJo10qFScsB32oIXPZWI0TOF6eapBRhnhfLs5a5rabKqfUASV/bomau+hH+Z55KzoXuSxt/NM
aV1D1jU36Z3M1PuObyUs+ZrSpzn1JiL+Ep22aX+5C18LXYEev9VVgKsnRX/juXTry2syNYRkQTku
qji6XcxdE1e2mqsxc7pmHk+G571BRKxHxTHA4eTfNSI23/GVaWUmUx7oO3Al2NqZsAhz07+ct3gK
auXP+3y3JgINrNOegsj6jFnbhL9e29Hm4wIiRTlF/QXY4LddqtQ3P7em9y2Vz9AF5u6ix7j/SG8/
GHbISqDTn+IjrZxvZ7A4mN+bk+BVvqK7KgxbOSJwzIGAp+O/mii1kDZXewrtQJqkXiLGMD6oGI7/
5iTKOosEb13gsGiZz8wWgEntZxjrHADMiQgt7lRrGaf3bAtz9S8vMFubJaSyiAvBD6LMduqqo9jx
tZx37k/MgJ0L5w4GpbjhfYHuccAg/Osz6JnoJudhUwCRNfkd+IWzLVJgyEaYNB6HzIxfPIRQqpML
cI1pyo75RH25ErA6atUT5Tqe1UvSDBzKE9FiaFOs49cpPf6njGsTQ+LD3EQr/Qn+weFFp13N0Z0E
CrfF5Sn3/Si+jFGeKO2F5BCbKlGL1Dg1kgf6Zx4RwE/CpcV6/hociTrZYdS64FM8lMnk9WWcbJXj
Nm7+mRxXiWjiW2lIQtKyxho+bWq/bABTnvQJEuG3w3ta+9OmPx/DPicD0M49wtnUOTQ6OY6dPr5W
sk73N7gx5JiS5ohNepsMWDU9PwCaF8cRiSzu1Ysfel8iR7kpKAvEeE/4ZaW0n/iYWk1BnCthvyxy
HrsKMKtF4Vo1bKVDP656I9KSJGT2ijPohVJo3z9IREExwWaLMNv3UIMFBiQvaIajf7eEX83R18K3
owgpc2VRi18n1Ax5pgheiOWB0R701hxh00gGiFy4J1tyKHUACjnVflKOOUhBbFE57IX01r/V3y0E
U9LtEGzuc+MO4eX/G3nw2KKOzd6JU8yXt6GKqr2ND/0+ILY6oW2eC4NgWvFoJ3hciWlkx8MZK7Qz
eLb7Tx52+R4eMrGj4B9ZBCqQRORm0Kb+flkA6l6pOx1eXxUTA6fV+hA28wNhPLlZdNXmIgovTLia
ajqpFqYmQv5ztX749+T9/za66Vjh7PaFKdqs3auPx+Ewn890Qe6MGzEqkG4xccvgxaH5TC7Wr97/
v1EVj8u33KsICA1aBMdkIInQl1EA0KE8Kk+2pram+NlLM+bJEIgD/HPaF0wbM9wFdxi8UjOJ8uXC
PpLkpSv1nFkN5nlE0kvgi5WNJoWLEV5svO4EXI6iL3eJ/jfVAqDusS4Dp47ZtqX3RfLEmXHVyQDE
/Da+Q13OxIi5m5aldLpUcpefnelr01LC83OtMeDIVJW2HUfP4ee9UPBRxz6846xNf6fMHsg77+uC
L+Q4XKJn+lWispmW5l9UWYkbexIy5HlJSE8NCU5ww3yuzN6mX3/HCU86/iSxabFVkwCBYKETfcR6
+lDS5AU2WLhUldczNUJ4U3YxZyy4ebP7XY1SpMsvSP4srxc48gXHOPEbq6wRSDVv9klBKPeeBxMv
kmnsafZsXhl1xB4bXo8utIwmzuPrsS6wRwNPQ3doIbX/cdjpCUpWhqLIu/Ni4/SAfOFdpk6ETw6S
v9XkqIvvhwibUqsqKf+ztj7y7ek2rIoSifgHl9b0EczQzyeWuOM0hQylbrmm5hDo8F2gqtiuagXQ
9KS5SgN6Mkq/G4GoejqstEtVDOHzxiOt6qUQFAOEbZhoxDUMol28yvQZSgs2F7a7DyQTvNXXgJYI
z9+MBYenCnwjXEe4ZQraKh/Vbm58R7HZ+FhJBpXmVp/5c6OR3MQ+x/LvVerd4C9MShFn9PFs60IT
XnV/fgPUS8BjxvGVv8SWZZbFANhhHMoxRqPyy4YVMzIU680ddT82DgxK+dt+tVrbGL2hT/wGdK3D
iCd0AUl+NrOwWxns3cR3Zdo6i8MXMueD9eyE6RzqLTx17PMgbWFILi7ZkXk/O6U9YKnIfPhOFOSd
5NtQLvIq1IcS0zRuWVuRMS9QEjDuA/2fsTJUfGntZa9M3YkzY0EA9E4MxsjT5Q7di5EsvU/MXC2e
I+jJHc4oYdXPDbvhi6oF0H2xs5xIKPuplAYLPWMwSf7r5yuSAtwmPs3SJ5smr7K3PG/t5n+ZrJyq
Iw2WBT5pCM174cnd9kZKF8z+tudraC4xEf/svwaxsmv2FdA8XpqhwSOYGpPKP2CtNwe/QiQXamKH
Y/Ht43SUbkv0gZEAtAth8OfWDif6TroE4GO2izbQecO6IixYV9B+vfO7MJdNjANq9CrbKimKWufX
1YsEMZYeEYPFd45UxDDbGi5QpAFFwEwZZiHSoG8zDK+TIC6G0mV8C1JxbjO7yUnfP7J99cYH+Ldc
g1zNMHB90h5CViKpFePhYiIUXOoiaDj6SQcaVb+RbvvzpgOTbFhpHRuhV8ICax/9OH75rWIzamfW
RktPpMU1dPJo7Jz0wyHxBeju4u7WLWROSbV9+fzTySJEfwm0Th7/aATgZ5Iv7S2o7RCGP3PnfjUS
GRFYsfEFiG3rc/jF2uFHxjiKfmPE/KUOKvZS8EsgBqonrFOQn61HNiozyjmwhlynS426lkZFLr3b
Hj/j7BuCvaXWBa35sioRSdPQNW4hWm/NMCzPD+HSlop946XjiJXJjlgKvMDCeOW5tuxy0vm14sCY
N/3v0YlLHKKgXOSvOTFI9JAX4dpiV0RlqGrWb4YzgsSDXTNLi6jAtQ/oFeWNeFTa077jmcgcI/3D
CJS6YTXZoKRxH9KdGUrxcvWu4hnv3RFA+ZJn6HIH10saK023UtveRJcIn5C8RfApIpXtyaoROKxp
5qs6EJQksNlM1xFSgyxFIPKvcNUt+O1nk7ykBJYJ58wm+Rb+fyJ+fvWOsoanE+qbFvsg7Wm2FB2O
KSRqst+BT42O1CElvpchHz3j9j0yQlxCHSvAhXMDn3yZW3rFGIGNT4PMkt2yEt5qjILJFEY1BwRI
JBrke3OWZQ1NU4SrLvAeuph50XTZfTXV5xz5e59BcsRUlZ0caMuYGCBzuUjm+Q5bvs4RUfz8iUXZ
bbt0qLdAJQLIYT97dsQmMmpAmXIovL6DlBcAxDulowqK+99Rf4SZ00gYS+GgSIbE2Hu4kFsk5WU4
QWIPNCmuog9ojkqxvBzqvjn8HYhG/n3q92y7pD9b+c1rJAU1Kyjnxezi7P50Sa/Rs9RKGjdj53ij
NkmrYKiAFzUx1roPTUxfs7TdpycQTxUCIy8EZkR7X+W7vJKQoAWxX1pep7OyFRVRW/Xe4WoOB6Hi
iSjOHnBaV2i3tT4NuI08gZ7mcHaejwfiESqwGpnAPGFfb0pcLkVyJVGAfJeNWTOBpll4ZKEZCjWX
tYD4GLRN9WxP7wjA7ydpULMNpCfc1W+VecDNvaJ+atOVKa7s3gGA/ar6n7R6b8pNYmCbNbfGUASI
FHIligw9kXuzyQr7llVMiwwDFOWPRBgdM32NN+fjPVRUQYhif7DtVnYGWy0bYt/mFHQJIxe23P1a
gZJKSuktAlZWii2KwU4kp0FQMtyBXWmnIlmweb36U4PNC61zcSH0Oiwucrjv9SX13KKrxepKGXk0
pCmXDYVpRTnnndBEpgH0SFYlA144m40cm7THIMv98N57xWHcvrJ17+Qxqt4ZaorPmU8ZneGddccM
kuO9Vnd91lL+9/la4PDYqQvyzEhmdp6SAjHAFEFIrRUPNNXxRhBL4ICDR2+uaptMIqa6l1/+HxmO
o4+emUi/Ce3h4usZhh1Om32FEMEKchPLJAzUfXjAUokSessCmwCvBvw38c2l6Ih4z3IO11oojYDe
6x9lzAST87+IKyGItt0ZVKlzB9SvYK75VDNBRhppU9rraT1FeEyl4I8TxRW9wMf/uDuKwKGvNfG6
CgPjrpQNZhu2CsrVhye/fwVMqkhELAWsvmdRkp6Fz6KijwfmKFFOrD7ZwyLJ3P9WWqYsyy9Ukl9n
dGSznS04ksKHNNojN58UfwMDFAFYgCoeBZF/w1f5seObmi9uH3ZxV0hoaH10B/nXp7NcDWES88Kv
gQMFY5V8ZGVMhshgO0n1HZx3ka/fMX7ELGNyOIVYbqxc+SAVO1KGmFP154V8tzvHQ5LHBrE6pz6v
lnMhWsu7DPYySy+JrODx/1cbagNKiXJBFTDEvb6gi9/v8YSrC+0owRszFqkZVUvRfLU/bQYwNOwQ
kKOrN7MVCtm1P/Wg0Nas6hTB4fq8ZZ71kZFmydS5d8T9+a1Ebk9Y6Fn5Aej7dtn7oWD7z6W+xTG9
nP0vOsNss9GVfJP5UiZFHk56Qf4xgec4UIj0QMIjPyCDuJSKJS7dZqmObhJwI3HQdD0Qy88AFYzu
ApmrJNEqhGGaAI5rMl2II6Eiu1s0IGNoxaUiZ4t8iHgJxS9bB9Dj6l/fWNOmVNubvn1lnM1oqTvh
SQ5TKjPnEjumiMwLb3tPIE/2HNZBGy2GPJJeEFqgRAFXSZdKRka4+xvsdIhd4AbMyoI8eDx19bZM
FA7fmiVIRDbIRSLJSLzzFWDmxwsLgpOOEvRVg1QRayLLOj4OG6R4QZMM8iUDoMNROu+p3mlpNfKb
dRcvfi0g6K/Sw6uwFoOhxIlGGTiJLEsWKZfJc4XYexu+fu8CmKOm7ha1AEiOejIIABJdEDzLmSFM
GYPEgFcsqWzrWrUOfhMqNy6EZctXisx5CapzRIJ5xBFGKedfuN85LCHp8M+Z2M5apTU+B7kzSk92
vNv7wumxZcCpnIqWnl8gHKZD/O75S1IC0SzjAqZggR2f4fD62OL8/J+u5w0b7jTkPPVrcJRop/9V
8YH6cT7+OfU7alheVWutUBj9w3XdpfATiIBMlGeoxxPLmfqBy1g9KesKlZagQ4s0N5q5Ny12w/EL
I1iwIj0tx3gChM/tyLy0OrIIkWcpzWHyo+jSD+BDxrdhJi+VCIVSFlq9v0E6Et/GLJgfM711RmWT
ZwYCZUPcEcZ4jPJeZo4/sghPRQ0fjJqeEdjxBUfi++B0NGyERWn3YnRoN5jedWf03SwSpKT1MlpY
o3QqGlihAru16X8zUTAXQZCS3gbvdNzUlIUeCwFZE87JbFLGh93hrYoJOFgm1b9XtGNLRRe7bJfO
PVdbqinhDfv+0sMcaXAjuNOf5iIOGGo+xQomvK5e3Dg/qKfd/ZU4iCG3HOtTHzNxzkMK/7NZ3Hnb
owXMHUAlkyGEodZ7XfNrRo5Jr30OF7gNgUwZtGRT5YHidxCNfci8HElCvCngfotkk1xqrsYSBDaY
cPFiJihOnQiabQwc0GgEsWWQYhRlfTS7SfcBR78S2GVwnmZK7e4s1Zp6RlAWADLVzKfbkul91fW4
1NRA/Z4LrXUGvViwHP1nnbD4ZxHZQFRlaoCB1016ij9lbOF8R8yj+nvqxohFv9bgHD9HH72Z2PJc
iJvF2SGFgMRzgrMjx7HPM5dOB0At8J2LBA5OUrPruoQcmf9JWaz5dnfTv1MV4d/2lECj3Q0u0dr4
cUzsvZGeMg5gB13qB0IcnyXRRmE/qnPRhypaLY8YqFJ78frMEqm7HarQH77mbHqLeedGERdr3JV6
Bh2IVjhDOBquf6D+VH+P+k9sM2o93iNP1d6U358SHjqghuuzFrC9TGmkjvdCJQXLXbOcEqZtitQ3
2bvpdQJsZTZw4z1LX5JW2u+Ofy0UpmJWFe0E3NZgl1ZnOnR8yXu+HoBiGsSPY2XbJDwaCZ+2i2tI
vYOKdwtjNZf6H1WZxEXlkOdDl02niZPqT/0BFnRwjTGkLEFVlxNSgJT1V8uU8OSpOjVKWYycEwkD
x+7TVPuY8OoT9pFMTxQniWqad+ssL9cQGsav+xXhnF/AD/hnY8IgjG6PA7YlSWi+HtChtKT2s5Qj
/HqQ95gtCSWW3KQAFucUP5V19R5ux7WsGdM8zxZpH6qcalkzLTWsDtKQ4MqlzUhry6CdJaSqJMWr
NU2IjGlAgjOIN3aWLkwbGTSgcAk3Nf/SA0be0dE0bmW3UaCvTRaJIVLZzC/Lx9FKfejLSBqV0mpa
jT+Bfq9sMX3ZgkOjXuzIl5LzAbUDwfytETLtAUtDt37v6lj7e2mMn4rRrdzC25nzWMbfUgQD/7Mc
UMmXzOFc6zUEZrNU600YNCd7nhJzL6LGqEWW5AmRkBU1BL010ekGAkF4fMb9FaOiZDIBfrGKkgZC
DBCoSilf4UquaIBps2CQ3HLq93XsCrOCnKZyAQ94co41WcUj5kCch6lboRfIE9sknJvrPdAOeK51
CaGiTrfqcP0f/pUQeAQWXR0a+RlKDkfP/LvFcUWGwjM3UWXvONNpITA2wAIEtOUjl+RTHyLx+H1R
sv1bQ5/xlnlQvSc+YN1bMyCIlYX4FsN/RfnMgt3R9ffFuhkAchAwjVSyyuMtNIfTgWv5yYe3kSVx
aROi1cXeWNiD4lUazI0UjHsTU7oXBVF77odsDhM2WdqQhZ7e+AVZcAuOJQ+GCeqcDHi6cOMFgzci
UdMFtlpq7dc/id5/LoQPxyT7fP2nVrne6acLSMrLf8MNk/NQmG0ZVChTUH+hrUhqxxljsqUyKIlI
EgX1O+RolhSsp4m56E6ZWEX3olZXfqwt6hUeGsZ+IfMZLKlsegahiopmIgSTytOY67lJq0AZ8F/r
8wpEtiT8SYzd/3O3ZmQKN9JqkiEG5o8eRcG8qjVdJLiPSOwoH/Bc0Iiiv9acHMQRKo+1VXtgAtpd
+LVGv7NlYMpqmTogRvkJqCFqcRAzh5qpYbD2CNHF1HTdy+HCEZyNWch2i1ydZd2rOu0nt2KahFU+
gxGiIm9S0wTaKHf/aT4dUJ7jCxoRsAao8VgYduLkELYj6aeRJOpHClGIGZRq/dpBcPzLxwAVjkjh
5Tl4IEGGU29x4PMBRGvGbHx5Z22HSIkoDnFeSvDES7l85jLPWmSn1QcyenWE7s0plflLGzjDcxFc
B98SE3C1h5A1EMNvYbt6yaJPDqBCdAb8rjo8FO4OQd4I26C+ccmgHsR7UihFO4gtI1bm5kCotj5p
1NYH5R8xk6TgFHFfqNDwzKVca4a8QCCtIueO+9CcA2HjQRtrDpbEWWuNIG2BhIYohOK0vqoOyzK6
c1W0MuHw9po/oT3046Lgji3knEHjTPDf1Ol98z6nj+cnlh1TjfWWjnKZvHNTZx7NcR7wfCLrtuyS
RCpaoQEq5kZacmUkL//bwrYlU97T8c2IKvh5/QbuWnrIRndxRzAG+kSEi3ZZuuFgcGrFcyKnDihx
nzA+H4ncWWztQVuelg6piX1bwblQjKPce2oY97/6Z8GekSwcoomMf9XgdW6TBO4enU+XirxcGsL0
r/8vqS5kbJ/54Nn2GDyybpAJ1trf8Ea1FGQ1meHnHTvUhaicXZsmQXvuQgzUKw2ZYIldDdwBKCUx
rpuNmS7eZ8NohF24Kzui3K1gjkM99LgKdHCe6ZXhGjsg4LJOBhVgUgFtzYxHWvhHiSUlKGanlvhi
mshiC5WnDHaQWD0XpxCgGHBwi3xS+1UQWpMJ1w1pS82BOANW+BxEdTUNvwLu8kfduX60fc0Dyndw
x73sVo721f9n3pr8ltABtuPcMUhzjgPRH/qJlZZ74edxnjP4Fut6yHveB33zdV+UZnXRY1fOce3a
6uJqjcPF4Un08suosOgOaX5ncppDYuKjXGSY97cGEyGKLye7Ekg2jszzGpJe8xU/WQMLV1GuyvIM
kHZ7gz4guldOHvAqFL4SZIryCodZgm894OD0oTt07ShH7rxdXm/9vaeYBaX4tBRrlD7KDd05Gng1
HgUb20xthuLnf540rWQ0P7RD8VClDfNg5eUhL7SrxqT9PWcS7YX4B4aBMMdfdZ1yosnRbG4nPtTN
zOcTy1wkU9g0KYyyLdFPWwvXryUl02hqqOIAVilV3q9TMnQbptcA3kCbhIFlLOVOCgzZQKL46qku
u3WzLLIVZOvLOEF0yiL8i1a9vOhSldkqBpWAhV5X5bxzqpcXrvpcXN+AV5tUzUhxe3dIdf0k0tBj
FGS6iYCPeCS8rGQmE315HuPHJJxMHfkOla/wsfFxNWmwj5Gb1vf2Ggqtr8FC9TtGeyVlUjU7SQdi
0GsNuk8CJwixbT3o3UrwWjk6CpsIpSYg4Kqa1nVB1XXI+2hDf6Dus7Ce+XjdUAVdLLiCcRrnKEDQ
/3aQ11YXOWVM73tIoeB1oKFFD5yW/usSKyGcw4VO/KSeWAAyMgfJOqcFrd+jyoiOBcPm9NY7W8vv
BfI0CMbD3Kt4TIYcMeL/KsYBSuXVPxNRhOOdIvS/yLfRc/WYKKvDZ20s2f45dn7PAPqWto2sXofW
wWTibbgfqv7S3r4v8K4I6DZcY4cRHQH+dV7m+zmqr/feUXVsWhl8aiakkSaXTlaQT7JH2VpJm5oM
4vJOp/yWI1MfnKI4B+sCeIYYoq5C39G0l7EUzsKFC0c3Gzw9d0rfejyiYDU2DkccxrhESgJ9fpbH
A4aZ1sb6hIZ/sKxwNv6GDPlI6kKJ9ScLNSFRYxZPg2I1CaLvhDEYXcQz8b2lDjfRWf9d2ItjF52/
qxytbVhnd4U+gOtHBc4ynZitQgw9wKPupzY/+uVuuaRsbAH9VYOLhxWRY2UNVJ5sUivtXClGv6hr
PdZHs/k0I8ObdaQUDhmfSbRZPMFXsgmQpKQCoVMkgfHMCwmsZY7PmuLIaDiMx9UOBkdLg0SFOjvG
hhcvm0/4UabUS3E6/VCYsMtOp9TwLktL5i2Dd6Dcgv0uS3Ql53ZiPh1GT/OSAICvhWKRDuKZxuJr
g+V33eGx8G/rpDFXjFZz9Xvp4ytppWGQvRawKzpdA1CEMpvHrELLLR192gYrI7vG0r13GA/KlSgA
Pl1B5CnoIjPA7+MGwn0hHU8liugX9xjBqZB+bZ7+8++MKMUuQxcpsWOakRexzMhB17ph8NLDNAjv
DLjqniu6DooWtwaKPSRuGU56ZvWSuJbV7UHwKlGDpgh0dOhmDUDPSMCaz45Ha6q22MAJ4ruwd84R
9iml2idos1tfzMPzgpzZ2JpUHsBp/cBnlfgEWpsraXj/zdpkSSUeU13V08zqud0mCzaF5jg5aldC
lPHPTaf7sv4h8DqhX3ieFnO/O6YczbCjXBEbRpjYEoJOhdno/Ypg6wAgie7auYf3lxmpxMcYthb3
S43LoRPsUqPEjGS9hW8DMCjuOJ2Z4nVZnAWwYAaoQhIqfpFKC6XxW9DVAKHELpb+dqgfcEX20dN1
UiJcAUvTwyc49RYOkeKRmMTBYYm8ToZAA/zqmlmSQgXOnBD+uaqnKMJTXizkE6L7Kz5lBx/qOANm
+GHiRE1KpnPQYxfs8n8NrjqCYd6Z3panWX4u8wQZspiog0J+p9JqHKPsDcbzCZ8lymdnk2M3Xa4o
VwrhIxl2CP6fMIsaiFzS9lk8KuB1BGDwubk+HQ86pkg/OKDNnikmYJNMQETk6wZSJGXltZnXq/3w
9IB3lY3DVe820b3PcrUAlbLe8MVX/2OivI4RtDxJhZKnPwtwjVfUY3qomfLhPAUunlislJ30tcvO
8n1n792drp8nqgWON3Y6RJBFYprsYnrZCeXxwNRVt995uils8gwJR9P1BRKzO4a2mMk9freYZm4b
adtxUzYHRq0V1R2QJkzvad9oKS9qZggwikoQUdO/ZRZXoIwa1Pc4A8fO5JuDpzyj6cndsQ+JDeES
XCnoNslBrmsG2eNuTo5Rn8vANFUJlcSmyz02jKXA2L3nCyH4OQFZmjZKX/Ltpi/ozybXTF/5VsHa
4lGBh0oQmUSwZRXasgJxqpgMlzfhjIc+pEnr8xhlOG8rNReAWHg/dRZHFwOXq6rTxLDbCLjcZ4Wx
5bSIot7oTlppCY0/Zib+Be7hlhFfUztNntv6mCWPSBPNwSgNRd1uy/yUjO+h4fhaTWMHgDeQ+H4y
U06e9am62hPv6blPcJUuQpqMGr/acFEkuhGAV1kWDs0UeECqffascahCOmRamrj/fzgJoJU5ZRfk
He8elGN57BB4gPIVWKuLDr/6uYpeWwW9C4KSRQavePSOy9bdsyrG+Vttaejy1t1y4r+Qhk88viev
fe3n3kL5sp+zcriPGTNXCwjoNH5N3EQoTss00btsHsA5Yz7HxL/Urz+j9HutOTpdQtqyW+W0moWX
4LRNCky9I8CWJLsSHs8p5pGWcfqIugknL79w589HEvyxesBsp6rMfKfiJQp1n6rp6zhj0ZFz7oZz
ZUQ1eEKJZ1TTXYP22fczW8/1HbBBFqkR0cDWiMPn9CxviXfrpOC/IKp4N+MRvlotwLQ6/IMnalih
cqzTo3kJDe5qBIJ85t4/tLlFIfxgLjB3vAekm9PtG3R6L6F/s3R/Npk41ZM47IagJDkiyTEuDngY
NyApZo2tJ85jeDL4n9T/aRBcD/NOU4ciVeJE1tn4Xcc73u0Z4WixcbZoIpcFGe6RrlsLqDeh2kLb
Y2FFEGq6vi4wruFaRHDOPzQmbyqowiov4K9o3yt2n7MFgJm/mqE8qcruHygjvZhjwuSrslgya6+L
vR/LKEMaGPRWNLTg6dsH8tNKNBt0+K+C8FdvcSH4ZKAJ+YG2RbFIZdeJ16HzSqolZiBl4HrQVxMX
L+PQ0wt1C8OBaPdi7pMVGHXv1fC87aiCYkWGzr5YtfFQ7a4tBxeNBd5Upqi35PdJX79gBxPswFEu
gRiO8sxkybdv2EybDflzUPqFpyGGkJ7QmNtE3qt0co1it1MPMdhewrNy3BhKSffPfSxQ8A6weI7u
XnfaBR72t8tw22PwFH1ZoFR92OicZOEwLSS13Wmj6pCr3rbDRbrPotfpDG96Clal3sISllI8RQUZ
Pd9sRcC5mvTKxf5NuvpDB/RPPHxvwn8bikwazvCFAOerWfgRIK1gTsUgKcGGudQ797QyntvH9lxK
4QZ+3JqfMzlMvEuXa9tLe3RkcZ6SjTaK75HS+YtIPMBqdmMbf8/C44tcSaG97818w3oUyssZHZoR
VS8gCxLhek+YMOYXzvIiHMUuCyvCFNNbnypw1E2/baDxOXve0o6l+0WRVP3mkgkB+OsBMRFrDGG2
R0qsk7CxQFLovqpFTZ1Fo3yDqMYnfFwFROuMDObaDWC7HSegy+oAoG7NYdYEsxZ1XMgUQzv7ki2x
nALw7I4AxsyD1q5dEPXAAGUiU7NbXD/iAO/gb4NfTTwQxFvyf8EQn4vkPEsLW4+QaRYteGjOSGP7
IgkotcWysAq+av5y1NyofuoabC4Z5UPeZa8P1E98T7Ev+48f/ia5ht3QAmDuGAD3zlw1eMReIn0g
Av6K5kA1nEQTgI+JYzknsN4Y0mKIEUQVOTbRSjuI1pArCQb0lb+nzLki8cG8bNW5OZsuOl8/sv+o
2IACgbnOney8Tk5qEHs+rekSmJs5S7+Cp40MYRI59N9wzDpBhHtWfCHPFfZD88oMGxwmN/VLDxst
qvrAzfRZF9A7/F1Bir0HfVehtvLxDHoOq0QyHnYnzUJnSBfBPBtaQXkYa4aCZUGvqXyKr4NTYkef
iSAVxLgNNp97xpQNsB79mRWz4xJArWs2ldNanP7iWeto3hN/y+M2fl+T8ZpNKnjRXxvnmCVonULx
/tlKjSqbPwVoUVvrYmFIJmfl4UoI8kubaKyTcwqLR5GlKLTiayXlVpU4iFC34+o+SiPVYONI9Ryo
SpymdfSlB4NFW8Vyb0obgUfDrSBXa0yCeURqPn/hc8eLl0+p+GZu1+MUfM7d5dIci2d0PSoo1O0Q
a/yGofuLceog7qkxvBF62NYT+SCDCVJY42jO2PlOuJZxhGZDyeQM43qCbEBfFmV8XWy4ms8gJJ42
cfvZPvwx+LFI2lsH8pHzz9cDjf2CwXH7SctlE865UPfCLC6hxiP/AcJHjtHzHORMlyQkKvZjQtCs
P520H6KvIVGxUZ+PHCwEpVOaY8rNRuhzFTV4OT3uOsr+3T8n+n1Iz62IvrxsrTqTDqTsDb3TFstV
+uDWpU2orVl2QBsDMlf7cbWNIGz4jvr2l74U0whul+PP96X3xLI3vRdpZA9JAemoNziJFd8pN98o
IcLz+ninBJwALkB0mL5LCXhq9to5OJ/Z7tELufFQM08NiUL5gWCIQ/ADshKzLOrIKViE0vDkGDPv
QTktIyRHXiDRB48rJ65gdeIWA1+Mfj9f1pk8ZQoDM44PKecMbM3O9DYUdeAkEJNXwyvs/wzK0Lc4
5zV49wjzwL22l0yCyieJYpv30+fwYMqMdtKdLkjlquA3ITO/LZLjUUehK2k9/acForzyQUJo6D89
e0wQjxYHpcxsYYvEHc+DmpPDU6qTFPQdfWGxQrjdjAntJRPHjYqmw4kkGOavdNg7/m9qmgDP7C+j
oZj8wmeHOXCI2UZpU4a1ESAz9UEfVy9yPXuYvM0MmLNa+nUxRL2jZ0zoOEr4pyz0iENvPXQ22Ouw
WRpIlf9uNTiZRTpC1O+ui5IuzLufNQ7eQ+ekfQo8osQfFGxIRgUJM3mWtSEx1Cp88DIuXo5XhXYa
tbek16IixXlxedplHFXqyFRzQQOkx/gS/WCCFpyXn1wU5TMzT2uKkzcoYeZOex7APiRfwsqV4n5g
/yPJWYnJlsoM29b1Ei/+UsimUv0tuTHcx1d0iEEsCNkaABu3sc49ycvXhyLewKIUUDJxOAG26+XI
Y9lE9DlcxuFODDkaXxY5sSaNEGZgmP8Ic9s+9cB2o6iAKQQR+d7I0gfTML0mPbQ0dTSNGXzp4NAu
ZLYO11BtMkl22rUZP6XK/fM2v92HarLhjwJzYwbU8E84D54qStnB8xbEmCZQF4DfS6a+y0POwCAF
Gh9dppQIulkyK7zwAREKWLiLFhIMMCMqMbPNYFnURb8IjMWEYNb7IfDQSjJpK9Htz7/5ZbSf3md4
2VISCEZE5ckej5unlxUXgKBgq1oyxBobDlojyPM7Qqs5i+vGDBOJqu37ngw8o+O7zHmyegqHd0MW
lD9O3YxTweDdwAmHhTtqjNwzAnIXuw2xqW/qLlFaQWZsqPTzqwmBS3Q65zmdzXex1Yzw01wOT3gJ
nWPhCKgjwF8RfNnfO08tjzsl/e5bWJ/ZKsO4ju8DAxYkLvHkCM7pTK+5koWydYEMk6MsEbxy84Go
vFaxac1DeLk09CDWYs9b86DkhqKGczKcVaIBgSIAJVrFb3i6FT9wNUN++vpxF+rUQWpeYa7mkYlX
MZJ+NeHs33vnwzwg33M1fOZFEnrQ184nS1QCBZuX7folCn7ayjpZ3gyDwAxjKaNCTZuxpz8ia5TQ
Kff+tYp3IFcuB+sJj793yezbfA2H3QL507xVq8OMxDDMApt51CmDEjTvsSYO1Kt63aW9xFNEn4LT
S1OQyN8E42upyJtTq+PY5rh3oGiJiRYhUchPNZvyBxY2tbEmWpZ7c5FVO9jdjyASGN0jPeWMW5bO
s8wCLhdtBPTEf4Y8my6rZVqM1LRkbTT2JuhaI3wX9icbIWYlJL4lek5UBGW/WylIN35sObhZ2GnZ
Xf+4J0qj9ZHB4/Nw54OFv82Q7lo5+B6M5Zu++ywcTckrVqexRVuWgD/i/WNY8lg1cqbpARzOLWFN
ojHC7ppw3x+fWSHYnWNZnEmeGikJEQFuk7HCR2qydb9nvtROCArdtSewVBKspo7qpRpUPv9Ra38M
r3kW+d0LZ84J4uMzrz6s+L/JD7WmuFZOCC+FbHL24xaJ01zxGGT9qTLTn3uRuQYwflA8QGc1WBdU
cez6Q7hvfWq7ukuAACi6y2K5+pF+WH8qOUgohosRy+qQQ2XhxEUs7MKSaqHZoX6ycLWM4LHtp8pE
YDZmn6+jc9GwohFALJ55DzKCY79c+CGk/spPVtggdYKyTQ84CUjt9Gf+mu3pOb/CtXKHnhwxAnK4
p642y8hz2vxKlfD2pZekgQ6qW1fArcBDp+caqCpi/UovO3S+xFtz4rMa+hD58b29AlTqsTnBaObo
RQEbM3CXNFC/staQ6Q0fwLwhDQcjKrqz7otB1Yhz5lnMkEWXJmZd8E4x8jw8gPg0ZrMbUQIu9sTw
jR1Pd/0JFE4MugBU9bjcjV7JKJJK0ioJC8my8nmbObCBaglQ9Bf8m0RAIJCxUNXWNoszWCa4Ivgc
SnGfUkU/D3wvjXl0NBqd0jDiw6AtkteaOcpLolBzn9yzsubJSxZAsj6XZ570WIA6KuRabTliqQ6e
QUGAm9cbi9t2jWwgCR37mVq6DstOct5Ygj4ZckAVayElCo2DoOeu2dU52atGdlCyKXebvq+xNCVD
rMbULvgKj5XxpeQZLM8fjlOIahbBgBX4ZmTUlyZ6SGueELOBVl6OXG+UmliTdxYoSXZhnpHZa/Qz
qwuq6JAwj7l8RcCCWpnHkezqER6UXKHzt905aW2DVigcMeSCmCssSV4YLmzNj1NxHZcWGx0If4bk
+JJgd01gqppjs2DwVPirx4/4RZbVjC9yVYibOMg+DwG0k8ZBvnwm4aQzhSM/WDa1J/drbx6nZH0P
Mv2pO5P7c+BZdTBX4JL+qYPGarhW//dJaIs8rDO4xLgMrkSxWUnYZLIr4tkcNrNkkOuHGF9T9dTP
ppO4f54k/KEuueKt3NzXj35QWbh8yCfBelrNUB36itZ899KWhJ6mYxGV56y2eq4BYGtzhqZP+91A
MVpb738J271tnLu6CmEVVPl0JK6pYPjvhA0ZZ9kBONhHaVeYj7lI7TsB9pttUJEk5/sY3coY02bB
8lXWlXrdXOGsh39tJJ1ssrF6OK2AFVf7sAYnJo2V5l1DIa0DJp558Ry9afsnBZ0tTmesXNTv4LZi
IT2NAqzewTN/jb4K+ri+CkY3trG/V+v7Uz7puDRYSM+NhEMGmX6/kEbM3mVePFsJMzo5yE4A3FDr
7+c2WlsVybNpR/Kg0tB/4AJJKWHk3GMdcVZyd/nTsGyXxERxzeWf8S7e5LqcDInuknoInpLiG4nX
CHaxqdBz95ZjoXbsqV7X3ZTxvvd2Swe8a2eZUU0AOuCDIbRZdSWUb7Mp91APo4uvx0rJktSqg7Ns
r5J5kEagdk/dVh0IoiPpOKFMY91aIsrQGP72m/MoaO4Z9wlO/5ADSrWZKRgGJ3g2LMNu1/vusM0v
CVkFLCDpDjgL2giYX6BXYwzk2qbpGi8Gq9XYuhRCYz3rtupv9GmhxDI1UjXqiwjFgXj4qc1hysN1
NkAwZ2lfx1PH0l9dIGtVir61r4l2rYEy6U91FvMuBvN404a/z6H9P2UlFgL1dt/PLPs2EAvb1++T
hX6h3ZNEg4JHkIccz50RM79Q53LEsBUSa9NpEnGQcM4R5TXrGjU49o/ci7oueYMDDBwuIWJc4M7C
uopyj1UR189ndeC2RSs7rGO9Dcdl1ZeeRC4nuImK87EiCS0bHvIIlBanr3AzPRPEvBkqxyCsJGbh
cFh9mWsFd9xctLmO0zSnv/oz3GpYgVJH0o+na/N8u0B7i97gZ5M3fXh4dyyH6Mdy8MNNRn+ci749
Uf0701wvKfueo+eZvsqgUOg+hIeYLBiAgCqANU/HT4Q3JmMJfeZNR8OAMoJ6xKp9Oj2pSiVWk+lq
xf0M5pitOnly+e2sSrkyeaFUi7ndGZ49bGZekoq3xD4zyNbmMICmiBdiYiH6qOy/kZYl+GvS0Si4
37pLacuIjoofIIcYOROjd2tv6pshBDPYqQjeMB6bkiLWCZo+UkygxyTNfboQBDg4S53PPvbhyfPa
dJ2aYObroQL3LfJLPzOd9y/A+g8j0GHDKWHEA+WYwIycz0jYQJ0eRvhqi7sH31uk+CFATtyyuYW9
2YLJDrJgsSeBl00SCOfbfSU/2CxHj1J1FzFrAghECHmm1qlDdjCy0/2GDT+HS364NHJFM3UTtpUa
AIjEp/pUwKc0rSCpztwjzWZLYCXTc0RwYnBAftCk7VqWkTxWW84tSvoozEXUfH8+aLnBwecxdjix
tfXKMmNovj9t2amS2QvXjGQNu1y8Npic7rCud0edmPRbLrbIwzM/TCCMDnx59HpwJAiXp9j2+8Bz
D+Ip75IW64L5k/o+oWAiS8IJfBNyc+Ih76bQ/0kl/2i2Po7C5kx+eEwXNNz/7KO9zjyaxXOOPgYv
8Z5rEVU9GueIozty1G6toB7Dz0w2FfG5gzFSOup5f8Vsmp9BLXx/3JVVaNeXTVOw8CqZvqu5A6ij
lqJSuVvaKmiatQTUTgG773ZnpojCy9v+dvKxLjYIuS4MdHSLcWxItHGnqW4HUC02uevbAEr96sL6
TCA/x9/HqA4V2/AC2lqk4BCGGXoTsu99Uixn3CGmCTKN/6LZE6e4h2zCNoxVw+eoiSGhDpbLKyNG
CqSHPLbVYZ/5pSYZer+Tcl/uyF3uhZG6NsAVVC1zYoOc3friruqMdPHnHDrR6BNMZ/PVunMFlpJH
aEJ1eGmQoZg2DzH9X/gMneSeiC2Bgf4I0scxWgjOaXt3eSveo/ncXM+yWsAjWcDpHAbFiber8Giq
tMz9sN1ypwoRK49UOarqxCYOfH9DnWld0/NC1WWj3OSnxsVywjjAOdsUjlo0rVS+zP+hw62K+hPh
aL1HHUH6r0JjGsiFdE7gpY6wEyhHLfYkI7Lg32xEptLUbjQiiyUMe3zUkRV0LSsNguetFbqUsVDK
LbrDoa2VMbfTTVZjsGFK4crQ2yYs2kYnNk5Pe7T2Sya67u4l8ADPcKTqgaEohrQltJY7jkHWbHK8
df+R3XGDTK2BDlBLnppQwTDphvedInmwjKC6rN9I4GMftqfqUqijW0l2xAflOCAu65ZRB73QxdKv
rklp9npI7waGB3oT/2Av7IPugtv5Qd6Rk70knvpFFRHhJGGichC30vq5/3eNx1LjGwqt/rVZY744
oYQ8nJ+HiXCfeCCdgCxP12kq4iaTAftLmv7XP+lAGAeqJR1HkxRJa7QmCPvcK8XImnLPSY6NK2No
+XhJ5b7EFVdS/Xj68ORttEoXSmQm2imtRLRiAOXqek/B12w3UDLYjntKPKcm56yld3ZP0/rhIyFr
LyHiPOjqjc4Pcupy2jpNE9wFlrvUxKR6sQCPBz9VFyRqrzJBla0GANl/VBNDn2ZPTFUguoLXOY7g
rGqZUCsztMu2lIFMtZFrVxiH38VbMQBHJTwrUEqrvjnAbBcp9cSX7nZwg3iRDWfrV1km5+0fyLWX
AEhHqJHFScxdrz5S6JyyyN9m/Qj3n/BIELC3E7zNqtM2xcXkqLmwrxKKQla2g8GO6ezcPdD6RDGh
GmadpYUlIUhly/3sXVgswlelwxi9xv/hJ9bzk2xlVCqpJmJRR5iY90/S+xozAsfduBwdJWwFwGl+
xyev/pQqKL8hnAE7VtRoBZDfpSdQlm9tgWdhhG/utBps4EOjz1WphMK8MtoeoxZAKXge/QO6WbKW
HxdGENLUDB6y+q1C4s5gtznr3oswYJqBQSxCpYxqkHo6ge/EVGG6bV6oPXQdP65qoc1cwM4/kToZ
ufGksvK9Q8AFIW/30I5bzCgyw0/kVeoLr9um8H5LqdCPt/752guuaL4ElLGI4sqHwFlJmMK2VXyW
NXbV+PCJFomng+FyFXqNEI7xYetCAq8qC/3NU3n2B95lpWoSXf1xkaFGskLdOMrSGzSigmSgXqlf
8cMBaU3rxaCh6/7LfZg6DuyLOREy8lds4b/M2zMvxICDxbAju6gIsoYs4pQ2LpSG+h/L+db1HcEQ
V86QHvVSezkTW0q93/eYIVGeCzt//C37k8hc1V2xtwzEoFkTlJJrbHYzwDi3VnawCzaoT99rnsQs
MPNhCiO4LXiwfOEhY7EelZS9D7lV9N1BPCiNlpWDYe3qy10NJb+gkktCeaRuK9s35QKAhbqYGw6B
4z6PgSCOfOGAT+Cs4pXqw/6jiJDNZUQ6Dhvt4KTBfvN1ZgSkZe1njspzcQjP0Cd2YQ9F1CpQ3RMP
zvMYrjd/fJhhHo/EaOrey1rvea+Ho4FgCeaQC4r+Abp0Blb6jOku8gg2eD0PeSgCDEL6LaI+uXiQ
srsLZLpkd2lqzeJlIxd1qiu+IMGeFRQp60aUdlDIVyX4UQV2Awjb+C423wb3lncpcZ5uGv6RWvrI
5pmE1pWc9ZcC/MxzNM82Ujb/7JDmYPUAeeyHFmZ2VJDKKg1sb8ON6zo4UxNX8qMNAfJ+VDxWPDf2
cZLIf33bk4YgsXf9Gf+qFCsFNAP+OW/rtMxtI6JCMsHYaVtxXHSlE/ExmQnoe+5rpcpqIQMoOWkd
5J96o0yTwEgfhTiuy58v+QXSu+gtFUDajyDumvcqXKEUrZN69zkYhUCbP5E60R1hzvhnOoNmz9oh
q6HsLchQ2vZrbSXN2MAiQlSrE5PHhuwL48QyKV2gmQYQG4kUKqgsoY4vmM+6KeB+iicBnyuzU7Vs
Itz4gh7lR9qahguQQnu4TQ//HNT/mY5fJZCGBRyZ8Go0FuRO0KkcC6JAMuHnwbzQtw7oWRGrR25e
WIGasz8wVdsKtVykvuOgtGMwLqJKHPMF3wckRfukxR3PrrLeUA+PYHtgnmWJ8BF31PXKQk6IA2H8
gGi74dhJYscquQm+SiXciRNSQUgJE5KIJz/6XhZHmvPkn/ZLH7gkUlqdJbyQ+10Bcg8aREJCH5il
XnKsL9OxtwjoiMW/Ji/F0XnsIYayZ1oQjBBwlC0+GQ03QxgkVZhsjmjfrkHY2l4zRNLQRA+/SQIF
S3RiUdhpIDf9mfepZ29375wbgAt6PtHKEHO5hfGsmNUAC+x/FPwLuLEbHb3VeXRqq4Wrco3ezj/e
BlTG5pn2lwCbYdSb5JAiBp7Zr1hXEMR6H4A04G2wK9un9B6aLhZwTGUelS8v2izF/hYILcJOZbHW
I5oZIRhnxtBq7MGckU5hQaRSBFHsKu+TCtq0/3wDH6ULyr9i82wmaEGcAdb0+bOdIPb1LkZf+EYy
azCfRnBBiKHQ37hORYWFFpk0p98TZmSnHIhq2AeqkXRlzb2UNcdavQF/3mIiVYIAQjTNBhSwKtRt
Umh+HAq6WGhb2zVZAiZVxyLv8Molx6IoyWoJJ/1IVYZDslPuJG0IncNVMw3w5YG9BiSalMPtU3/U
A72RBreaLFXlEuRQ96lBVlaDqlntOij1PulCKJJY79zVgLabcIL2gOJpVSnbEzrmubsJhnUhmMd1
WD7mct+BPlTw1xrTnGpvzl5XNkxqqpHb5AiCmJf/9HtgwgkxgTV3yzY6RM0rionTgq4AH4HyeAM3
InE6o7gjHlknq5xJWa1UhcboLsyFY8U6bmZWxBMlgkbaeLAxyyu3DMsi5Xdvlwml26NlO93J2+MZ
Ot4QC2Ovmyl38B3+iXcQYKz7+QtwUvXxvtkC954+OLZH+KnrToT6tIgnrUHhgCh+tBTJJyb1LzAQ
+VwZ2+beqWJbXxb1wDbAchc3ySw5xQw5VwiD1F+d0Sskj+soxtNuRxFnlTqV2XMzn3w+UZFaBHBG
8Gm7Gbnd43UXNuOlUoSLNCxaHZp8v34sCQQ7zQHlQdB+/JiVaPZsK63/cDpnkugJYz6IbY7obSy6
dbCzd5CFPacG/4zi6EzlDbZ4rnV36wVKWuyWINUcYv+Rs1VURT/O16TcidIkDurREuQwJ+ovCxqj
cT2C3pzYPw7kQjHlMX7WTxJ35wfmtQpNnSxA7Gs6//QbFIVD34et1SHGM/Xgm2PVG1VkAxNnIwkl
jSu0nrpMG0yPgP7VpCdkWauFI0X+Ta7TrH267tXTf/wC8YN+z5BtNqE0ZC424wo3oeeCpHnMz1KM
II+ZqjzgKs+S7s8BqX+PCoBkwk66TQLGB7JpfQidbtUHMWzoizXToKViaXBrfDuRxgn0K3oDWj23
paZJHhMgFOnVuCLbj81jFCD1sgWRJiwnpfp+JOx4rl8/UJDRkEhhcIidi3L8UScdfyg6imiyW88T
gcHO9VzUHTiir/uCcoBVLKQiUD76Z5jN2QzOvZWMk8lr6Ok757DK3MvdoLa3bpKmOp5SM4xDvn51
+clGhc8RfTebDTIqBohHPStOqB4LbctWqJ3Zp2ZTEOy7nGmk8dbNvLgXmIM9SFfBK9sWkC4CP/Yk
s4ZHnjC44Gg0w0XknlOpxByGK01dKklBj0avnvN3p50BNNXYrEjOc6V+ThGqO8dt7PQarNTwg+LL
bXH65gb2BsebBQMtNvee+RI4VcKzPAiYXoM6UlHzX+hzJXQRVIp8Oudbs5OfaLAJVISgiPsM4zRU
3ECWtqb/YpHkaW4pnTfabNDbW+gp0tf4rUZ7j/84KYOEkcnwMOH4gbA9a/V1+nx+P5KeoSYlZf5v
o2Mz386UMh+nSGOp6YENYq5/YU6PP2NKuFvF4Q61TTlkO3+ZUaqC70oUjNle5FB73RxGwk0K8pao
OX5ovrQM8l2u6GqEECHCSVyplz6lJ4J8oSk/7Qvc2jhEmvFDPvGCCBnZH6ycXVxqvHCihacmiNen
x+fikQ7gNovecstI7lQ66wrtj8d2MkbZpmGN9rxH9JKuqqTImgtiamWfuUxeYVasfmyuEvRuhtFT
liN3qgezdSOI4hkiwok2Z+2PktFLZzYt7x8UV02eStQAwD36Z7mb39Uh0M1nUVojkVvOjl4Ei+vF
HMSMTwTdXI38iJjPXgoxpyYSgIsRowMcQkilCrdYPeKQo7IEE878Ufy8uZ+LDlqZGyXImtjiyLUg
U3dzELYiv4N9ppoE1aGUa6UVfmOmqS4iTZtfkyONEHCqLOc/addZ7CEWwkv/jzd7Vu4wMGotfRb+
HckBnLjk6SjatkgRBi9cq5H9kkpDcTATaRJ7+5hUkE2LSoRbXIHtkR+qn1n1o+ZZUe+jwvmyLH3y
D+U/hbuY1FHlw5S3Y1XEET1nTbfGnCTJ28sBhPRQV3eELoBmyClX/OB4W6s/auz5CQPrG7vXOHau
E+ABhCNqwdR8n7GWx/HOQeHFdPEFFpVecneT/7UBLV3zNFortDgSBMJqKCobAwFRzDnfsK8qvAEJ
Stmlg69/ncD3Jkn3Om20KhEVH3z3jlaCBj3nGvIuayqyqUtGtTKBZGqNRDc/peKzX5/rTDSoqd/A
skXsYVW1F6UtRNoSqRm9k2aZeRNGSenSZaYRt1R1AYXLUHe6WPZv0PeG1Vruui+7MegHCDVdcOhU
WRooWXRrkbXIqK2828aGsgD8mOitejWxYz3VvOmQaiXWMHQ87gs+WiyvDVaa1iBbiJidrwdAm27d
+zqIKUG7n77C6QLFvZ5RNpwWa5/MevCIg5L6lX8g0xqTnKysmukkkmC35i3gx2sFINzFO1H632XK
s+N0mSi9+b1xsccBHNk7Tad8VNKF/fzV2h1tZzN9CbXs0g73ZAWH0YxTy8JAh4nt6lBrlqyHowtj
b+IjA4ViPHtoT5wr3hIBpovJzVFlt9wYU2XioQl80fxcHVNKL/M0M9BDpbKBluG5W+x5Mm5WzSWS
PigHsCcqrAbR9MVuRRbY+P8qFjr3koj2TVJDXTuiX0igJkrhq3LAQPR8TeFx9S7f3AUiVtkgfBBG
eiH5AN6qGXygXq0a+OPxfClaSKJhuDW0tTsJasH57tYxyiuiVOqvKSrJFhu3hZRl08rWOyxV1JfP
3SdY452hDpSBThQXc2sO8fUJvHsXMyRVMJpMgvCRReE2GjBY6TfhyY9kQRNxbMgXx78XBqoSEA3F
7/bAlJ1DLrnFOAtPVaWPgzYu76ICS9+k8o61t870hCZHfvMffL9jwItfEDFDzvz1S+Y2jk2x6FTI
0xPIYCILfL/Lo/4a1qhN/PfFnxL0IeHTtDccf5He/ZiALYXRcuguGP8FRy2coxzpIgGbAa+4n2m+
8AkQkno/JaZP/52YcbGQGxaB8hNWyJIzIDuklm9JnSUF8zFJk8lpP0L7r2ZO77e1EkC4F5ffxY6F
W5Vrj0RKFaqfJpNfegwYEHg1JhYfBAUl6ehq1omgk4+teqxz6JtbFBoR0ZUJVccLLWFeDE8ajaZI
H3xEAPISiT2t2fbPZR6l7KH0XbYxbu6/wsCPEP3K6ZN0gx57oSsy8Bwzd73iZL/1nePLGXhN6hm/
w4CMo+QfygyHaxtU2h5UM5KX8/HBM/dn2Hbj5QZiMenDm0WxWnl7DlREtDajhxMSMdfQWcQdsGni
eCeaUtueCE3OqQ7Bsblsiydt2iuf1KSp/6j0KfcTt3X4wMXnf/2i8jxS8in4FiL+MndwAPrYWTq5
YvW5SWRAN1ixcpGCm9wuHp0ShJ00UlTY6qHBo4FAms+SgIK7gMuzBtYjqW9tAVzgyvv5gflkksfC
h7le4X9YOKEuEGKRKVBKn8w1rT9lGlZ+V/UzUHYmXOjazywXcKU8zYICJZK12O8XtKeiZ6Fgfkky
ZZCzVBAd8uC9gvGJ01qK4uJepJAqphC13df9InlyFWRIW8CMPVLyOlSkXJnygSRji4mE1MN++fkE
rZt87NwswSU6RAlDUwDa8vxft5GXrFLde8jzTPV3C4Pbt/vOsmF0k8Ik4anJAIg4hUkfUwWqj3Qv
uZGalgbEe180/2EYaIyBHKN7th9w2nr/Pctwc5XQAWuFMyny8+ZREy/8NofPeE7XLla2UXeqHVir
oeLbdOdEVjot0o0GMMqMYse6iHLcp/z9uZ2lPLvC3/Zg1oZFzp7ckKAnLfMAQq1j4WQEKPNdEPdj
PxJFiB06Kpvk43vuO1qHr8XSbhvTcyMH/Ra5+85Oy07wWlWK0yQPTbFWLL2wyHGe6I5TRo2CGyYI
czrTRV7kWaNTu6HTrbZ0wPCWpzry4e7H2OUsD6MBZC18E1HRnhVlm5YUqJY6ClD/9S+5HJzGkvjb
kheIWwuelGvF8wZNJu5NJxLozJeM8J1w3NB27gSvgtXOjnsN7H0OdbsC2Bk9e65w7FXHeTeOCLkp
8IqpNEN1E+vyvpKe+9J37cpj2PkRyzTBCrHBre15nvr/8VfGLrViB89qS+cuF3kTl1cWRZsV1AyL
Z2sjVoYbFaJ4BLdzxyLZhlYNrF+tUYb80taeui9YTSODIe9175Q9v6NnxdYQP4q7yY4HsvpWx0rk
7huw78WStpvGOUHmsJnZGf0rAWZlmHufTGtUa4fLahz+wGP4mo93nGektOSkpWG2Se7Sb7z/rUwo
BG2WQFY7AR6SlmfFZFkTnpIACAT3GIYhL0OKjkHG1HYY83DuAdwHO6VLii0NIkyVpFDmu7A3Tpiz
CT9LjePydoTRX7fYVfWREZexhAkVb/RzPtIxi5TEs51QuInNalfCePWpSaiAWw08/HjRhnuuv6rk
VjKGw6vevsJb+83LFWrf2TrQ6Q2n+XHQEAL28/STFl+OwarZARlV3oBOXkz9DRNVsyfN0DtBKgoN
f/Hcha4Xw4sliDbYUbos6wL1TtOLv5ft0lg2tu0KgyjH5RLEnWfX5vPhYikZI+1oTPzHcF2zwZn2
iMHXmNFJYpnvDMA38YQjwKMPwCTP6TTHTd9j8pV3a+pq80TYYdlfgrHbZJOinzD4D9HO7qr+zlUp
KbKTMAASrSEsNzCaxf1Cvs+hDszC42KCaHjkkzdW50b7QQuvmwxS37Y20DthaqMmOMklS+TKpyER
daljNPpWkRvlVXYwrFhuhDieJ0JlQaLdRK3P2G0B0/iKmQvFraKz+j6/U5nT/BSsovs83xrt0gxJ
MiJQvHpBWzq2Ve/vwGgcVc9V8MBLKxCMM1RPxyR+tj+qMY5oGoy0hPNac8WDsGxGFmXOf0btzo9K
1FyJU2EN+aUC0ruWrqeIbJGfSMWRi2gdmNIbbZ954GtkDzJypdxsnw2l0mW7uIqySa8hPihthhp8
x94jvKHzQMhr55sFQAjPKH3ql3BNU07hOtS/44sBOMsrp703AwSsYMkYqrPub0GhxgoV0NW/Ek9I
riU5qWhn9gb0oev7XtIbJ1LujJcEb/DEn2NisDzRjzrLXEQ0b6QrBc3bBQTabigRuBc3vzQemd5+
HssTnq0e90FNwYA4VSCs64ffFKS0Wnfpeqt4Q4yCrXqEzGVnHQrZh/fz92MJI/wOugVrV0M0snzf
iBmxD/EmPtbD3t5mYgrUPmsZuV7RX2nr3VsleXAFIqK2O4Xr3WvtOsjELoUlpeQcFBkm4y/v23T0
vf7hfV0vV5EBvcoaLMrlLppkQ7jQ161SVtRs7u3V7ZSftGhC5QZ+nw7Y1l1aJjW+yxl6ADgGSvrd
D6HsiP/T3/QfrqXBYpybmB2Hb0eGvJP5jtwfdM4SibM7adUYh4uIhchNcUH2rmMZX506yfGD59Ud
sJS+hmQ/nadMnF8bDUF/cNVjJtDFXu75S7V+WG4c+oWh4inr3OlhuHNbYn/5ANp7nRgdgVCZ+TBW
TDDLDyAIQD3gPgH2hUQ7J11fsryhsW3kJeT5A9y21LK8gw+9v+g3B2zQGjAUv58ZPM4TcMTByRxd
DvllYXKk0s1MEYUbkVntH0NPJZJfDy5Sm1OOsLXGc67n3kBZpp2DHlwglihILL2WQQcCLeQFruj6
uLYzq6HY1zce1s3S+LGKhJvhKytR33++f++U4eBS5wvOgj/scASVZwpCuLokzr6R4k8xVo/lLJP0
mqUBSCSfiKI2eHRbq707yBp7xWm3HJDu3ZUrrS0XO74z3Cj521LE5nJOraaly+j2OaAzqMoUUpCd
ZnWzE+UskpyEZwRGnj19cXtKUFJDV2fv3Jn+oR7l2YUCQ8ed4+5eMzqQT6n3ypz06cbbSJmKJY7h
NReEQ8JgAYeue72KVC0tHGMNGpg30yqsVQ9xZ2Ru45bjdW+6y6VFEy8xo533FXnL/zAyS4/3JVFl
NPvf1ZPmrchDODyn+yTWTB8FlxCqoK6/l86pvzw1qibDLLwArKRwP1ouCh/KFuw5wcBd91sqM8Nh
Xf35Oh4KoBgkQiyrvzRE6WsefUe8yM703H+ZuTsVDk6wiB8cr9bjFvPYgGdv/3Yx2xrjBqo48Nr8
O0C6yuVNHlQXS3HQUpyjYV5JijCTtwARsuveTx0O/rI9L7JJ86z5WHRjEQZKljdCodQffrh9L6SQ
aymSEtDKleVmhWBkAz/7yf3oqP90E6JoS4gOp+3TQwhyq2yGDwoUBZUOZCW1BjdThQg6u7aOtP/X
GvpryYkanqGD073ITcSCexrgUB90T8gal4V/0CsdFqdaI6Y4qBw8PZfY7Ffd9LAqPr4JAUY87fCf
ABxw6MeeF+HGozPF0ZRENsMPBK6yRpggrtpwun498QqNkmMrTlyxxjhVWoVITft8V/0F2YeeIkv+
7VBOoedmxVtgYvBWyPd8sQdQ23WlqzQQrzSBneMOvKWnlPz1chFWhYpFD5CEtzt/wICCOkFx8lfk
9jbN44LYbBDEvh41vg3ErGsXI8v1x8VXZlc2jJmr+/cNOdeFEW0csofnJblLdDo/twHmfxyHaf9/
V0RwHrN50QXRI+/M34Aa74Ju5ZqmVubv4rzFJ/eITdDJaNeWy3K3o8cDhyCwhcD/tMgHpF3PVawD
6wTn11zenpsSDo9+JKwPuAcxntiSKWf60xZBwRweoqcRap3V+5LVv483IVvISCLY7NYg/vJ/OXdW
8tzj+pGxnW9vwwy9/aUVvJPvsRGiwNHTkkPrrJE7WqaqVcoI/JerMGe3Xow1qbWhnPRAHz2NH3aD
WSM8izIpF4WO/ckiAktKi/i3mD40GH0eBEVrVQ3O7y4Jk7wxcmwOogXOlGOhrMwGBE2tdq3UQTVU
qJEtdTs/obgD9Zh82VVzmiPFqGbaUCE8IZRenbklr3kpAGuMPbzWhgL8IbzkJWrORIhB03B2UlOJ
Mza7eDcuU0pN2cHZT3L+CEZgvxt2ycu/U0jjo33ZI4LdTLTap1TssMSA8HvuLttZ7+2Qh0FwdNJl
F8cC21zCKaHyIcx6WFj8obSxvtzmoFwZYwriTJ0y9fS9tLE/wUuRq8qVnfu8J1aT5pAnVqq3AgQ5
laAOpkzTkM4OuR03ZD9fMIPMG02YihHyYpoIAVK5m2yz5Xh0GHj0vTqh4TH4OMqB9yhv5Jn7zhRO
+9FBeqvMvwqXjjsMGKIHTTT7ZmCwO2QeReER55GUD+fTUar0zAkMKNJ/w6Q3UfYWGRWcevR7ne/h
HRF8+DwMneBUrMyfcxJJ3d8Prez/uoyZ84mtZ36IS08EdbfHzvChG4fQ8P2Le4jtXhZwvjAJMkSk
HCn28c/dbm2sw0PFG4YEWncf01w/RVOforFKqOadKa1kdn3KlgcN+yzJTzr3z6WrZup10HN7hJse
US1//XFGJ/j5EfZH2NtbmV7TKqwzy6bBA/etj62vEqEBE/tq2uuwklpO7NPhKaqs2SOIznPI9QN7
/zysiI2FLY+mmZJ7I/6L4CxNj3ppDqcbAwVdCNbHo1pe11VarI50ghIVjr+Oct5E5JOfLJpmCX/5
Pc+bjfAdKFeVui4r7ndBtevKjm8wXgI02w3gJALI+aPIYDIA57QuahSRS0MnFs4U4NsbQZR/2JtA
553jKa9It8W3aD/W3L4zJggMM4QLBQulfxBuQoNi6vjCaUMMPkm+xn+GG4BQM64hXVScqNsPc7X+
pain3HqSqqCgmYlzeth7zYQfpQfJHsNIVPiO4oK+cNpZWKXDPbNZK/T3SHCPRoAkmDIbE9q4HXLM
syv7E1Xx/KptHuLs1cPZTqnI7YcmlUIgfj2l1T7rDcmIlV/2BvTezryKPqn4YcysysloxuuejxQb
Rktk8eOt6UMqO2spEVt1PmeB1kb4lxDO3gbitvJHO/k2wRfxTbTxnujiDeJQNLvL2EvlFLc9YbKF
8OtX8HGaPFqtIeJeGt3EKjN6S4nQUVk9EnLeb6woefS19aU6zTfv8AGYN4T1kj5z0mbRU6Zevu0M
LNsCrabqa2zBDxvSGh5+Fa/LEPqEVpwjC7Oe+rRCphBBjOY38fVWJF6i365yr0bNQKYbaYpgz5wx
fVrrxbwoO8pW/B98phC8D6kEMgrr42dH4uWWQD9Ca3HrxmArsd4kgTvWr++VN+FfB/9aXPo4UVhS
t3i6xJUAF5kRUmMjDC0oBo18n3n8
`protect end_protected

