

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jKLNR6CFLXNaFIX4EgFderMxPnKvpk4F9e4rB0Z3eM53MFOGJNJgkVTyQHI3/mIWOAReZVwoVOMa
CdAhgWGvBg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9g8iGOMco4oFYFI4TkAP1q7tC6YdaKcKnkZE7b8B1VOvr1zofUKAItPH7rdgXy1xJT5veYU9CMB
1a6xkY/7hrMk2un8LzBXxNY3CU5Bicpo5xvFJFwxXUw2rsZfzzw96pA+9XCQOKRH4TLd3b9RF6St
0jOdYl4JHV8zrfKdmxY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T9dmjYx2RI0RbX6wqo4nWU0ad1An+UnLDs5SJii98PTuke7wRIDUcgwzVXGZhnqgRDMGrxGdV3bv
2TG3EcxZKQwTVnAC6QQoZX/EtMHghnA62m/5NpXmoLwh5qm/MLJ1GcevcOyCUPonSVz0GOgxnvwj
ooQgeh9D1jd4jba778m7tqjzyqrMu2wlx/9bVUabKnRucVtEhLrCSutcfwtKRjcjEslE32+ANJJO
LU1E9xHWQKY0Ykt2thHoAW/gEGE3TgPPSeS1uMgC9gpn3KeR1GWNFmz/5i6v7Pure2Hjx7n/xHnI
reb33XFnLAOOS5csVRvU6rhvZeRoqLN9Ju5zBw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z4MAcGwOirs8ueHe0/LAJt93fwBMCERy9UlyN0pxTk9Tu06Hakd4P9cZvnfzA7zREYXMIBu2NDPA
+322PzRY4McOROTi9fUMbDa3sq4QlE99HePrmhLC9MCN16iXhbU+HBEFNxdCuVK/qDkcEHSOzIkz
ISv7GfjVXM9ytGOZjadyXWLpl+dtetGHtMec8w91cjipLXbo2ywr8DccFy2Q+uIfn9whyWTv3WTK
w8NeftqkhVPZqMJIv942kdyaigmw+FAOB+eg4fWaELYnDgvofFaanVzUBmReOY7/b3LQoUhotNip
TF4puoXTeoGR0ir2Fw1i4DrX8pQhZYrHf0g2Fw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RhMVl/dQLgd6Em3cvXWswCuyQybcYHVY6fBYkTB+0qwPgxUd1H6xUy5MSLur1rc0+xMO7DV0gkc9
m7J2qnyE4PeY648BXoQQvdkIDs3cDfJUIMzBSJRhAzANt/GvnCfPAPUqQ+RK/y3xKJwLsMukWXHR
t1HX/5OpB6TQZHZYE4vz2lTGPGbVIW3QDoyrjz61tA/jsHUVGJvZ47VdBmfldxPqiY+Vh9e3dl75
JmttiC9La0yOzL+SocwWzDn/QZbcRHMsTtLWlhxlY2wXUCss3GHmb0o9kugY6zDzV+5nG9yCW628
du+GA9eci/G4jwl4JXZ6p/WPZm5Kh58Sk5SgqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z6wIEFjRiUpcYIEu93tUzSRYb0cut/OLoYvuGPmJyBKSi2zPwapeByA928Z27t6xeV5W3znd08OP
jgjBqsSWHmyKGPK5eXde25Rc7IZneNvK+sw4HV/jPYtO1qybQvKRnWu8hrBhMhyAA1aL1U4QhZ0j
OVNZp1DTIxg4hiigHOc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M6YZEFH9Zpi1+cHBSrOstRid3w06pA53vGHrYgHzFGeKeyyHqjgt7TSqiheP5aW8KTNRQvg6odJR
cQXh8v30NMYu/jZmXni3nFsFUTUEXNB/ePMil1PPUrf9TNxaYXBqeX3zB6GdK72zXdmYAQQJsXm3
TD92LB1fEOaj3R0/tHYpufRdGd9ixd+Chdi8l5QOJjm+yeF3y5TfCTs0lUF+EsV39HM15hn/yqbA
gT+ibQT1xr8NpGHcWrdEkzmjH4Sn+dW0cT9kU4XilATPF50SYk2ecvCzISKLFkmNR9pfut/nGA+t
DPxZ51VLTruJmPjK9LFCbh2X38O5lo+z5+P8tA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KfvJFdvhmWTKbQ5Jxri/BeSIQO81bjo+x9EfkeRcMGW0X6ByjZDkAzxfNMlSiensyevMJMtYPImZ
QLedqWGrPYexifiq6cCXFqk8Ltq9l5wruSZyV43D0ysRcxj4KEmXC/8PpzjDp5HlvFJFOJ+D3g6t
NM7RYRIRIXaF8CskZw0jsmkaV1T83Anz/mZ/uZ2VBOchUsPeuvhUsVWM+cLnpjlbkKWXTtBltE9K
o4i/EdrpFyh9UMZS+xmXkJ+At1Ky5wvIPoNFGMpkkGQACazCdVYLc9yp6bpOYlB/gizgo2+PRrAM
svam1uLoF4FsN5wTcCULaxZrksdIcF+IAZUtMA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
yLKUy8ccHHlVHDiq4V0aMQl0B2rIci6tjvLAbh3dZDYRy2BceMbBzp7B1nP7mxZ+zKWg1+SA3qZU
1YuflIuD+43Ii0Kh8QWAbTyCgF9ldpUQl8zir9K1yF84M0re0g49wWw0eZv5oY9yd/7NX3hNLuQU
1vbV6bc9Q+vzq/sN9RpxCIG0w+oa6Jb46pzzvbugFOJhwpacVspnpsgj6yYS7gE2X2bd4ig0JLvF
8f6Mc/ADSzv1WgzlLUKdghit3AMANLOaRUXklOF6ON4D8LYUNIWGACGMfBbcumapfDyEiIJdNmQJ
yeIURurw629IqWUSl03vVNOxv2n4IBXipYdEPzC9V3z3Vxn4X2olPISF0vs2nnVFeeiWL0SBC0Ui
k/0/X9i/kJGMVnEr8+A/1hd3nJrIG0zYOo8JxS8dSjZV3ONCEB51j+PpLJYEki9Mfs8SZQw83AIO
FvVC3KbDL195VL9HfGzDcsABSs5xb4fnhqpyXJV/am51yJS4mQ581FlHDJzh8WKWRmHoS95Z1COV
rxUWBBEjRdki8DAYSZCQnWhcETKeLyCMBldmGC1B5nSoMoLeFO9NSx65iAq8PuEwp70JRu0B0uAI
9Xp6QguDCysfKPnZJ8RqQLRFfjT//fO8glDL4pN436WOM0O1sxBCsSnPTHQVQ/iGDE/0oxEKEH7D
QBZz7pDCgtzCCUrWw3rkj4O9KuN+qn38MQz02e4M1++llNXUq/ax+UtM/vnZ+Wbr7xpXaNvOkm1h
H8BE5MINv12TukLbm/b2aSom2AxhZwzhiUt0qljIK6X/IPDB5QN+jY/iGadvk5ZtNw1Q5lRDIwWR
SKM3LzvgEAFBpNgLcrK9xgpn6HitBRttCs/Ua+xBQbwMVbavwELApKSmqVqdpHmFH5gzwQiIGHUZ
KxRmgYO/eeSXwpaW9TJNjfQJzi+niT3I/ulHRevxPKBPn3WAbiXO0mfI/QZNneifA30XRqgHCsgD
8oqb30XE1frVe2afGysx0SU3E9ee7gEtg1GXZ9fi992zKDEJPCcwh8/s0WdnfTrZzQ7Z7b/Gn8K7
RnA7c5OpdFGU4SEngmaaLJ2t/XqCzKyfwNbR60CxYie77gMPhPAgBiXJ8lW+ZlHxxlnJx28BMAIb
NU+Hd4auSrEuQizzM1wO/PIqY6Up/7V8OspneSAGfRgLLOLc8LV7cHl+U5qYOCd0CzrBUzfYHQkN
t2F2X4ZJe/XPMTAu3QPTtOm6/Xqxa2vN3z9MXfcjfDbyK/mHRntyQKLIetLcNfJYr/vhgopT+ksd
IC7aIl1Ta5Yhb0gwmYGwjw//FcaUONfVoY571du8kqlegRGH5TuVwLfV+pYA9Ragw0gjfGvjjfaJ
M9gqL5HlNutX0R/IwQMHLhAaeS0xsB5EJMdZRKbjO11W2sF3XLEjqGeOaYqY5untuiXVslMFsooW
xFtuidHPduWrz3VdKsbxTQ+RJMGI3TlAbVDn8YbDGRaC8n/QAVfrfjHzDSPSfQELGXDdO0QiE8K8
W6H2Puaj+z1RCHoCcG24PJDHqAHOcV3hiS4DLRspso2xaIku61UbC+6Q3IuSDHxdchXhZErzBh5C
uCYLcAahKt0PV8b6HGYnqFTnFb1oCheMX/PuUdJE8eOX2bEqvjyX06m+TojKCOluy1jwQfIV0V6y
Cw7/WqMD8ds1RVs9e8wAVWLB5WqAuVIwDN3qEylFUiXPgq3o6TRIywVZDCxKy2a0N7TX5OV1obds
b0UnVMN6jX7WJRcuOIWcnB+7aSGgsBx6nhGr0+QefIo9knJqN2J6JID6X5h3Ntxbu8XVUueHWu6P
+wvbENesfwskjJNRK+GQfnuRQMzf2lev3ijZq99vQs1qBu5Pxf9EZq5clsXmYiYsiOr5JYWescBJ
6/XIilB9u2CLkdK04Q809MHRnF99uOegYna55rtQHew9brhtvqvEQ3dDIYT+yhrm0AKRnSZW+K6m
6HQ3AJ/LDridaPt+2XqMyUNOOvLE5RzoY98t2L8v1L0EzjH8x/2Me8dh6F1/eaF4vP8mtzzh5QRC
zGhWkvvXgdH7wlDWsV1VQLi40KyHeQSNya1tRVCh51Axa9uyxTOaUSd+qux4vBNxqt3IxmDD2Ayl
FXbqA+RtPByKVQPaxm0x3gPtzL0/sbW8kVR/wXvLNKm5b64qKvR+aN2wG+5FWAVNXCRTpf2Lfo6J
lCXBW4Rm2tagVOrdfzf3fkQD6YGdIly6KMsBiAtR7ijoOMyumhGwYGwO4CLjOFxGeTpls69GPnwM
OqCtrodVBaqzJnNr3ZIUzubTqYIqHpHew4o9W+7OGmpK/D62q2tkPHUqaa+Soqym4s3qfW9o7dvp
NVN5IUog2T5JN69lc3NzmYdelOkfEvztgmjb/4OJbCILi7ldjf2uAtBe9Yu271aGdNddceWWhhyj
T1CJz7tosckJYv/bt83y9IZbO5pUC37/JaKCHFzfseZO+XzHwvo9Ua5tzaWUtZqMRahRsNH5x5rd
KVRxDeC8yFN+VL23GJaJLRdwFZDpZtn52Fho/EcqtSDMNLpnpSh3/wzTtuTeRLJpvPySz4UTuKOH
BG6r2/JNDWHn2yMU7tzYtPQfR74PilrHiIrIJC1zSH1MWCRa3c3TMERYy4BRvMO4mYvCOp417ZZ3
pha1whi9giMD2zNEM+fP/DiQFzSL5vag5gs+uLS6/Mrf5CoRpwBjc9XqpCtMJISwRxMPhujNmvj0
o9RZNgj2Z15IcWPVyl8BB6BwDgpXWLysKmN4j6evM0XCRXkiy+YEumy/aJQfiI6/zky+hXI+cZh/
Npcg7Q+9vwrmqu6q311kg31Fj+ViaIEL23dUa37JRtuZuHPN5kXKIDO3irfsv5PGiCXfhLBIMfsQ
jU0OqSKZC3esRkDyVbp2GJ6hmDPRMVRYacS03KL9uwKiGaFdM8D0pEtbro/J0LD6EhoNYfppO3dB
jw1sT9RfpMct1lUMxE0b4HMcvbr4CBxx+afNuHu+4UYxlCGsnZLESS74Mm3iYBv+WzfokhRxQRHv
riTCc8evo4uz7QNaa11ykhSY/VCVLciuIbZ7JBOGeBMpZPkaHb8EqdjYFw2EPViFvMK9MCdTyV+i
SFsZjhLOvryECHPAQGXLkPakT1SsSzS5VhxUbin4so8sP9Aiyw56MlpSaZTTBx/sKOoclRfjWbMP
V/Addxr7ZVIOr1vrPiDx6TXXxEY2ce/7xIPSRvkGmj2lwFWdJcn/sUn+14euLoHAfUAElUFhL6xY
s7mOqsy+vOfgouCb5xCBxhhYpVFjhUuW/7Q5+XnISoox9YAMHz8M2RByxe3qJ3MeGE5TTFpwFec7
pt174GRjq09pmRDqzzP6iEy0aAJccD12TvYW6rZM7yaFULI41zPk8TBmRVbCfg8x5VfLzGbPFZbu
dn+Kr+IxTB7Jv14WsQiJgs6KZvYN7++m4m05rL/L5b9eaoZKAYL7PZhvpqkvYr0Qsnxo8s1Xq/ZI
X0dQAPB4vUZzvp5W9ZfB4yV172KGkP5ubn3LZSMa8TIFLmcTzmPow/bVZCyO6uZdlcJ7Rw82umVU
9963yfajPyLvOXNHnno/oNFB2TKOvzY/RIjYEQBHTQh7yhMHUuHd9S2Yo93yBB1PlcFqaHCfAwQq
lXFHsoxpYo0wwHQIqWONFga5RlM7boWymP/kEuysbGuYf2ccUEhmxf457dolaOxO7FqbsH0RiAHX
srNink7xJkLXTgerOz2YL1ItmknXi/gdMbKyY+JoolmauSzanlxMkzcWBXCaLSWQEmzHoscNydS2
wVBaIuYpyT5qSUjEhRXsr7GGb8f5+WCEfBsy0rERirv5E1qucd1Ay+8vDHm42gWuJkIe0Hy87IYM
Kdfw6FDwN4mPMtrhgNCAApHOdrEl4A9/GH8y3Zyt1FXgwAq9rafKF7biEsnvAlhiiK0QBtBp1FuO
/rfJmL6IbNrie6WywAgRKcmY4TbffLERZgdM2VGEwrFNbqDCeGpmXPeqtRT2i0vtqM5Ao/99nU5x
HPluKAE9qKBUMtmcx6Canc9WPszhajNZCW0j92p9DeyfgjV52ucp9B3Hrf7XRYRYDc3jqM8oUz+/
I6ptlJSmalQq57JbAN7vFazMK6hEspCJcZ7JMIv1TSZBEn97wu3JX+sL8VkJjwr0qCtbAQ+cjDo9
FoxC/mRQ6bYAZ/McDaRnfPMmVSn5uThNCvpqRWiaQD0Bj0VMzmmukWclXz4t7wn9tpNvnnd0RpkL
9BssFTV1Qx9PptjPyx0zDggj8U/jq9UOtxSoqHph5qGGH5ew5mXDk2/FhsFbZ1xphSGyF16jD6XJ
cPRWAVAOyt9j/TqtBJ278sVILHsQTe7+8QMuWgSqZdhVf3IVqVTHDbLlyVlEmZwG6xFjMehhmH7Z
XdQC6QN1K7uTPSffC2DLWJDtY3nP0EDnc+7utX/OvfRpyr+nPYX83JW1BtyY2fIrzpMetpL6coRc
QGcTUf1dz8IuQ000OjvmppFfWS6gzzUL1VESL1JEbhyGTNx6/JjFehQ3YgEMn/2hRhclPYLpEgAH
Oly2iXdFPDP2sQf8S1RbJ5uf24aUWZ80ZEtOTZlBn3xDhRyVGay6cF7s3X93puA6Myhj7nFJPSHX
gMMmJG6w8ZtNs4Dv3ZPof0vUclncrXIK2z1X9FTkBxfkq0nxHvbhmBIbGeP3ZaTkU+Tn3wJ5J6Qk
34oJNgATEIRSgrhVPFfArJIxNVaiVndLx9b0mkbgj5IO0ICDqcEFgPGyxmKxmSxc1DhVqGjSISor
ucUr7G6MkhjGrkj8G5n1yz0tx4C1bO/kZTCckqycJf53e2ulJBN3XWLK73EpTQMxG0fS4StU7+4f
3REmy4n1ynbXb17ZBkgi/MStw1ppepONHz5AIXCgUSaxokL/7LHd8nDCpQ1MoP3VS0W+WNvQE6+q
7vL/cr2w7ypXxRxQuRfvQ39guTdfrhBLQMFKZV5YVjmFwQIN0a0f0axkLC6ESgNs+3/yUrTtpQ8f
sR4ooufR2jsV94/J7gDqaxb1EAkVmllx5WUCIe7PDwHkZjEU58SmH2eDnXLFcwwsfZIXe+m5+smq
7195fyDJ7cHVAaE4zmG/Dd3nG6oPBjRqtKgXAyErU3T20QIWOAYzcR1Q5cgowudoaTJkSo4or78I
KrCiERzT+dFdC+jRz+qdcGeoGXRMn4e1jdG4JTBvV/G9D7Nu8jMBnhzyNU688CgOSmtDaneN5q+l
PquA3gbkMjRWTylveouHWWYCrgfsaKDlIq571OfbJKva46BvYUvIe97LLVA9TyL/apbBA8cXRz4g
m/qRoJCg+AdyHN3pgIBoRyOfkUZ5rT2jG4i25zZu50KKOVvNsmz6eNHnX19KVf4cxAmdCmMw7xWs
eFd5mP/R6vcvHmwX6djBdgPzyUAuU2JVQvfQWg9b3F2bJPoKMImSwuc536P0d/jQxQ9MooFFKO/0
m9FmFNSbWlzU/mo1kOpVnAdbkzh4r76IxCp7Hu81I22xo07ZE0nH7YySSXtA0TfxZNPd/9Weuyjw
q+ekxDwVqo+Xg9qUoKimKRijUemq4PsGFKCfMkdgMpVo2skb29zmxp6MFkmdcA0XpaKM3aqgcqEV
a63rt1KNVKAYJx6hE2OF9L2FY7eIWGt0vz3roJJFBBRHi7WjmGr14EniMc5rBbonuS61Z5OSU5wY
cacM5jIJ13tuYCs7XlXO6tdY2xOdpgbnBoKzGry0EXGj+ZuJfII9ObfBDZ7nyIEQb9Lhkreqnhxf
C043TMxEtiOhOu/UIkehph/EhPQ2SUs4lsy9dFIhCpziYrnTO5eFk7/KttpL0FlxsM4x2UWgDYH0
xY6bXkEGojfVhRFQoLoP3wlfBSOz+mQAqzdBJ8RB2wWAeAMOndWY//mtnCWJE/q1NTdpZovzAGQA
60enyQfFkvt/vJt5tfZTW9l1bjWkJkqZUmj+4tqQx3MJnW4jMb3POO7EYZfiyQUWNW08MMawO/AO
RUV4cLdzQ3vo56MrV9EoCpo5eSNUirMgxDg6FBPdN+qjZhqQn+qtY43GtN4X07/xOd17Qg2NvlyE
1dxMRY9EZBJKAziCd5LZKUqBVNNS39Z7dhHxEKKFp7QI5UE2rrWtRfNe5v0ZNZRk7vyEyGMLyMBH
CAua1fxzr4UdMWTdq6J8m/RWvpKC6P/KkaXMpK3d7l8wfed36m9AVsvo5UCG9Mwg+/OPZt9Ihfj0
9QhhvylJVgflTZ/78p6mL4w24zfXTnU/3ZWMi91d3YZHkn2AcbJ3ZC06aV7LZzsgmTRfA1IGxufq
+/K7CvEoDzVy9HwMFk0a7yBXeGcLqyVbgOJlMUt2QcAvgPYJosbysk2UZkk0vepBqPaDjbUqImRZ
H8Dl8ddpauFKqEnqoF4sFCPOSpvSanbzJjCMKcA7AQ+C5auEaolclSb1Of1iOsF565MXDTQrCr3I
mu9mj6VqZ6tVRP/G802b6ZX6g3ZjygbhkJxWvTEzd5AomdVMFDA5ZhqddILDeyvZfvHF78+3h2uO
hwPWbVcOlhCS9hQ4qsGlGFTov4AnYPltg/NO3Ycgx/tX2Ez6J8sB7fLNS2WdUwCnYNMQaMX8C+Bk
2PPcJvhUKZaJbPrcECpEL9TGq00/rcerIZ+HsGvfbJrAfHls97K99NNCWgxZ02ronjIFM9czcEM0
30M6kzj+scjQ5olBy/i3v9r249RE701vIMqROj7ZD8ixs3yZAukEophnOzoM79KLxGfzHHiICEMo
Cl4gzaSpD4VTbw9GyxyJh29VCmvOkfqXrNSEaDfNNtswXHTqfLeZ2q+eubxeJrd3oljD0LFPqLna
L/dkBiOR/vcLaZEP/gbQYIHSgEmRUtDuvkH7a4oeCqATjQ/7bVr5FDAviLOJNOCYkv0DxtP/GYRX
nGdLQpWH1qrhyBz7ZgoPXMiIAdlMFtS8X3Kgu+Nuf2MYEQV+A3NK4K4x0bZne1VC1N8vV5uTsGj5
nEr4yam1d5by7T3OiFK2bWeDqDUtWyXu1mT5ZXliIMmKtrEQdvriXHT602DjSbYtD7iFCUwE13zm
m7TKy4Der1cfdzUPdH4+XOP9dGO74PQoMZXYsMc/r5XMTDCG+HNAinyOEmJVZQfGUto5zcoPMrL1
+2FI+jZUN8kRIWePadWhygLFqWwADc0GsY8uRJYgs93TWNypdncIHqq5aaL5QEW26UoJjt1vVPe6
+Co8z7XCT971kbbwmxzuHEDrgDApdZ2Ybu5aaz25A/fNNXJOwdlQwLix4o7a7Jx3QChJnIGgZtGx
1ldglWRUqz52MQbYHQG+AcYEX2CxOcC7QXeaFx+5/IHhwCrfrW8nkUA05J1bzmt70Z2cscXq5T64
SOzJU5MMewvnIgDfUjXENEXADv/DHn/Sv3awJ6ieJEE/Jb9Sb6VOEjiAKOvEbmU6ni3AguOvYRLg
pPqUEaf5O/YOZqBWPDp0Vb00jdyENiblzZhehraDfmwPNQLYyk36TMDCyTwzcq0tlePBNeSsewlJ
jCQnCELa0w8lOvjgaxuapI/+lo6TmSGo1XNPKGIraJTOl22WLmx/j+n81MTixFhRYioM1f8Jwc+V
+AiOg+uDxBgig3YsFWG1WiIca3FZGXKdOWRjZYsyjfnFY1vc0/bKkCQrwnr+7NDmiS5Zq/Pz1nCR
GhgmBDi+mjXI0iSSsVP/ExgtITuinOu9zPk/KIbK9Au9BlSupxX3fOHAtOwYW1t4z9I63JB3Q8QL
gcxQCj31dIlJIr4gmuImRmebMv6RX1y13ahPZCmbexqV4nD4ay0apyu52i6+r9C0j2dlQqQA8ulD
XT9/+d3Qc78WsO3uQljB30aqo0YJsGumVaO/PM/emUAylKsG9XULHcHzQL3DaRZyP4Lkz/676Kly
dDFZF0jPt1TeLTUz75Rcp4vQfiGI85/MqNuBJQOL9jsbbdcH/cimUa3rZUMB/bk2/dLK+XM5X3+a
FHWcQpgVWOrFCyGG1H8tfM4XeQ+u1sF3tgEXjQROtr5U2In4z1W5ndmxWVDR+tFqXDYtOy6VVkaC
4/yb54nZNiymTCBnm8b8fMjqYup2KevIw/11LaoueiAdayZE46kbgd5lbTiXwpEGNmmRgOwpkXBO
cDzax6f31pS5IIGQ6UN3MOQodF1IlQCCPBIf2+x3uWujKG25CWDSFrg8sD+k5Pa4riXWGk0hsSyy
7fX8S6OpozRzzGdronruwcX3KQxXjTyiliVQThnVIXuPuiIElH4U/lq31fTiHMvRIpgSqfvazTaI
VNhPp4pCZcBDQqixk6ZDUL9DvNWFpAIIE27OpuBDvZixlFrkdA0+l1Cw0gBHpTDnx9DAIDBBnaHa
QCB2WlrUZyo7MA2qP+H7zLGfwLtWV69L2P5dCSQCl+ur7a42OmjCSwD25kbPrUX2FNnI3uEqbHxE
u1SBKYgmW+rawqUVFvUusT0kl3GmBVnCb944z6xOHfVneU9/qE8mmmLJb9437C0/PSCStLa7JU9K
r2LURPAUDS4A+PHzO2PcZAy0mJTggLOsIhStP1XWIa1D//1bKUlSwvf/VzRioB2toFA5K7kGjetH
KsuXUV6QCA6FuipupoPmt8EHBSFbxple56NKqBd9COP8ivZOxKeK3AHWgWsaV4Zdg7TI48FIX56q
8gVF5Ad085/gU0V5t/t5OzRJnMwoJ/D7z+eNw27v5CXBUpq1hRqcICeywuoCTIsEgKQEL7QfLhpp
rm9sf8RyzkVwnG5A2E1/43Fsh4AyPoCf4X66el0byJwTOKeUig2zeBxeEm4Yev0aE9vWTPta9KPg
mPDlmniNCF19UjmYbYUGxFP7YPhMjIsRb74g+p5Jf6tdeGW6lwlp+zDqo3guyulQftGSdHTePXk+
Frs0eVxA8Pyp2Oy89PfWvOnJKSs6fAf/9WlyqHpZ7v1NX33WioBuAHDsMxOlmS2txs60XWkgk+zG
3s7868VuJnPrZdbiGoHWMu9bXYo0p25BUFwOrCOMkPOuKlu/YxNavc82s5+zpsXw4w4uSdtXwAmW
npnGzTrt4JzZ+p1Cn6mvqmdO74VRPcUzuepZxJW0IIWEYcjsOltAkJRpie/osVTSuf0PPJt3QJOs
GLjWG6gqaxMlr5I3wA1aCb6VhFDLUCviuPjEgRbU2ERcfYkkhs6bZsZHBDGR/A7WawQFEbwBQG1U
gXuCcmKkEofHsG5nojPfeZoA9+/UdW54FTHwl9hQcTB0BR6GzFU6AHrRHKkyhFlwAx09ybOBs6yb
w7DHdqwhtasO48A6EJeapTe8TfhjKEVmhlekQqOKCHhzYKydLpPR7PbCEh7hTL2ZZ4r8VFceBlxH
55SBc+gFqgKKhBnbghksPPfSYZlwtMeDc6LcYBtlv0UrfHntlZptBHGcLzBwo5KAy/TAOygo4fJU
0RnTW0C6AXiCD8tg62AxFriFkvB0fb9jWJVp4o4r9uAaFPa/9BDYBMca6V83E/61IcrL8qJFmyS2
xiKr20pbnj5hYkFjy+NPNMqiaeEFt88JMN5lglPSjCYySunieHC2HIubq56APGqXJo/4fite1efc
8yWp7lOiaybWB+5zIAV555qYS8v5NsE6hreCnaYOj7AiRYc9U3WhKXQat4LKuktpLJAc+1h3JqKi
auJ0Ojqdfxu6obTSJV9B2y2F7yhhLdTRleF1WF94VBCDcn0nw1/xZetMBjYGG1hlfhVAejosXbIZ
5Lh5YcW2HmsIOw7+SWLtBbgA65lvjA77crGZ8OtpWcmyUdAMmbK+sdP5cfoER2ivwyJvjhJDzaCk
PotmG9cVeMBvAOZOa7O3/BkmFBiDseDKiZ7KYp686w6E/qcM7dC8hdJ11PX6Q4TviX5jykCkShL7
rhFU7XGc09ZS7kNPAV9ulN5U4p4hZDvILwyMYmmsMuJS7kIKZvh5p6BKmyrlMho2YMjluC4sWGWE
NrmzFNkfgi1OqK5un3feO3tRxHNbUj9habF1wyIaiwAOGyP0mLrtbGJ0tuSzqm+CLbgcG1pk7xxq
D8TXTk3pLayxJmAAcaKWw6fw+R1DGbSbfByccCNt+1vd6FDSDPEdS8Fas6lBZzgwq5fbQRtVrzCq
QMmNTbdSy29wBGyWUomN+2mru4S23aKadWhmn+xKngcbgej6Hrc+ZCAdnOG3oAu6Ai+V/QsSqBaS
YqNFnk030w/oi5J38CeS9eCc9F5YQv9zEtGsZT4F1qnAbUfjtxnoIw1cq3E0GpwV60lrfHsJtOlw
M+/f+fsjsaBMKaY2Au5xzJworCKO81EkFdybYweBPSlGWDeFS79T2heI9HWCQykdfRuNkX2swsLc
FnnE1ICBYqkP24fuVQM/CiZl/JPbPpuSUt5cNS7r9QXajeQMVavA/sR54MVyKLaWvxG/zqMC+6ea
aM0jm/+8zvW7dATeIcCAseYr1GfaKZRb5B9AzZ5h7eFctPUlREY2vHGU9QBDDQeuRZPhc69X3mjB
1uSUCOpzFy/61yfKm+hnUSn7KrhZEmJbVQPEX2VVsF1eYTOsMlNysl2QnU44mc+12TLo+AsJbThF
+O11Y60Gkf3mdPk9LkRQMIgh4KtDkFur/ivSQF847LMibbADf6TVSMgTRP+RH3S1z+t20xGRiqcn
QKIey+yq/FFS937KEAmGEUGG+xaRBJK3Ep/Hz/ejdmckTweUmpqv/vWuRpe7WM2T1jtkn2iy2mSY
jWBtQyC1fZPDiUEKvF7cCooGOwOoEYtL0/8+s9Vsapq5f80X2PSfYBwObH4NvNAVDT1xK7Ehn/om
XY061YEaeIV57A04l+JTfcbAvUNZMOeB2ECi7fGQW6Zf+KjoQu7HvCJvCXYyDiqXleLiLHUZEE3j
sg0Euk2HwqkhZi7nzk8IyN9HcGNjDY82lUiULfTCt1a6W3I9Pt07N0e6n7UwYYrUEWls7zStMB3X
qoD4Ni9Ykh0Ipls8XynfvlPHlaTTHKzpnIvVQyofWoq8a1LJPkUp0sscVaR2XuttY7CeAUFl1s3y
KeREtFPwq2p6UzqcFWB8bqJK09spUcU+3JgSUd1/uc+lFiYB3VaEX6Qi1paYcZAU2iHzP+pFOZls
o6i8W9K+SgV0yit25VW99TBcDeGrL76i4voJz9sYe4J+K3O2ICqWaecfSyCQ1sSMBW/9dwv+ENUF
Otlr9rv6f4Y65plaxDJk6nFSfVn6ar6j6G/FB3cpy6iMQN/erg1sTpJpbRFd9yz+VSdBNpvRPAq7
Cq5GJ1FyOF1UmdH4A5sy4IapyZI4G6V2FNnGgYNLJReBu/lC4kZxmU1T43wtvgJKmj2lLZkYgGwb
yVSvIl4UuDLNmlt2f55EkB2CcztbEZf5tbydSFS3pjnshGBPC/BnFIyyRnNRmPqIKLxXS879BXSI
MNSzeo8dnSdFQCbR92h58Vm01FEBjcRDJi2FHp4Uv/c6W+tVEWcwJ4P75t4Ard4Qo+KnMsg2/ycH
JQZCLj/3hyyfLPCAADMBpJap7b6XHjwoHvo1p2kCgIM+NTFVple/kVlpAX+IZuPzIcAOjW24xU78
NOvg4OoEcISsec6PzMa7Zm0ElGqWK9vs9ZET2mDxH6lJtZN05tR7IuvySUz5K+OLAmjp8t6VREM6
6bsKgS11XMr5WQl90vmVo1PuT7Xh1pGawyO59o73hZaaqS8m0F3MWdyHukCTlQXOqxIXiu8E5Cp2
0AxhC0rHZJmQv/XpPFlLeVV5+ZDY9g+LfV9pBzBwKJvgH1pyKF0feF9VWPc04vaDlwQ/b52NGCq8
7w4Tjml8uJzT5MY5XMFeBZfemE1KQPDtdWxo2u+mLqZL7P9UpIHskY4SVl7qLtuDtGdJ0qo6Jo/z
AdMvytVnL9UlcqtOv5p2vhtuAft0SpCQNm/ogzuh4KMu9WKreCj6A69I1bf0n8al+vGqOWrSAk4u
AiA7oWeDxBOdwvc973XqTnY+JTAEMFZmMTlwy/Z7PPnrE/2vJPqny73fnmzYim7jiwtqxubbHJLr
S+twvTIlaNz0rwu21VJUxHjrO9JLZHq67TmiY6BNV/wXX7EMqorhn5jCsWMzKMu42FGme32R6S6V
o3N35EqYKrjvTqG5YoKTdo+lC9q31FWqwMhMJ9metJdA4LEgMLM7w3NH1iMT3g0Fj/QLYbjdaPuO
HN7kmC++lE5hV3qm/my0MCC26b9KbOcofhShX20/QddPPOTD63QE4JFa7C8b2XKPehRP1z5H//Qk
mhMZCxe4g8xXzb6FTpYS921b8GBJ5xuIVKdStaFr2gXDFu8IuwNWkc/sMro5LCoHwnFM0d0sX+dw
KyvTBwmCy/OpgdjesY9bjZXKif4QKgTaD/YxAIeEl+lIZyXslb98dP+ikNCx/sVo8KTNgnNUCafH
OH92xITMRcY38fem7EflFJ5f8abx6inYRtZrg1b6BaRQAi72iGYruU2JuW59YnpyWxRiKO7NoJo5
Nefwsvz6x87Hn90r0UeRFLDQM2Z7z09h2Ia9vkl2xqI77SHcml/hM8J/b41h5mNQ79AaEO5ZGYsT
xf903Xuq5ohGoo4CGcVd5b+R2w3P05Oc58e8QgwRSe6LoabLY8hCYOoct2C/3Vlh40zbYCGPo846
Qbk6RzGXEFtzXn+imAg/NEE3E/JEHu4jHGQD42PSoZkZIc+37Zujsn7lu0JixlKBjISbTFNmlqia
EU8q2WQVBxnKSUN4ht1NU94E83yJ/qyDPogok1p6yUuA0/CXpUmDPqkv3yb4eMXjtx1sbfDAfNCd
xcHGvh4XCdUttmY6Bq8FkejEMpqVtXbgidJgufWlkG9j3R+AZaU1dgNaI1kos8u5XTlM5L8xnP+S
qyW0qlroiCU6P+3oOGDip5uRSwsHu5Mv6lzeu7OU3zi5Oa06wrM++zbYZeBNNNSJDr8o7deAUWj9
pD5KvyYQ6kGShq7PEz9lZ7m3XVu8j6h22fdGBY+3wlvERFHRKZji/GwDvQS9KX6gdX0WuzCeONNQ
R2GwGm5thrmdnyhn6c5UIhfoc5CmCNQ5b2tX1UD3dArEBDuB4DTwTP5iuIX6NPrjSGkjyq0oPh3A
CdN5HVu6gQW1Bv3kAC4cbKRreN2z6djdlElZrF3SovUk0+wKMbDLBO/iZ5TzpwWJoyQgV1f8KU+0
LNrmLroeZTOGZIoaAioB7jp2eDqC+dtCSwCmuUQBOWlBadMjO+Fu3idVCLA5179jezD/N+IykI4n
ZjxmhRA7zmNYv53TZCX6JsQeNNgW3/6ftxdf9qVJYnTMW5YuonMfIeJu505ndAAhdqQ9w9z39zol
GDY/xRuBzGuH+ItDVLoBuCGyjvafEpT90iafxAUey1FwKgXUgzB0eeWahafS1CD2qChb3hEQfmi+
PqO9a7i2f1EpoRS+iv6T0/z5EPzNm2IcKhJZ0jo2aTQEKDg+D65Mm2XnTsxoKCuQcRDEKWlicA1H
b3e4uQLoM2yY5L52BvPsvaenSg1gWlmRS94Z6yu1qNlcOMs9PaOc7vr1tnIR2v0NyHar35O5D9tC
6GqrOpQ2CsQPYyfaAEcK/tqK8nxtucMk2ZlpXEv1V0tXXFimfjQEJvA4TQ5jA03cs4itTBWBLpXm
rivz8HxLI4o3mXWqE4plgUPUMN2k1YxeYkRe9Yvd4S47PqKxt/CTEdTFmFzRjOlZdxzJB2KnNsSe
k+C2ub5+6L6+mkCF0OC5eg5rpocQ85+gSVv7uEa+qHlM6kqE9Zju2ifIpvjOaj7Rq1qjNHMba268
QBCq1A3/0KIN+Y1copk8yuj0oUxZzNu2nInvftSYhoysWECNuO8HRTv2l16bkncZNOIVhgHxhiTo
megV8XORATOsOmxHxGYArLmCFMsbYuPFANXUysxDZLOQPQx8xgbFEXBxiFqqSVT6kPxgMSidkzQo
6XUTHcwD+OPPZjbhvfinSrJLmLxQ1TZK6zRLrpRqKX2NuTtUkTsaCbD2qQSUaaamQUZcq8Cx8t/D
e8Hvb8sKu5XxgIYhSpNKIKR/4lG74zdafYJRcFMandVmb34/Cmh21SXOiOMYc9d9nJBA0ql3qvU8
mitcMiQcSkzATeGgrKJrBU71oFxjw5xWNOC16Dzc+IuEGZUtL+0Nl7QddZMs3UUPjFcLCRBKA9vt
UWcPE2lB1VE8oHjKDwlKZKw2a8MmVLcPFCkBkUm4ObiOTPLzseR+cuAgLdEUwW5it01yOOoR2jb4
gDp+YSSRZbBPrYVvpt/PJbJxWqMGsmEf4djxkLlmBp11/uhd+15I3o0xoLZNQ8NVyQjTlxfB4kLW
Al5wIG4SY/CHSYaUGp17xo4GA+cPkHSEvJTDz/BiAvHcV4zwV6joxD8WOKyisqYLtk+SxDrDoQpx
uJH6XF++q58agMy4bsba7LyMqKjCMmchitkRcTQGJIPPzptwwwJ7JYWlVhMKk7TyNU7o+byI+Ax/
5jaV/dzecLWepHZSLA6ETM74worjuKP6Mfs1GMZt6GBz+BMPxugFfyVTyCnJfQ6sFBoLT6lDNPy8
32vyObr9izNDYujyQa6OU1cCXfuBR3mlpxxv6/DDrEieNowRQSVOabRIlSc5x1Y9aAhQRib2P+9E
TsKI1676zo1ZNzMR1hIkoryVgzTZjqJenkJTJyejFMLqnZutfF74PzICqqaSN/1Kn3BOhnaWaHsO
emoF4F75huk2jznLYdN3+R5dv//QVW0YH7BgZ/j7lxK3cva8liLpFC7+pLyWXc0RB3VF5TeyBwAN
cn6wlMXYsFyRXpqP9alGIswl4UC+mtMRTSnqmiEWz0yxOMlseOvhrmJk6E4cGhMJRKDeQZQJDelH
fdy8Nr1h6Vy8bYSEE+Z1F+at2FDOybYpCcKRh7pwgfGs+wmURwwqc5m8mcPsZNuiNIQOJP+MtKDK
bciofvJtz9Fz5T9ct+0jTm1/2Ci8bwPNg+JNd4RYDXOsjA4KJbNprGMhTmNtHs6RdPcFscKVQjNR
y7Cus07x1NLUnYP6Cei2nVHs46fZbqX5aSG6OGefwQXt/49lXpMYQ8CY+p8wxeS5kFJUS1mGrcFA
6umSvTM4vKxTb6J4Z1gYQx+mXV0g071n2+fsKWecNlJzKsd2UPl1u3uI9fHMmQ+zWfPgVvWLUn8c
QKkwt02ABRjcC05JH5U/aXEYCNeRrGrEXcf+F7NtY0/WRC7L/c6/7e7Ow49Gd7/ME5hy/Keew+UV
SXZljjIVKgaOlkb33NROlCSboZF67m/dQyQC16Z2ek63Z0MJqDUCi35xb1Sv9cePTEyPqNtOELgv
7FEqqXyjla/BqcRwMnkqGhZLUn+jY9CcZ20JpuTjlT9IOlyq3hO7n+q7cmtCQm2STmomiaaPrKXE
zaXIjy/xcM5nnFQ2ctXePhBR8mm1515kBMfj4Qcl8xaBn7xfMM9WLGmdnmSFmm50i5bygINpwpAg
upJLzGqE7r74+CVMYCLDsmR9ZOWYBVCxNR+f/ki6gMnwg3zF1DveMSnkm1x1aIil66rioEVFOBkN
43BK/D8q6rdcfdavAhFKEF9dXl3MVWvLWlByRiCR/KeovG1IAdDOWZKwhZhyt0JkoZfCGWGkpMNP
vCgUzOE/TtPZC0sME6+LcdFEeyNZ5Dud7yK84cm4SSwbvF4YrfbiUGEKLBCg9wG5AQTsCN6as83/
pNe5VVY84l9k/UmDDciovacqVrhIq75KZud7zJp2R3DxOZKfHt5WqpaD84rGDWCTTYDNc9k9yQVa
YUoh4p1d5CfOzgsQT9+Tc44KiakeE4Gq8faxYfU4Uk6iwA/kppQqC1iz122GNifVdCVn30Qx+zDt
0F56CX0K7+eK59/Kz8PsYBdduTG5O9Ab3VhodspROCRuLuAATnj8qv52Fk+gi9FUsyevCcDsxQ0a
sGeS1XOEypm4Z4RwVTlPRInB8Fp6F/gxogcLgN5lgNq7EhKH920Ke2CMYbq6QkuzBBKCnqn2SV3h
D+k4Kprlt7C4V6Dhmax5W3+jDYSbD51u5ZxrolhFflgKu5v5oq9wninisXmWSv1Ay6eM5pO9rJof
dVe3uBQEt0z0I/x/JVkg8W0+DXBOeD0447Lg6zpeIyphMmYBtrIyOhoss0eAEK1BWVqOG8qocMuB
LIjxvKJ/R+HPjNbe+himLqSmph7HQOoV9jz4TqfCPqfqlV83ONrCpRC00vnxd0mIiaDWGm75/HSj
4mt7fSC/ontVWr4xrRtnQFAw+LDUZU/LjM3VisxHbV+anzHmFtFWAnIZ1GgGz8n8gdGq6tELKl3r
terjZw4v0VtDtsuGoO3V6PM1UbXIxq+DVZsantdw83nGJj5W03oP/cY7fPMuMaXINGzaCv7Hdnz2
muZT/5R05GvtdmIamNYHwtMV54c3jtfnfQuXlxp4jopPNiakPFAN+HB59znI3PNP3uwK43vY52eC
L1c7kkV2DiKTl7hrnxOI8Y2PRRZFVeADDvWMf6aJjVmEjMt4E71RwxIb+JZbwW+tbdBJ7lcrR7Wc
6l0pFTtSHPOrz5CnQMX3xkCYDWst8Ewj6yu32exxDNvX81moX5jougPpZ3Qs2Z9ofFBklAe23oDe
QWav5QprlAjMN3Mbfz7d5TimXufYvwNnmIzd3m68h63kvshkvvrVH3JR41yzFDOQ1HLja28DxdMp
vk0mC7Y+67+sd7hgtlkvQkM8FT9sw9lE8VphqXD9/v3VEvsf91Eu8KczQV/eaVr9XRZIXhh+nwu8
TBKG1gKdlRm6mQOihP3QY5YqphDWCT9I3qyuxNcEaJRl00Sf99RgYdk4PypMTgA2+anBRgqAOUA5
dI2AYUN+7DlIgythg/LSNnb2tNIDx0aJ2z4qRlr8u/acooCsGa8HwZTG2tk/xNpe+7femDq8g26F
E3W30ybTNG/Um27AFp7gKkJaJ26XquvFhelC14XtxRrVG+VjVCdo8f4crkLgUiS8KLP1Z6fBcFZn
JuQQ+YiPZpeLtDmnzpbRgxv/kVszTL92CMCdeIikdgGMA8EjSkCtg9b6uj+tkYbQeImCZYYVU7p0
T4ItY10MHbeHVk0FdZftuIrGDdovOWDbizClXspz1lf3i8VWWH5wg6iIoq50Q9cA6FiMDhd4LE4a
2Kl5eSpfeq9UHDBx/7xGEtkVWe018dB/6nFuB0VCZxl2/KgtytkK/GmtLsYKO+Mcj1gpQGKVAilz
I+WL48bvrl4nkSL5Yg8YTAqW+/b/yh4fCvEVDWdY2hbADTsCpR1zfi4hFzf/0bAtOOOSeO0tm9e+
pjLiJQZRabQWtmvEqf8t4ib6tsoEoGicF4RTMBpufaxJfY68izw/7i+a9ltr2wMb58XzTvSMqIQy
3MDAxHHif61l/9a0Mhbv46eJkwEc82iBrY+rAcJQJtu+9a4bmS6oORPLvliQEArph+TdpIN+6wUK
Tp4dN6JVuXpAyijfOh2uSa2rSJ8kpfj9VuMcH2ZqgVgnr8KLPtoMMn5yfb/uMv/j0cUm5EPUFV6G
F01kRfXP1UCqA1cce0eTLqQ9jfEekwgdRdv/9ajKWVwSZ2PNI4bIkfNuhn3D/jt6vepERGFZYN85
lDvcSQwvT53K3zB03+B3koBZl6baWHiy7GVcN1zL4VtvkCskR8lxt9VJqQ5vMiT0v9JlebMHyNxb
PorQhI2gmg7p9QLegCbq9UjGR/JMsIoCypu8LzzsJGZfrqkFYinl/06mYEaFGDsFkwi04XIXGVDT
FHtL7Nwx3BT5rbzgrJ7ZrpiTA7WO4RKqE0vcOmkJ9vcDVQOVqIErgLg8toNUS5CdHGH2KnYtPzPc
Wy9jN39WMf+rq8C4LIYUYJ7LuzqNNrlrmaZiojdCLDBebJuTAIjLOXWiMIVZ1asJF+IJBY/fb1U4
izQ2n5nvlCD/duRVk/fgtBcWamPpD/X6AV7DpAEHgg80Ri37+kI2HWgUO4tEbaSw3dUqQ8KYTZl4
HLvQc/c0FpGQSQTpdCrOp2pIOrfo50JESI9/CZX2TY+aGCqiw1v+9l6QBiWQoNkwAwvuLUstwukn
cif1PgXgOKtSHlr9Yor2sY2lKX+UKUdhNCGUjenKaCD8cEGTOJpksiPfwz1JJQWVOwLtl8dmtLTJ
nbNgR48KKxbEvRX8mz7hGKroy+bckFtqBKgGjn/EWTAPUex3E7ZVryiHUegRVcMT7kzn9eWCkvP7
mO6G/v7G73gDRgG9NLnk7CGYEc64JZmYdy+QpHC5Sfysuuo/OCkO5YHI8XBrAPxFZEOha65mL5A1
RaZFcQbQtC0YOnemWpMVHFJlEAjPxIBquShs1VcBtKlm+6D2KJESI17gLLAs4yjMT5cFA+5e5BIu
9VX3zusV8D30yfL5GfOF6hN9M6b2o7QRYVrrRKkCg8jOkZ5643qNpK+axytwUnq+xZQE1ZThXKBQ
D37RiBldO6H3pAlzmRT2tKaeDQYLBP65WvpPcWZPvRMFsjyVhFAdHOfujwxnpvMR8S2rxSMmsN3Q
OdbQgHxH8PazYRQfp51EVS4s5pqhZVo+RLc4nH6CM5/MusSZ9LRzFqGeh3gvYFtBjY4Zu+Hy/cpJ
JwgvKzBNLO2yj3kT7RbUpclRg0bgjOGyoi0vVDf93oYxGa4z5xdF6pxrGgsE/2BK8OTOMXQ0a6ff
/R2XpbXOnqFJgwBGq4ZwR02ESnHXVE4bjM5nLgcMYlR85tVncsij6CY6NjXNs4wHBXFLmSDe7ybC
EgItYT4hAYIa1JiHIa87wkKz3WVV0n9KWg3Ik5xcyox+dMT/0qTpOACyQGZipe8C+emZx5kRrvym
PqcZJN9OtGW91IE6uusvFC0qZzVG7hWCCjoErBxo79EpeSJDUay9lRkSp/eu2oDEWe6rlczaSUGV
0CaGFofxvgnNXVMrp0IZIiproQlPYdKTMzGMJ5G+ToAoLEi6KkBmNGW4Wza1LXbE4Sj2UZIYRGfb
KVVjfREP/rrZq8+xA4PfI1rlUM4FBcSEHc9JrOZwOpaZG+jW7Pu02W8qjBH2AZaM7/D5Uus9O1ZH
MlnIYbIgXwSgCu11x8BknQjpvVY4Dphf5B1qcyoNifKgiyX0D5Js0HpHP/XuKXJO6EYgR+0mVSjC
RqSa/U4rOK06mcGiGGsrBPAt34/b5oihqtdN806cI6BFM4eHA94b91H0Gds2kR3lKNpZN4zQwjjA
NJWMFc3GLH4t9s8OHVYsUIX+TrASEiJvxMx+wjjBLxwqlHR1kM3yY/WJWKIGrmpCn1y/1nLgtw3d
646IHBzquLT5fweVze2ghxBnlMIM/Jr3NK0PJ30roDkhG4t8elGl0qgcJ+0SQ6vSgPfrfRzOqv8n
yDZYWuhtYT6m3BAasdLwVqmwOjGUSSYGWJdj5P52Vpm4vKzspiFkzD+Qh6Y4MlCS+J4u2E7XYFJQ
xdYlo+jWb98EaQ1kNiWg804tWjqP6oJmhCfub/P3c975elK70SYGMk1mRcLQV41Zyc5j3X3pw6pk
VLqSgPG3eTbfk5iWGNl40eM8iJmpfdis1uSOGyJx+LDjpqiKAZW82Y8moktYl51XDgOZneyCJNmw
0GzsZlt1HRnTVEtaaqC3b8inQC5UNw+uOh007/lYcpuWw4O/WmvVf4rIBNt54jxSdh3Cg6/sKcHW
aZ64dhIoQIrP06Wsil6f5MOrvcajaInCt3iAN/zm1NjCTWd9Tl/Mrxi5HD1QdyqpfoTM6HL97gme
ouuEXZ3rJoqAN0ZkfS7FRg5Ch5IwyPrAJLIionrhP82aXJbFIcVTFNiW+Qx5opht/+tqnYMwv8Co
qLxRrjdV52j37V8+ECLkM/6PXOjOvsRtHla5nalA4GYiQJCQf5pWn9xml58T+iaiwc/athjL9jCl
x+HYd9Mj0ryUr+2eT/F8R1MJ5Z5WmNhX/8XqC6qctzH0tlQncPjK0M1Zr4/iqbMBAsrOY1LuKq26
PuOQDuA/RMFYS2xmHWq6dAOX9+v3Y7YVeDu+VUTssI4gUVs31OHz11X7U/KifOYLy4OKpki8PeQr
16WQzsgdv+eo2IPAJbIZAHk5NIO1np9jj5O4sFnAlzqRMr+cdrHYUVAVsksgRx2LtyPgUydK2i6I
CUTbRTEcZHrtdJLSON4ne68f7Jp85W2e9cabfoxCKS7WkJ368o9TJ1YPZ29toLJczILO81b1M28m
NyPMQ3d8ojLcEmrBKhhRnlXW6Pyd2J86NjWc06Us22x6d6JaF0ivIqNQxYl6trbjxQxr7BWl70q/
EprCB3a8YgqEQHwaJl3tIyWO+BKTT/VRPrK42AKfZTp4GWRnT7k6qrSeuvsGIiepoZ/v/yzn9STe
W5DafMhYTuZ4SQMIVkfmYQuJQ+LLuVkTV2HViLPhC1Z9HzjzHBOQfiayvSFyj4SG91rYvLgD2wlj
wdgrfW1sZlG/C9yshQdM4on8LdwIKjeteaqDKqJLoOnsWfRNVEv5wBc2sNG6Oty+McsezQysPpVn
Va5thsriBIvwgL6gKBpu+0tDSn8QD0JhKFcDNkd/BsqUzwSBUg2sV/Q41K7/sKK0JM5FfmuFg/WV
MxhPC7jGZaZyh4y9pSCEWXKDdZ9skuDE0ETZwX8TLTZXgxHCxLpe2BbiTErRMzL7KsAJIt0cpt1m
wtmDx5HhJFS5009RwIROcSWJazIPcAzXu9Eq9CEnd3ZkcoL5SC6oSfGWUmjIS3JTFPgQ6BKphobm
Vr7rbt6QGfXmNOH/1mdlxM+mBtejSIqiVCYk/qXZ7/crmT5k96R3vLHxvXXT3J85SPn920Op/HOS
t1y32wnfCNcHAPdM688Lm9ZKSPAkl84rpaW2TegoeuA1CX2bqNARfWvsAkZTiSDg72ngizCSYitz
OyyB1ZbX1pHbuMUd9z3Jf2jW3d4TpmFAY5pXD4b2b3+jDHUeNtY3c3TKIlDVFauaaRSCQV8KQQhk
d11k8523wMrT8syDrUXP+sfsrVQkYS7l29tRl5HiCLqrxxLnB24FGuRyfabIzSGQ0BMjKIFXvRDy
KH7JIs5QQA2P5iq3cZtuJCc5uo0MloB5SoFqneYzQaPTJuTKw2OOZK3z6+frmE0JYIWtFO9attRA
Lr9iXARzW6TVd3Wjnbfuc4jHAQaHa53Tl6PP0ebCFuvnN+IQMRKmz30SK8eA36XlH75YtqilASp5
DUFl2aZGa/fCshF5UF8iiyWM3kxwhfngLWHdoPCX1UZCPE/RW2CQ3Qu7JlCzmMo0hHz6dvoz93cG
hZifMItRonzAuCFomtmBoi1xjeHKBsnPfWeEkaElIBg/xnWfuCcwpce2fHRq56fBsM9isIkacTMe
QkrVZlP8snHTNVcQ/nDeWvCm+fn8fYACDili2XEA2TExyZgsVXLt3uwuQFK1GKv3DCRRE8r5QpIk
T+gH7rk4J66SEkp0BCfassCDGOMPqcMH+u+a1IUhprb8Xv95XDzc1kQHBtuv+fF9n2VG79AltraE
U7H9hZNIUNO9MvaM6wvpay2k6JmEaSzb7ZoU/hyDknRUqhGQ67UPcZrSrT9xyXIAMY43CFrAgSXX
ryP/TqPpj3zlYjDm1OttMuMkXlh7I+jEGGCqgY7Wn6fo6HVQYCBgoy0OdKiruS+ZtwUD7OKYELiQ
R+P9ZB7RQgf7aXudtaNDF/j5zyjTySUzHgCbwNCj5dUbf8y0NZM+bKZV/NCO5y6vn4FCREq5wjcN
B82OlQVH8o8WsINWvT4jStfNt1Vm2rz4fRnx/HAPSGZi3kAMOBn6Wuor+rNtQzTdYEnS6ibzbD7b
5T7icYLmoBy5ZeRhQL/VHKP+nHxX4k04w9rqg6OrTX15CUll8Yn1Hz8CwjxpAGA3mml06/lgfq0K
pfcDYt+BCHfha9wTAlmxCq3HAmuv9jaF4qspFMoUhh9812igq1eOEc4Ue4xwOKCSALVWg0hhdobV
a/jF8pOVJueKBRer0ei/WmYcEpoRPOxXUNTbsd6lq0LBbqIGrSmVaArBBVHVSgYBUX2Lwiy54juJ
qlK0ucFrtYZlP/FLkqhs88Ep3MMSEW1cubCVQEcfw6z8GS4eOYEfbScwf6xh+7+FWq2OLI60APDL
WWgiyCwE5Zwi6ote24zbiTWIBx+Il+71M1sfWe2+4jsNMxO5USgno9klSZ0a0TQiTwajqhXGBC7x
CSGz9z9406vGRES9lPs8QP9v4Q7841SD+KBabTZuVjLPXNjU51i4hpkVDly+A7q0Ne/eMLlXAomO
cp/GDS6+PEWAm983NZZJsP+Ch/a5gaFgWjAJAFX+Y5pqeHTozdH9T57+sSJMmOsPCtazqABvvd90
edWu+acCnLKYwqkoJuJSw/Xeaq2HzRyLfZv+S+WBhObKvAWEsyg5NPxXfgTlBZAuA+8JsBTgNw31
n5yIK5If9mv2+AI0up9GufNX85MCTpQun0NnLcPMyKBUpGrzmZRp1lhEEBt9jG/fCI9NPA1tj4K3
c6x7YDqGaw4fsaWkecS4Zh4/DINCsLkZyfiak7utJ2X04G/RoE/FnwG01Xkkek1x7jOTATIv88Vq
3CxKE2VDnOuS331EXPrG3pqv+8I37OQib36OVkm9hG2SQhZI2yxLHH8iZYSe8S6VRxLHrfLQ6t6u
AoqWVIhrL3cBU+K+5BAlV9PLcGMh9OEDfqug1soPJOpvvT2koI2TA6mTHaMFrowF5d6lbZzZ3yAS
sUgM3LLn9CQGWlAljzTNx3fs9Va0LP2xMYyNwgv0X3l+6mFB9RpBOc1sAyJu00KGcP6vhFjD110p
HV4K2Di1AgLaHR0tUR1uZFI4EsBFdPeY9Dm2L+bPiDq+8Gnikd/B4zTvWggiexh6kOj5Q9OC80Ua
gkEngS2ADYFxVwD61ztgvN1rPiHhvPiSyEPqe0xpw+xlRlPR61HkImpKxRBs1tkZuYz40EbqAqz4
T5FU0z+LkOnuTjk+KlO8dCov9cnaoIwl9omVEF1eZZPaKISRLRWT7O8PIGAY7A7WyA9vzolb23Zz
NlaSkwlTjXX/m0LH3Os1nQnTOZZxQWoxOH9VR9MuGWytP/UllqheYub56lKdNP+8yniQc38QqAwj
2s7DdGl1VQ3xEaT0JikUgYstIi84DabM22HBPFj230pJAPesLfit2TyO3KuZk4RpBEjvHgiBzGV+
WJyvKikIGjYeSaunTVlHLhTsWXqP3Cw3TqdZ4Kdv5B6HsuPzFeyb3VUEcWv2vDQVEvY++4iDyca0
XBPohWsxUyoKczHXU+D4g9NdFdhsdtTq1j2ZmQAiiJPeCV6mL9jlEcam4dojMlNuOtgOlgAbp/a8
AdDDJlq+7lKezuFSXQfiYldki5Feg5pRkJEcT4AKTjE8GcYBsM+kI3grnGJ+Wpd3ya9AV8op6Xdn
kIbx+k09vbMkmhSKasDVY971swscJfQlIibIFpoqD3EYzHXUIyVQtnzf0Ff1fwJDjJ1aD9tk7MIy
MOml1CvIqdZ+5HND5jBUKxcAK6iPDqStyW5zrK7QAIrUcNtQuIge39b3uyT9nOEtW3nvscO9+e9T
O+FVzsbecr2++BJ6Hk4cD1lHoZgL7rgGIatnztDlWsUQX15Gcv90wls65uyDnihqDdUUE5uNuNiF
UGu2EdBT+6oMUDtMGTx3LF5IXpsUkvskbZigFlPnMyOeOWGlzt5OSQDpnTP6u0DShAzd6o3Lx/Nq
DMHChVu+2MIQ4Oa4lljKbCWSA4VIQ70z1YMf9pZPhjyWHkBwcZY0e3U8aCEdolGkV4VAIA1z8Sqe
q318GgM58ZMPZ7gR74eMU2Bd6kaEkQOzZY3CP5sn+rrHN4RkOzaGhaPqwiQlGQwWzS4NTL1y0/mZ
DWfnrVKq3MZ0rgQDlylUMgQTRp9horI5cTKISk9i8EGImHOwrtMAJLudZ8D1fTSvArt7lj1hzafx
mePZi6TkkAkzj4Yx4W2MCvMoBldKVNBOBrrueo/+UkmLEionzUug5Y2CRVUrBOQYzuqaJjK9SkVs
GpnsX6nTD03758s0NIo6LuVA1+sKV7mb7LPfZrpi/oGku1zELyZnlhPdFY7nvCHGtTGiLmMH/XZ2
y8YDebVeZ9yACJqDIQk9LDQ5c8/DjkCNAZ0v9yHIN0qPjLYMwwO8TPuqkXIlw5xAVDpQasu2hba9
2eH5urwh3asSoE+DLld3Vr1+r1l+94+zlB7akLdtRc3xhyT3kC4Tyi1Y5dGtbGVUwDVKv2i1/QlJ
18y1pUNUQxWEatQr/ESz6IMD3p1s8pTHKBBTtYypc8EahOWZ7uj3jVTioP9qyKhYPcVqba1gu5xj
KyRXP/ytZlNXfh+vEZ4+Fz80hc6BBdZdIpyloJuJ3LqBuAYwNESiWEKV+uTY4Zg8VXJ7ST07g+K7
/s1+vNxTTtzE/IPBbiZGH0j81+2AFH8PKb+fdo2aMIafKt91yKOPcOVDUm62fk+LizPNfM265PQN
KphxQskYO+Th6q+si4tuDEtnYK7vvkSZN6lkTl+RZFRBT9tyaT3Cd6IW5IemwBy+kg/xwi4+sdnQ
pFiF9Zwj4fXjaEImIhvz7SkDFeiP1Q9FFBH0IUCDyPS2hJOs8xFDfK0r/1QS+VA7rzklWEa1eULa
+Jal/daomkSjbdJnQ6Nz4rdh2kYKxv8kZ9d4GTWZPIAvx1L0yLOdDkmHPLSTd67qAvu4WWPuE4Kr
Q6IXbYCbMfjO6kcn0PYItRrLQsTSCBA1/rkVKPMOYzmEw62zw/gxd0hmhb2KM8gD53Y5FnWyr3Gz
dckySYiUTdz6Rn7ag+hZ4wXKo5sGlo4EVwgF+GNIgtK5TArdzrSCFC6MW59JeoKgUjiUE6E9cezV
WorsJg3BlWNYJjzwRUEGQLcfkDT8ugvLb59O4FIZdYKHKeR0eC8W7bz2CTyYm6yDk7PZHMUSex2L
nryTntK8aPXIZNrB0b8iL9xEuYddJ6/8o1F/XjgCIjBN1oxC30KmZ4Lu6A57mNNA8z/u0tNPxDRb
r6sDUtLjs1netFupcpeQSQhptuuWYVS1PRoCVzC1iiQpvlNOACJ/l7LqUEh3zfxncarurjdtbNoA
bhUOZLUjpiyjTalhVP8hsHsV/VcCK/WSMbRwORpEjhqvyfNlr5VulcT1x0KsvKQcEamfb3QTgnwE
gWMD1NiX8v4C6JN/Ajqd5diHwq+D8UA/x/HoPCYZazIlJFw6oMMZIudSnBErlL8H4Va8FfWS39UO
XeXd4Oq62UWPXxT5ZYnO15XJSuRK4g+9jrAvHjpVkq/51GrlKGx6vl/s6JtEMg2zNf34XvFNpQJ6
1q+LbxQJSLeNuDYYJhrZBmnk/eE9FuQPiwkwHyOMgrAw9Pg204ifij87Sg5DqibzFTzzgN71AAIn
8pcwbJhPn7pOx1g1EsrIOYaPgcBuYO1k/rWTYosi/4VmwjcYvxMmGnXQ11fV3bj2XSExfNtAsUVH
HlVZRLiElK85La2L+dQEkg6p52whcez47wPOs67tc/8gKIdDaHrY18H3uFGa6fiWA1VDmUTEw+iD
IxFFmceFVGKoggJGw4ZJCS9swcWQSmGhlJZbuTbn1Vsrh5WdTJGY1bDonDdN67Vkp+WLDMH2S1FI
mD8LFZ8u3FMWSXHtlqhbsCrZLUgXT7Ih6NawVAD0bboW2A2eb60myscX2lPqzIoFJQKzaU0q3IUO
dKPYx30sbc31/Bg8D5f9sJGxdD0zFRWFciAmuENBcy5FIAjdyHGXbbU/vuN6dR7IQnzpciZNAnyk
401/YolnBgTpeF/vJ8zmYZCszGx518HiCa85uxe2XwuiMeH5ujwuP6sauruY9921icge223nGF6L
K8E9BZS222F1X6dFO0hTE6cJpKw1qHlyxyX3Ni15sMfy1entA2l+alvlD0ijXBSmtc6QqalLENC2
ftni+pUIkfLJLlSV+pTNmMVmqkWPNzH/sapjSkXSvtQYvKk/xUXn37+4c8SUjAMlf/AaPvzE9ExT
NofiS63GSMgZoGA0dI3dvoA/9IW28rrw4x6a/5Tvjev7d9zwPf6CiDInMJWnm9XLkFpCt/mdvEDb
UJTyjGg0jUI+loftPrnlofzQ2ZtUFMyxSRymyYjCIEcx92fWp7MQRM0odDja2/YTPyUsdnCcjsoW
EjzrtHLzKC+/CV8gR1yfu11Ptvj74JR/Cpv3vSKaOZjU7F4axu9VlFcNKfXfsvEFyObXCy+rVWiM
da4Ch11w7k+HZK/gJwWHyrGd3w27eNRbfwRg7a/l0k1rH5gv3TvBv5sr7PzutHdxe8B/IqN8Z4x7
17m6QzNMSDgp1XggOxt3mSk2GGGiwU5OGedAZidArGRj1xv/fVaGG8fc8WU2CEDOYLt/LeFGzNlK
M05Gk2Wdf1h84nmOPBMSOG3xAufb9v9r9d2kZGp4k/gvKdsc0K+hW7xEZbalKulgyFEqwHhr1xii
TJTWhCGqGLCQSx9Du0YAKqPcUsHeXZaZnN244RPJdJ9IK1SFOZZrdA625LDT9J2nPLm5Spmg5tzn
8jsEXOdwC8L4D7tTZfWcis5+X3rJW749+fJ/PAMigm4aGYLYZHCJJ3ydJIN3lFjEyTlSDZ6X6RLo
AGgAzFQeiYDPSqJLEuk5IrYtFE7eJBtv4K+w3EQbONf9n1sIHeH10TqAXmAXCUwKG1gAN1CB5QjZ
cwqr5f4cTzDK6ptI1jApdr5o54jshxwWdNJV2SKQ8Ki0hfgCZRWid6XzmyW42zfzG1dq6SkR2uBu
qPVM2ts0oNcp5n1JjR0KNUm73/2JxuJFW1We5DQ3dUHdt1zkgGSpI0RihGgC+M1qU/32q0sSBmT7
uMbq/0xUOfVDj5SWvjFoaRqXwmqXbEaX+TBgPCtIKyOQIB84vCenZ7n0yTZwKFGRl1lt60GyleCv
1HyZj1pfShkzpUVGOCJOb0sM2ons42D7tA7+OZI+3I1gXGr5UZlRxFPZ9qUN2K5SiqqbjTbIaBtr
hAyqyfjs5vCvQYNh/TsC+ixwrpMkHgb/pSkVU0QXg1FsSzdlYCPDexNCwVgOiVTcIqgJI4RkW6L0
cepVKAJUTNnKEQ/PdstwvQZeS9Rld56gxo1cBdLOBWnYaSon53AB1xLYbutIPJDY5IqYlTneboRj
fF/C6YDx7ZOYMahiFINrI5LRLBJSi1/NfHCewTNavuvtKTG6KlHn6G5kzHJCLsn8schydxugntEn
m3GVglWK+5GrgPqjvhkoIIDhZ3n6j8pf8oNxaWznGLYV/N8BOG1hhEYHInd16MPHoWxV3KPNFyyK
uDO9Umn0ZJc3q9V0fAIQdb4Tws91PMagkLQjjWN1SfY5S428uo2TUwd0Yfmyb+H/qGvGWgXEOmLS
DquDr4V9NDd+qLJA+6t67zbPg2+WVO1x3uQ3VOJMGmjaRGoHuRCSJaIPyHoox20EZqkzLIsSAn0Q
TnjOtFCF9f9RYtz8AJqj6xxYQ11gvn0YezvhVgWjos1PlUVTmaEydaEpKhoMKrT2Fjxh8Gb/YuXz
UR/4ykeOGtIIn1hthU4YF/DzKfKlzaWHitkXv6IRJBh0PG+5DYR9vwUq521jIx2Txj5Z6ASyQHXT
o7BudkS6gO3LnSAOQl5Bbmgmm34UydRXkS+7yYW3NzRMXVmLT4kWJSmWePu4uBmb8IGndPUmzJBs
gU5I1E4X0IN2u/yfHs/SVvLn8sOX8Gwa9h+j3i+VuvHLwwPK0dfsheWaesCIQTJ9HVcKLzH0LMPZ
19SPOMsNApvhG4SO3/kjwRRf5IxpwvldWxHeJlC6NkM5ByKk65fvIWOGNPTQzajCUKpYKxxvQil5
bNTstplRgDSTN5iPirAlBu14s7KUNM7s9zeyjCWecmYbm1i+7u0GVxgwdBLQMDVTSRuwYl4JQfxZ
qxXGR9e0SZUgvF+I35jwOUPuQ5+AieRPASF/Qi1xReFtqLzqA37CMRgEbn6kO5L043xLYgF6O+OT
yLlKWT/sMNDwvID4MjDOybiD4Hv3HTHXe5iR3bVLXQTijuNf4Qi4KqyLoAnkmWYc0HoTPoSjw9Dy
gwjRehOHDUT4KxQXS6he0TbAJJIykIWT7OaKlPbJcPlWn7dUvnH6SVopoUEM1vTJHwcaHNKlPuR5
Fd9M0wriiG8ErUl9FfsQxB8gsp0nNK++X0bZdtg9ee8UwLYfeCA02o7z38NMUBbezkEm/OezSzXI
XBfI7H4uBhMu4sNm/f7AcbpiVsDF2aJo3lWD35mWpUxQhXmDSiohYouO9Vy8iKW3lcXCBmaR1knO
DE0kVzxsB66PwQBQ7A7ATk89+yuX07SHqN/b2jC4l809QR7ekkr4G1+SY31ko1ujRcpDvWdKjEXD
bI9lvyoYCaez4WRjOFvlO8qQ7k7uhFblLujfBEH8iX4dEiiCItkE6gFK4qwb/Pr+yg/ZdU7Zafp2
vfN7uz3aARAMfDn4bZGTwg0VBJ1pXrSCAcr9+5xGkPKhC2CO2f2mwOod10bhEfaAhNCmlrSWQjGp
owYwe1hTP5JUoscvrbdDyYnYMhlfZU/XQEpcWPI1cfOqlcXDY1b3DifxgM4X9vL94pG4ueL8fr8V
v1IDw497miH7I5zBfUKL2yLbrTSFtiepDbZRY0shbVuZ46zWzlTzaS+PwFLd4RRwjxwgMzlOz7Vc
8IvdYYxg6r/KVxUdYxKGDbCIo5CqVDXsOPPFB6Rf7Wv0+NdsGJZEjQZCYgvmGtmmaomrnieldoPb
Vjk/0I+vfkU6J41opiw7ebBSB2nOUqdEtK+BteqN/rAKQFO3v5QiEr9qE3rrbCfFm392eoUKk3qU
awyU7hsOWMcjNV6Ua7u6hLxP4iefblwLVaRQ05ES+2gAtzzNho/aKFrPy6ZcTE0DY4VxdAkTtQFM
1rNXuFBT+e8D1Nbzr2/O1K27uhff5VT6zNSZwH7YK0ZMO9FlIp0BLlkNpQ4ylJz8PseSGT/6b3H1
+Wf77GuNlXUMBjhFppMxfpvkLLDjoLVXEOWK8D+QAJbf3icKtum46X91Ua9++jm3yHhudAA+WzhQ
zyWBnK+wXi2wZ2mZxEP0BOnNaFtv8+mY056K6JesvmpNMsXC3ATxSyZK2g0CTGMsWC/jVFQTu6YY
VYLs3SUzVvd2LAAf2kn0yuXNz35Zo2pZkkQ/pYzrF2lsRY2XR0FmtVIjKud6pR5/sS3hQke5BnOz
1+E+W7duW13NN4sHMI7EaweDTqtpwU/qccBgif51U0KJqAVd+qm5Et+gppkZRbvUY/pnleMQTCzm
OT+3DcVBFc1yajvx9gqo8pGfsx5RfvZI/7EOvErLKobFAQ4J5rhQexnds1mQ3tR8dcfSLWZ+HQCy
Y2ve8QEoMy2g/zhmTwQJwQe0ch2qRLKrXUlHzMzFzji8ms+/x1VVmK/U8k1gPMF82OPh/0t3Y2v1
EvqR1FPuUK2qx3HiKf9xYErpYmDxNGJ50W2weh61p5xrLEvlfGzIuv9HBIwBVcqqwNqVNfFf38Hn
a1234ycfPFNJJgyV2nuyJd4Kt9zKKT/YnhVqJpgn9gstXri9/Pqb79qippC79CnsP3YRBPdVC/jm
p3cI4nO/uXu2W42Tg1VIOsxv9FQmFbRQg8RH1p0zFMybubXuLrfkUL6GQ6sdVQkLlmesRiApI8HR
PsOAvT2IGXmypR5AUVavdp8q2rxzF80hSgI5MuNecxOxR7BPrtlYMzqPJT6a58PZ07HFQn85aFGr
2IKWPhDLbWwqADoMPxnrRRT/NU+gKUHxWhqVsJJ4M5f7C6k88lOBvNbbm7JxzBScEZmZq16Me6/P
qJVz1TZrbNaEAmIn0TYVWcajLfJFgVR3FrvgPhmFbwCVQf4/zCf/EJ65OXr8TQye4vWRaVWXTpKV
8+QYOrtPYkURi6F+SKyPb7Zler1dHYwcVsZo6/THfIZQlvAOP3+/kdzmuXq2V4akytIgRknbW4bL
EpapDMNTVQrBJS9fItBYNPE2hNX7ro1Fr3avQ5sktl0FFVh9fJbyLrQMrABB/rQnGPV5340alFpq
QHVDQQcdTXEASKAejF/No+tBa63N/Do7A0gWUmqJ4ArhNv3pmGF0KW7Ft97Gm0jKpPRtaTZWTw96
zXl9YURkB6xOsfu4JeI9yxBGd7SDM6d/rY4pn/VvVYrHogucu0OzjnsbO7p04jW7bBs8FnGmd5Qb
fj9sEdKXVeOfF2xFslNfo+UyQ2iys7nvwaBpJffklJ+LlnW9CtPEQjhEz1HMXy0ZhtWJginMcPWm
tUta30QO8C8IaPXaudPFrtHmPzj28a9B6aYB8kgv8H0EnxKYSGO7/o60vuNUrogNbCAHsx16OEf3
+Iw05fCkrnuZWDjd9XZXXpbfYM9qh7/ohDJStWlbfEVnUrR0M3aYdnYRzsME8t/zfNOosrQrdEk0
QH9b6uy+6Z5M8BuqThTeVw7cgQbNts/8k6Sfm9+t00RNH9Ftx2HPYce0Y21eYwRkR95Bwflot2PY
u6kfC+Kz0LVguwUyji566P/laFAsCn1RM2ELJQw1Oj5RNRXCLUzhmjtDCPcXuHNJMQIvVsGloSeX
3T+c42Yi+RVMcCO0QnDJhX73QDup1L0tMjAfGiDmrsZgX/EeiSqLqT4Hauk6qFIAZqhDlxxMiDdj
SApGgS0xDOkLrwZ3tJAQhP/zTR23FTYpc5mpYhjxlG0bXgcRssa7KTR3T+kmD97isOww31EGKtsu
m1hlBfmh/Oy5RZt3u3/sSd7wmUZSZy9O9YMRe25tR/CbELeSuXLcVeiVpIXkWCluIQKifZ3bbgIY
gtsiUhsFihDc9RlCZ3VtKSjIs7glf+L5cHFutfJntIIs0TNmrmv6p7+NYFiEuKrVWbM28awMM/7N
Zwas+pbvMB5rrjSXtpwMlKm6MoSMTVU5KPMidmAA12LKOk3gprCZwLvOh1p73vNYnHqGLGdu79eV
0F+7bGnjEOI+zOtd574hV5bg0aQeJxS8adlCVJMspDN6VAWiGuqViwYj++OsRXA/AHOSNfVZ59Eg
WaSeLkysatUOUJevDY20egf8t5eWch/g2FakeeGxqdyvAzMfDQnY+PIwqZciBLeD7H2F2bYn9ZRK
iCaM+IpOvR0If5rVkfAElui9SD88GyCmi2lnbGItPTHBkvDHvYiCQkihgtCjln4eWhMPJP74Dw/z
t+2l/XEEZlL2RPHotbRR0MCvBJt38xfQwE9kHIHxLdahc21ZROe8rELH6ElIZeL03LdX8jIlkG0x
iV3Vy6QNHOIpGNTw9ON0103t++Axz73czPnNu1ihNL28IfqgN60wtHljGH+WXcCyP8Z2hJfdbRqc
El56eiCdW9AJEzPAWFJlgrPgUTROYVi6wXFfPVaQpKWS2dQJI2aPwibriq1WjVSAmehtWJhaFi+U
OO9EJYJf4pkiH4JLiqPOB+VK6Vy6LqJJgHYIbhn9uPuL2gV/v6KxWsyUmyLUuGWtXC958S2pV//a
1pbUWXvkgvOUKi8ga9+axLxcvCicEabGaYPBnaECQSnXbMQqSedWp5V32UccWL3pkp/rnRubc5va
KMKHGlBPticY9eDFYxzgxV5jCrV7s45wzAmZ/o9+NF2bF5r1YnntVx89ZxZ8WDIQd23kYNeEGz3a
+Rxa2O7RdFOP8qCAM7y+W6aAaxDRXGnrOzciRNiyGPD/3CO3IwAiJFXPftodBjHPbOR6zd/ISHxV
Tbvvk47ci3C+fRMrVceR9fNAEw83ewzg7r1YNbhsapDu1ja5rW2YHL6rjdJQ3dITzk5TIk355VPV
DyW0xerZkOIn+zWDV08ptgyM0nCjcQGUu6JyqWz7XpOL4RspOQ17YPcdghIjF13NoaNk+PP1Yb+X
WD25Aowp9KghnL7og4VVni0Bpu9FA51wx90P3W2SlLVWcX5CjXPollxlN9mRA8HQzhHPR/XerWjP
AOVjYpIgocyXUaqdE4cKbVQhp+pHElf6bZzGJAayQ+uVSIUz/uoV3RL0Quazrsm0C/GNbEiid1bO
7j4ms8WOlwSytI79fBViO4ZBsECIB6QfLIu90dHBB//ejpx57BOtOtfg6oYREaOAgb15SRuVLRmu
d0HkRxCUaEjT4K3dvywhYC9CK3bxgJ4B294hf/kUPbkuefrBIBZH5ztmL+Fzt4oYHfcyeMluwrgJ
SKI9mq/zyOdvaUANDbRViFFHROLr7kBT32djKnNwgJ962mV+asezQ9GHBZKYwQ6NYbcl0Kc5DuKV
7PqSLIQ8M9GHNbUKTkMsMC3r3tN02e8c3L0AOk9lnMRoyB/TCG3Ao+vDemJkoHfdwCUEIPEfhvpm
q2IFnIRuGz7Svn0nYeBniImFQkoAeyYa14Npsjm/Kt3UfMRvh919adE/lGxNYkBD/QJVUEkxYTro
ZgQGAKwObgeqcnorVttT11lATpUnnXx9Y/MkT297ND6CNa0gI2xqdo+eG2Jg68M1n7ibSxIXNY4r
m81v4Ofd4JqZwLPbtvuZsRrjbVkkRyvGhiUDW6gc4yQYcr9bbixPNGAi1c4nMm85P57p6jkewyaH
wJHY6Y5NVEmDLWDd1JaR6TMDLc5Z3gJDsOB7ZMg9I1meCSV49vgGxR/NSk+xYf8bSUUQSW8AS8bF
uXZeWrgMkJpEE4ZhwSjvRv+hhj6DDoTQ8Ia3HoUpYWEqPtJwINnPrlSZ2SxmxsA/AK94cho4Do/n
Gax1OUT2JQKN7ElrZq+sVbxw//iLMnFhiYYr0/eDUuNei/DoMEYQJSgENqaxVS8DNvKKfpFS8uJB
qp1M3Nwjs+Xp/ag/Uj0mN0M51xBvKY68UUoeP/dAworzbySrR+VGZPIb4ua4sXLmV6aCKERIbGlW
xX6Py50x8vOgJChJW/2Xx3/GU5y1HN9sTduWC/g6o2Eilj3+JvkSWWT/vDeQB1PXDVKY0TpFAbZJ
TJz6DEXVAPFbdNsPol0L2d3tJlKEq/oTSgN8BXlcu0q38jYGo6PN0DFZBQ3898h4s/leZtdPg/Re
hk9tjam6CToI898c5W+JCSlYsXu6FHSEzvkfjuFtObmy0agsPs6rYHCY9yTtd6DWyJJyLH2rRsqt
LbypxcimG4DhDsb7EKTgRAPoYsX1RvLxPaqlef5CcT2MO+VWnN3dXLfrc9AhBZCIQtO3Znk/qs0M
koT6QC8NStjz3CZbZWBJbHChD71aaqo5fmn6YZPQ+lGiaj+0PMe2KQNCGABRLHztc3NB1h1zul1I
Z0xytXewa92rX7BrENEv64Pu87+a8OnzNXSxGtLhroKgaNveRfEeuYm88LL8kN+ToepQSE1PYs6b
81oox2uNLrd+W00BHNK1XbvNXSHiSJz7A4Iqhsa+6VeHi17R29UbETVPcHYG4WhBEExrZqmwu8fj
AiM0YcnXn63x2Jm1yn/AVQO4YlM5RS3UNJHLJwnNnGRXHIBGSResXG0gI8+iJ7cn4unXZMFTgYK+
RiX63eVdQy0Lf8QFTUajnZpyNHaFMLVUKginemzM0ZiCaF/kYZ94KmAe7uA32L8WCkrJzKwiigXy
fSJYsHf70fHIkbPcXO9WUlKHS6yA6HKCQWGBVMbfGdtkXtG9bLsqFBrrRa5+E2zL75y3Dh6AgVx0
866jdzZQKt8/ixohzmSmMvVsiJnGLlszbnSLYRQj6MLS2iGCUOqWLQQQc5ZDZtw6QWi3edtBx/WG
hbUvm9Ui3DKbCyCkri5j3nNwY2ETkb3rYfu3Q4MI21QD2O0lj0uBBjU2kneghGghiLGi+X7aACYM
KRdqEuG6sBRBYfDzdvK7/XCHRSlYsRf+N11KwsttTwnWm3UV5uL+1zR/PQyneLvwoQKiXcg549RW
qVQdB9dj+MkWECrJ2gcMDoRmIJBJLLP31a/HnxbPwo25HhKtzZccyMEU9L57gK5defmClIuROXTa
K0QmZhd7JTNFJgOZ5VAtF3Myj+euslr+iw7vQjcZgX3z6wyfOSSy48hK1HGbiUFBlx3sMcQU64vn
ZUB0jJjTDBCVy5LhyH5MlH9cl0li5Br10xrnrHP0YmSUCl030eXHKgncLVrTilTV0SmAEhUI47Hs
H61DepjfMJ4JIjMrLJcgXNWbQJKpmXNDnmiAF5G5CxjLBRyKMXq3QqDEMtODz+b1rK0/sOBAO/1R
nU6WqUmU6Dr5JHmFoZqRHLKJ5kBlEOMAuJlkkzpL2x+n+2vrFiwgqxRYTSti2zI5JzyePZhgZq8d
A+5QdokHKNVjFCPWQjbwB+TnMrIdIWF5WRRUyNT0+ZWEASz7t2Dn18n1q+uKbmE6VbpbbtSqeh+w
Ya2/YWSLyltheop0gRImm/KfO2BW38t9Dmhwg42UCvW95SmGNfmCViamSJ7KnpsKFWg/UgpBu3Wk
+rW0cmTwPcaIkS/CuAHEv0U6GNEKyw5aZUSQZ4s3YSAMd7dynZ39XuooWDJcYfVQZ9bcGLKz5oYx
30tm9AisGQi0QPuYqRmCv145efTQniwUeJ0Rx7p7oV4A0oTooRWyuVUzYzZczzIM/XyGaGaDpZDI
2nyKiQQaiPIyGL9Gm3MnY7keE+s2FHTjGQxS2XsktdmYYPq/ZjjWsqmYQDDxvyKSZ3CqPMwmmLTi
cvev9dIXuYdctrbB6C7uFG6ZxH7Ya5i1jMxRQoq0d2Qt9qppPaRrp1uHm0csu3XqcZ+qIolFlVmz
VdgzSfIb0C2NFFAsOlBOFcGJz6/moXbE4iz62/e8t921/Bk7SqPtqIArQqhinBwA8vYbSXmlIy42
ryQ2JaDhYIZ2aGRAsBw+wf+iQg3SuCnFehLk5bGIgHoEn/9f+6rqOJfuA5knYNkE0gpYRkLlNkEf
VvCsjA2ucyRxLS6wp+RXX+5YXwO0oQIidYyTZ9M32ntpM/8xZoclCaRle65EZIRqcsonfoBoCRac
w0Ml9T0il5HTlvkm7c/69OJX4Eb6L4vFOecN+Pq9sQngZOwegdaYnweizhHkweLSq/UEPEcdLZBm
fPFxIE2ZLe/oQCE7Y4zQcOmHbf+KTpDrG/7plDAMKDbpTUH3CSRZLXKBCBMtZ4J6COR5ec+Blo4V
3tPPlcHqW8mDd9+32v7NEWtfRrSpb38ne9lWhX3P5EC0LV9P++SPd1nciu2dFvdKKXAQweoWglKp
sEkNMD3dNL3xJkndQTgHq8fJr+h3dpUI40WylxzG8i8U36CfpxrMS7BtWxoB1fouLWgsw79vXhEb
iFgePE8pDW+9gd0w1lUFCGvJIxRr8dIKNbFYdUrrlokwAOSVLSR+lOFy33Z69xn2960ybh9svKk5
/qHS5vLqiOlmP2z/DkOAgTxYuFMWXTzLYWQSWDH5QO8eXzPUgic37QJbkbavQ/IypfQ7e6TFNlS9
a6aJjkfcWvvIDgVkXFB8XDfgVdwIy1eLWvOOR27fa1OzQQVktVk2ezKTpzuUs3I9Y1qripvm80GB
XKqSw73uwBQ7C0h8DrY4Vrg2qKxOzXMIGsjhAwgEwxq7F6LzTSLnPYs2D150jSREI+v2bq8If6Bs
GsGZaCoxFpEOPx9lFwZTV3hATvNAtjSzrAR2VDq3UaaPU9cEFzfrYcjyHAb7OSRnnP5gpcA3vrXY
JHK7Et1rToulFs8m7HQPL6ttxhBnUeArHn8n+7S2ZEUqo1F4xAorHv+Ok75U8kNb1d9cl9ZmAlpx
Nb5PiRVuTATGuxH6
`protect end_protected

