

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kIepFJ6jqif2Z6hQCi7T8MYfP+LI0sdmG8lsu5wSq/AxCNeKlihKZ8YcPR74jmxy7mTgHLdfZrbq
A2Kyc+YhPQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XFGKoj5BxP9RdaEXlRCt73HCgihFExQ8sMgDBn06/Q8b+F1zZ6I5mx/jTlR1yk490EZba3ynyP4t
5/4eeeR+5y8yDRk7Vej23u23a8QnLAapPu3MH6JOMoR9TcRmUxwU7GrGZ0xJwWqDQ59+WH9II+M5
qp1wcwmTlT6zAzv3vFs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YjHf6DWoJJLnLxoBfsKiAoXggXY8GOk1aAXMosUj0I5yJ8xXOJz0ATMRRzdR0fmoMiSkVNyATyIO
0CYY5VIsQ2e5bWA/TgGTgc2FfxCtlbwVcSUyFqhLuxtdGqvK+mx+jENCHlWLLVc3DPSq9ZOgBukP
sZilCpMmOOnh0743pp98LzW+BB+BMeSOD+BfFPe2J+aLBM9wUmA1IliwY6yG1pPwSvw83zcip1E5
iXQG7LgPBjBIxpBUhpr1Os24+Vr3O0bfhJm9I54YFVRjpmdDgd7BZn3JBabE5gBMXOrkH66/uvey
7bHaF+o0Y15GX8VxEGDww4Z+sWiuJ5N2CcKd1w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SRGphz0voa0co2qA79Q8Z0RPvTHJboTdEbP9zDkDmblZIM158XGWXVBFdW7hTxDKQ6sbYAkoBg8g
brd2dGcWbk7t62ITmWohVgX44w3tzjPRyZ2TCmoBbS5DtjtOExDq+TjuNCnAlkXOc3rKq1E9idTK
CLWjzBpNlsgou2FMTFQj24/UHn1/wzcIfxVe4QklIMWngr/cCRCZQnVWO7yXolY2h8wJtbVCPTCS
9VCpj+fMyLF/fW7P/hxsuw6i7WYBJKl2AQ13A6vXee57rb4ZpKwd8wMu3XZxfBTe/uXe+TKQZnM5
bSVr0GM14tYIULhUK8kYgzAFzXegBS0CUyN+kA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oU8jgelAr4yOf66g7pWNXMjQWD76kL38hwIQKewr+Ssy9GGSk0ttJbvsslwxIvk360eJ3s2tuTlF
vWUwBMH6Vv68S+oLWMqGUzC8rdnXi99SqxMvzdt7Tlc5ALZHTmBy81CVh8s3ZEZfmiQH1fE1xu8f
grokkMdXe4jhvLiHQ8EIUTFpFDtzSkK1x+moiCcoZOvESw2OsdpELt2QGwGEPEcs0xJ7xalEd3+R
J9VsahhRHKz5mQzYmFjngrRdr8UidlsZezhckSsKXZhWbxy/oMP4luzcg2UdHaSlsV5pGuT0IE+n
NgyXJFKH0pFFTcE4PzMOQFcrflNkxgOj5VygTA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K+SxpYPtX7YIYtuW2uIYAtEFYn3BIXrQyoxQi6OajY2BmZaNtrj/Zg3U9vsrPOwttAWzzzpmu3LB
lU/gE+8e6ISjRfrDyKvPhLAnHBYsEjs+QL6xETVfM1dLq+LypJ/ssq7sznHoHOSh668jBqaKZkei
ar/4OvcYNgPTbhjbm5Q=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L8bb8Fo/GJpLVKff0w0u/ZciZ3RdVcZRaygP2Y286r9eiCpUFSvALLGKcRIgVrrNndvNjZLiq+Tq
wkJleJ8RD+xIS+Y7aT6TqEX9FyViL9xjMwkdq/se5eRjhl+kMOuNlk0xKKRhqiEZMquClALtygBP
RKw0Q777WsCkQ7X7a6n4PHP+8graKR7DRp5OTQVL9BF8jeWxQFHdwl28CPQvmncAosxrkxX9Glju
/5DCrcLDqFQuadZE0FVCJGbmnURleugEkNX+PFIwgW/hDiPvfsAuYxLVYJDbXDt4dFINKeZZDE1M
8tQKruEt8x9FUJkxiqceCeCmKgbJtJX0XXw2ow==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DOFx1DDxk3qeWE2T5Az0ZiWpzeNbgcXYX/DDPD5JXspRYUMv4Ws0IBS9bXX2Q5z/9ve7LsurUlyE
gTayjUOM3u1YibI/h5ZivMyyg+QW4AueYYAtrVi8Ur7PTqaieP+6mQFYZO/eM481TDgsoEQE7byN
6bjzuXmQtbz6tBgkULcpJvfN0kXkWSaWOJQuid5j3Y+bCj7oAGM0iv12H6YoAiWCfbAm6B0aNH4r
lEaqcqoUNv/bcznqZpH1tKWMxDajmCXgMCE1DSl1R/k7ViAASrXS7uei4l0NAcao0+6dSrDhjDpt
o+8/J2A+FhbC3pud69+tFqRwYMUq6tLgL3eyQA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175312)
`protect data_block
HKXyhSGw+YYjIRYluRcpW94LjY2cCxeOgX66FU4sxmh9DeCC2g1scO6rv9eVJmaPMBrydFId2FIg
PLa3dB5aMRie06yoGFsvlQOY77vp0fPu72JY6pFECcObYe6leFj1JlieB6BrSxF6lv3PB0xyW0c0
qpHO8h6PP9YKmxZEAefrrMsDj2vb74RPZmUw+sO/R2WcFpIQie42qg1YoLkqt2a2PvY+bFaTrasG
dPmQ8vzNCRYZRLOA768SzYFsEap2kNvEIaQXNzbOfhnNPULYYH6g/blmT+poG9ucbD41RN6aytQ/
0H58+S1Nt01bRKFbMvYAzFzexdrzA55AfQSXL3VYr2jbok+5kIt1F4qhOeBgGjtNxlkvxAumtX4l
y3r0zgbCbB1JOzXDVZwguC6hCtKpnYapbTKSuewSRsYczs/O6QMLCBsfIIIXsMqEtNVOGQyr7GHZ
ZuCL3OZp36r4CIbRrrGQgrZzFCrXuXfiLT7BglsK+zxM99HoNVWRvaaZkwnUWY/CqEnoa70jnlvv
gW2yG3VeYW8xuBZhD0BmZDu60mbh0ebSdYt+U/cTwgWmb3WdFVjzO/AWgeWtt9rrUjQHSMWI4OfR
PK5t3Zms5CDUv+hRAXBKOE8ewd/DkXj3K7TiVcQPGeEMThyBPAV4BsHSFLagHQuQMpjNoqpIJa8s
TPSYHJfYuvxZh+PWA6LkHExKTi7Fb/ZuwrqFoKlnQSp35Umg/wuA6+fDy8i5/W3qpwQXeMd5kPCr
UoSIO4o3SJKas/uf0Hdno1Xbax6JNhZYLSRdbkODotk/fXY+zJOHO6IKzQoE5QlGbfCvnQKzZDZX
feHFrVrE3K7/1Q+FlLoHWLByOaSFpXGvyPPWi4/52j0wJwduaSlGGhpfEjjNGiPRA1B3qzGv3i0l
iiMYizO4sncaGG7z1CbRMoV1O7nxq3L8SH07e2n1C4jviwPuoeeuUG5DLqLl8Owf8sygnWxZoJNQ
BhgyabNGvBYFw6j8n5f9onLFrWd22vzI1Sa9ULPe/MsxYKyeAytErzYRv66AYOFEqR580gRGsnVh
pljDNpzG2S9+yR5RLder0E9eR01KA+Bl/OZE57+E3BKUxThjj9+4AMOvMQUCo9vLjdkH3bWIjrt9
wT6NXSi4KnQXkFwKdzk9+Z6TcNB7i+YvZhR7k14r8DyjpI1tyoB1Orv+iVS+bvFaaYJ+Ovc6CTw5
G5rq8xIt2yKYgYc4rAlpUvXpR1cuj04IHo3bld3TMWUA0TQLXuk07H8l14qaKxrc6U36GvS7VmfB
i2F5P3/rcbrAqW4bARaH9zG19FuTAEJMbUCtMifHLYQsbavitZ2ohpi2QQFaRk0reu6YGpETgtT/
t+paDEuD4RZkL7eJpIvu++pcWgwSGYxSVhgIsl2gJSEVD1eeCxjram9hz89ZqL+zMsbvyb+0SJ6r
0dsydVXQ9HHvc73/hCT8j0nT7Q8rOy7mC+N48KJhhmlHF6QNW/XAvAM7C6I7BcRLKkcA9n1gWbnu
dinsqZBqAD3zoaokdqXXQT0yDn9EoaZDOR/F3lUl+scr4m+Tp5W1f/v3ntqEKCNfVbiTa/Vtyln7
RC4mcfADkA1MFN1MM7VjEP/6syKKvSKTxfOTzSGUAIiFQVo8xTrjqRxq6mKXAfitehcS85gb+VA2
V/SsYJyHNPyXW4/S/AemvYuvxRUaaZ5Wv7uypcSQEbdQXxVqKjbAJPQq0wCCwzudGsBREqjpHV2O
AHdc5wjGGVSNYOwn/GBkzQBd0R2yZ8pACxGus4uQpbplMvvgO9IwMatrslWiJjAPDYAP2GNjFowA
SH1+OG9PI/er/HgVpUjdSRSWz5ACsiE/bNuncgM+PnANHHh3eHA5rJDzNsUDeY0JKIhVvu4f23Aa
R0gNjM7YY8VVkPRg/Vzh7hxJdfVY/B/wRekODoXFummINa7YSNMv9uliDrwqQCoMKQCDo8RgFbKl
96qPto5LKUYYUUGMk/qLlhDEH1h0JgfkmzE1ucXV+ISRAkPhtAfKuCPjwDQYlMnJMKtUwQ216xyz
v/xS5F1DRImQphviGEAg6NAgb2iYNEK848wiealU7Ha9kGNq+HGlsCpuIy0J0mzXB8zBpy6kgA2U
H8dyUNRgCPU3NEPYN7d71N03ddG/0Ml9c/+glD5BsuakKkCD96qyjqb9HMBqnoPep+ATF8UEKCrB
ByqUzk0n7dgBSq+Oq9Twx8e2Y5+vm+Xpgp3339JdEpFe0xnJVR+x20XBBAIM7f1zvHSgsJwqKxUy
1NDzhWqnhfv+RmHpwnQZMmwM2wXh5SqwmpFZl13jblx2QrtJ3nSR9of90Ap4GeDLEotwayThDLa8
i7qCXMVAwPTPgrsGt4Si0NtLEjhphQkhWU6j++ZQZLAoIyuG/VZgvrDRzwO/eZJtvLifTXVV+dk/
XU6OvbMv7WGKYy1yamB9O/ZRp8lQT8PBZK8ZvgEJKCTUjjwDqSUVGBv53x3QxvgmuNx4IFhbpbvw
yTYrj+78RJIdwZGke4Jpvxj76Yx8ANh638agcoQ25wMc5PEG3kJM62yZYezqDxITGiSA35Dn1kES
3HH+NTpb0sZEAk2qAaW0G73zoFHIxwdPr8sX6GnUc/wfA4PYxf+U8HeJTaeOODvpH/XIi0pHp8pb
5Zv0FbHV8wKgyDHPoRIThmxjaQxIeiAemos6acKcMz1CPfbJZNvVPN70WVC9w2KS8nsQuTLWDVKW
Par165xVOb/LA5HfO0w8fxBKWeBuQeQ/DyHe83vcm3E5iBSMrXiSJ6J2a+cMcUTUpwkSjJ9VCbQZ
X8AC4NyZgi7//7S2T1mT2u32n2GiLghyI7ypYu2jNPCU5L+YMj84Yp/pEDvx0h0XMn/HKRIGL5Nm
5fexvBxZTnbr/P3NdJ34VOQwW4Snz24ejaFlSVoYAQDaXhpq5kA0OO88qT+HxYrwwtp+i6JK9ODJ
Yns9jEEolClitfn2Y9f0ZyHgsS9C4EVzwHeRIL0i11cB2rIwRr+P5zQdUB7bgjeup1TaHQ4QsH9Q
wg3K2GPkAhRH08wI3h/oL5ugnQpJyEbOtWlhIgvzKckrqd/YZF6LY5ItN78/CAEKKvoxe9j9Mo2u
rIyTpamuSy+bVIrBzv5qzN7Nusy9sR8b3qB0YRSvwZBgyZVydawEG1+yDU7Ule1rk06+6DE8546n
c3cGR0p+7mPVgNJAUN3Mvtyr1TKHHhkMJBL9uJPuj6UKYZGwv5L25OsI/SiOVF0AfANvSiv+VGxs
n2oBBIju/WDaTJ47JIWbZWtkYSC48U8vUaFGsWnYcy03jVEsvHLgVLG2++6p+dDbnSBox15Z/AKS
CIbPUs3lqOU5r5Oy0ywTj+raUZvRGHwubfu2+MHFXo4NaKQSiwFBYBM1W9Zwhfa6+uUkaQRuSUfV
/Co0OmADXIH9OqeQgE0kpEMUUuOcLqKnOjS3ix7iIMOM3ZHul8VAMYvzQ3roQAHsI/u0PEU7g2v+
f/e/3hdRH9K5JOPNYzehp0bmqY3mxe3iKJ/gMWPWV3vp2UapM0xtB8HjHqnCNH797oKaOauKIDQj
MW+qhyJF3OpdolrVSxhml483LmZdswflX8bRO/YvOBzNJysxaeGtRot2iClPi9bipvw30Vry4bds
kGvDIdCGfAwseof6dBeopZZ799hhpxPnAohA+ryO3+BUVtJPqhIfL2kGwBiTaotIRy1lY5BebDtq
WLegdNRLcet4Hw6miwreVfaMDzhE9PRQqjMV9N/RMiVVBjEwvFNCUJGiB6SoroUI9swgSlN0HGau
EpsNWjQBPRgCBM4GpUo7IZVQ6myDcDUgz82Dcce0YtUsHYnqV29yaNGzeMzD2oew1xdXPaXmCyJR
SuA0B9rnDEMFwgc01FqZWw+xqYNfjmPNcYh6tIekVr6ZVe7JPnQXSLqvgl/zfsT///C1okevcTiK
+keV67mof6zgJTjbL8XEKCXScRkLLUPyIkafYU76n6mxF/UCZ6HJLauEjAiQ+JfVUQBMZ5mK74Wm
w+IPsReUMw60UCtgK3v91DLio3p8LvFSg4uTy//W026cv0NFldZqiV56lcaxNF8RYA0e1mZwlPAP
j//skZseqfOLt3IlIpBTXg9IPShLOYvEwgEmrf0txk3lLH3ZliNJszLYogiG3LmgdMcmtQCjnsJD
VKHnEGwFqaM9zMExIrg5/RZAKAx683z/CVPxLMWhRWbSVcndYR2NNJj2TAwZkaDpQacfh6FgDYV9
VosUxHWhxYVNmuW+/+g0RtATqnKHp9aWlbm47pp/Eo7Lxsfy5Q0/3zHLCIUlJxmA59BRqvahi4dH
t0qcxNADnPRdj9Fr2qBNO8oO2SkmZHrlEn7uqrtwp5zMkkuUuXgeIo8/qXJc9RG8jZAh2W3B+w1Z
l9C+k23nCESFkQ+i5dub4C6WKm4WRVe9yKa6vr4CiF0gvdiXoNjF3FwNI98u15NH/gWNUWD5MBVb
KlbwXsVfv1fo855Mmc05AUkMLCFnUShyUirPC0pqjSwqvD3YsRB6IZK80ddwZxKKxlVVsf31YXsR
VzxQylJ2zRZnxwOWSO0m8dGwuSZUVoBiDR45AC+zuK6bD8auRSwsckoePqZ3OFUYDUXMQVnV9hI/
R/lnEF2edDGV6r5Cug4tMGyDeq6GhlQi+xq7nGTG63AxhjZ292sU8egjC74lXBbpBhnVZLJq65eE
MrIDuBi4JLZ3tBTjh826ZPw3OmNmJ6d3RERxHy5CGHLret0NV8KXXESDrv/8I+2zx2KGJ6jDoEmL
OJ8sw0CI3rd8yY2zF3SisFjRfW7OzFn5hnEP5WSzu0wSmKd36Rkpluv6fCNDDJGJzqIACumw0f6M
uJ3hIbf+0R+/O2YeC9SW6/JhKKIxqgd+Wd5sDV7f+UhfqXdhMyO0jLP8zIU/XxB0/9NfZuDC9GE9
xGOTZ++WZ81mnRpNpcmVAgYjHPInbHQfHsh0J0slQSqzhpd3JFhxcXam2LuR/M/OQMXQ3PIMtFNQ
7NdHZRabaLVV5XRuXSz7w5A6H0xZK59Jko+E9uZHhAqvVWLPQ2mm4S6eNAcvMvxBDvEhWK2maLW+
FhCwA+4Vt9eYsK7vl9feorSphtE1z2pBzBaozXZrvjatRgWk2rbgkG8LEDIIFR57Q1eLuoGLKctK
BYZoFoM7ecfTwIZkQ9e2G0JlYynfmwa5gpxZ87V8/6I7u2Y/d/bHnoo2Yb4QHrzOF0lxEnS/d9KW
JfBofjlvl70SEQ+OkFs+qQtBUu+mlvV+eFreEHc1pei2cEkClNI2MJvROLWWhhklsnUpQnXV3ob/
E1Yjw1Kw48BL2iHj9GWw1JKOauenweiopwgLh7G3L3IlaXjPOW1zQpOV3Xa2tJHrYH3qSpAxA6ey
V7wjhdqRa8XjHFA6bkkqdSfKK3ggyngqG99RHh7sOvhlwG7GrdsKUXNVZHlKkVdYCusxu5s1p297
VwBm424g7DlATqjXx8pj4vfO+fgbbMAt1a6JeWNHkthEP1uC7XFgm43Rb+gwla2skb3SDA4qhJhq
vfFNmjaV8SM7kM3OB9mWYF1wOqE6A2Z6cX/LNShiIUbZuc86Ygzgpvxt5lR8+zovIOlnZfdcU2S9
8VenavSaRKpvymP3Zp5NziKCKMAkwTIRyAvYpe4QYQPfi6X3ex7Qtoi/oCVy2fwhtwmOSKuilb78
mMIgmwXRNH++U79iVDj5nHFEM3mcN2oqxplLx/7uHkzehWn5eTXlw8Fqa9Y0wBUjf4Sd9TmfR80I
S3rLNneuXjS5Q9uXxwrnWbLYnhWlUqrzmGE7NOhOPXfkEk/MeZGKzUG1syJQ2g+A68QOH0Q4Oec6
Xk3ZsMTVVj8NB935vl46hElPOREyzGUZ9QwseoXbwLOtiKIMlmuTfDaFvY8dB6rcfA2GgmB2srgP
KyqMTDtsHJwo0JyJ3wx157Lu0hzEP/yY0bjljP2bnP6/vpJCukkZsrfRv5c0cozdq/pz6p2G1kWT
ceqN5gdQFVYR3qescojXAkZEQHM+Hy2UxcTQbKUG/fHlcciuqDMsIMmnhbeJ4KjdHQ4z55OWY+5q
4Br4wx5sJWdCybG271tdFqk0l72VD4EDHIDWG6ePxoL98Qv4n8AVEERwAgnaQUZI6nXaGWmkB5aV
YgtASqd7Wbw9i5B/QGw3/FsdmP7bwfgVqnL281D+/Hx+/oRvqMrLQEnrB6W6NstBZ4F3JcJxVaX8
98ARHtLnw4L38gbGPlqMtEhIPs4dlbJHOvsYFh3u7FYTwnQSlVh5SsJxQeChIku4PhoNZM2XXfNf
xVte6li+QmNcCa+2LJNNg83cNag7Gy0UD/boXor/Ag4xJ0FI84MtBN/iW9AN5uFzUSVKB3HNVjip
p96hkRLv19EAuaHN9zzFFDPBomvcqGchQq9wg6GK/GftwsFfc3UY/yVlfHXn5JLg0yCTXTocT8S4
OblDcGbXeQJ9q/D1RKxbWU2CSpEqBOt0Y16OI9P7ckFnxHAOCjONEzZ2LdTM+kngNGi4DdCXOb9i
qI7/lX80/qsN6V3abk4PgcdO9P0TcgqnJWZyc90mHU7Cgm0+aqu7surXddgfDHv2L9osBjW3vUL1
n99wQW6dspB5QPS1Ae4PR4l/PZ3shvV9HMAIVHVsYZgdsQWL29WVXbQhLNzNTSaHAqbqrnO3HkDP
SbCrW4mZ2BeBFo+oloFh5g9nsFD8Kz+eCwoIs9Smn/HPz8T2rE3KiP6zdCuLLCcRajAx4BoLYNLC
lt7OaMINhhaKqN2ZLpoqM8hevvNzSQAQLVzb8RoJmlcBneTFxu/g39XkAMyz5GiP52JOlZ8Q+Blw
7cDr6EvvRhC+MlALD4Ag9wgN9vn+z0+W6BBzJC81kDvgi4gPSkQwauvBXOBr3Yjcgmxw3q1F8K41
AeS2juFArmwfbVF/P5adRA385OxgZzEx02tCdcJZYGwpexwkup6pZ8/yqSdBYrnY78tAIpByaUzl
l+w3eBdtWiW9P3OgCltKSfRodn7ykXiyUa8AFhP7blL5nHxWpdh+OJSg7bd6kkb5NoDZSSyc7fC9
nGMASUh60zlSbVeLdTSsS46V2tQuSPV0B0UlVNdfGzCIutniTjc6yOL72J4UXJy/yV1HwKOS8/9M
W31ubzayIFREc22nKH+wYp3jUH33VSxyLBMjA1B4LJFev6TNQKGwZz3wX8Di4FWTdP5ExH5aN95m
KVSMP4oK1WobwzOtNYCqASmkyXvAfZo9o1GzhAefEorZWXZzWFNHE4K3zRo8fpZzLyvtAfQi+vwq
OBvLaoOmTgh+2OXEmjWFMpURlSK1KSj+Cxo8UJ1BMPKOJyaqbaONM0AycrziqoPDf2F5HeI2LXwd
ARTPgY3mPtTn+sbBWwN3Hx/OY/E5aizXyOk8dxjwTCVLlwMQVgjWbffvTHzu6SYBVjicbFzVKo8o
wA+H7ilz+2LH4TyUH6KIu14JwCuCsnrhxJDgWjlARqDweByeA7+DFewnWHloaElItGC6Na6e6n4k
geAvu7twJmDlbcMNmWMlabqrqH1f9WfjrC9lz9iUN+sEYB0DdSgtejT6fqQNRfcPRFGA4/68kPjY
KMxWPtf5kDuTu9sar7n2vyHqglL2Dj+YZZfN4Oz4vigpWtjkYHirAknXQMkAB0lI3CtF1MkQrx1K
/+4P3A29FRNSfAnFwpEOfjVOllfpH+W4JKOG3ImDFfLLDVmDl0oAUabCeuARKQ8qv3hXaN3pVFwi
gjZuE6hX6axqVYVJLzzMqeyEVOA+qflcDIUNGAFD8ybiHBqiYg5s6bSOtrH+WfJSFZ99lF2GEZCr
YQSSmkoijH3it/IUE+270OJ67AOZyXOKfzuivLvy1KdzmtY8tRqIGej7g2kq6ixZ+TehnM1flDQr
+RvL/jqcxr6Z8q/2WRb8vUvfKuN/qmbjxFMGzVEw4+gl/74LHpLAiuE9XhRcCHbzxqvDl7fSu64L
EzHjUMVwmGfN4XBIMpXaHbGr4bKvb79L2RrVmVSaUAHx8eQ8GGqtQlw253rLFwq3E8i6dYcBy9gf
QiiwAvrwfmqIGLBiMwZBGKpOrslKVCt9pQmqLqyTnyoVm77rQ3YXzZpNzJK2GKZG5ks1VeeMab47
WzMPYdih5pbQQGSRAKlj3LRPPpIeeT3Nr/ha68veIzUzKXIyguvLdOtYbHgSck3giQoT1aw6Fvbm
p+vj1CnivAToN0iK8M6msJUYUG/eZyvDdzLKrP03Hsc54O1OnflWhuGx5s72OkEzVtyhxOhVCk/A
/Ix0GvkchZYOa27+AajzSHAlrQWtVm364Hw20y065GsSkLOCnQZrceXP27/1nbuPs46In/70zjQa
i32/poNBTOwqWy7NvNaG7GdLDCelGY4VIf0Hj9IKInEmHZHlVtleCpB6AmHhiKVsMfHxqpMZ7ESj
u/meNUtBzsWM3QVP56/NEYyZftF4m9MWXXD/piG6SpaSVx1UBZPLC9Swx6JS5Z1Ul97N4SxnFVUY
EWws6IvqFF+S3DmpOF81dN45DzPcqd84d091FX3HaoE28AyvJdm3Xjl+H00dq/KEU1ZYNh0UMcib
Md6kZu9mgSCWqMKlRWuyfbx8JktiryXCa6Ur7Sl3MB/vjutgf9ZevfIXSRFsWfwE1220aMXuPbzx
XBm8FpGPcnqqCligsYM4p1zy6KzU4KT6LFhWCTXwoxAWW99fIsgoq609JJ5MMyhyZFL5xHiq4ndW
41skFP29ZzXnN0c9CDB7lQd67PstmB1kc/oTuOkN4mF8Yt/eMVxi1QlT9FEsMt6wAHus2rGz98j2
r/8WJ2OKww97okVHZhr0GI6IBdLYEGt3lUdvF9HILmHoXER1qsf0CJ3PP0ae1H/V2mAwVDe+Zk2Z
q63TFLNzqZWKnc2pwCi4gsEQ7egFk32Gza8NPzHHaKSwUR7u9tGV10mA8QlPrH1Z2L+LVyUZeHyp
ej1gNWMDEa0EGPIcqu4A4qM0sxe3p2oX1UTJ5IR/Ff6h0ATZIOziW9am0nK48dgt4WCLdb5i2e1s
dElrFKzDLMZIFNx5k/YvaAWnWQQOQQrOYdHUBvOrUWElSnFn9WV6JhArP45VETHqnZfxvH/T4bDH
573SZs3T2zbMfvjbip+zgEVLNIgAxyeyGaYQjVwfW54c8dDf45U3i+Q5HkCc1Vykn4EvmrT7N4PE
96iOgB0ZXQh/xrlumNl/4XUbBCxw5+OKzSBPOQrj2x/hXr6nzJdeGnyW86iIarpmLgw82XgQT9Jq
oOHZ0WJB8ZbVhR0QCMZ58+C3coGrmQwOoNAUOGC8opQjEeio8VyggG+FngyRa3akYHo0jHujL/ym
UN8qhgQZnQOHtGgLuakVaD6gYav0jbu3cHg5S0hWeLSK8e+ZAjOf3iKzYk9b988XIqHvknfdoXlV
/p4ChecjpuSp5E/sxFStueopb3nMhE5oAcJA+pFbZRy8OyTQ7JS4a3ZNvYPdWptTOoeUcetOgpMQ
Rn094BT7VgQtsSVxUY40eFud3huoDoiYd2/IL+MDLaJXLK1EYbg4f/4K35rucfyF6vVw1+kTNrXG
Ac/OWes8rbu/B36vrY1WxJwAJodJU0RRnsotdd1UF9/R3aKkto53VI+lZ1Df4H9dO6QPUho6mPPL
n9NqUu3kSVsbg19KjBSeUNVTsAaMenR25hqk4Zw4HruNFmw1Wp4IbxXKEFwIUsks6u4naWcKgq6f
E1CnTmnPLWdLAIZUUGQi8u2THj8Zb0oihB7oY1KFf0XOvYFkV2FJi839qId7g4kdZRHZJZo4IJG5
7ktg1RzzkyToD6Ec7zuMoM7V3dTi2FnHFFVlXdQQHa1pjp7Cjy95Km75SJRGZiKvwFGQ7l/qKnsw
c016495ZOTU3xzw8+O60twjmSCWgd+1lXC3xyM6CzGmzfP5rp0JUnNTYJ6UCXqpEDfM0UsWWKtMf
ggTd1OHyzn9i/0CQoHSkNF5AYvh/RN9R6GID+nXcS/A9MFEreqlq80/1z2z5h0SD9h4lBL06TA9B
RVqDtiQzJsoZnIc5MDlH6tYEchCh69yW6/B6UbUqeyL6Sx+r7pVIG9NBU/Dk0Ie8GLvK8JUmG5dw
hXXtrckYT7pxleuDTe8pKWIR1vWJSajn1zjv6JX2PlRnnb6iQozmZY/H4QIFDN1OT7hd+uQLQO/3
n0umt7Ls3O2PY/8iko7UKZu2s5JbSyEBdltfdDdmJmuiCjNjKcvWzwVMaF/Nc9QzqvIZiXbeMr5J
vz2SVMYzRCudOGXQ7rKDix+QuB0y0LXj58RXwHGC/4Ail7RMnIld5pPFU1uwBWhT8dYgH6oufDob
RgjkBp7/cUb0xBJuZt6M6zTtnI33TDdXcbevFaFNVeTj8JMC9LcjhZfuooadfFXpWhhdPjD7qJLC
w/a2ELZoHnm9ISk1GG+DzID+VblWPNh+JTVOIZfIcQ4Z7/sWxRmrm9IXNdQnIj6JMe6t2MkL3HxL
ozxM+v7SQyOAzp/oRe05gaoCo7CiXgRbLbmNaFHX0RURDfaIRj0WU0sUyNtm2OIOZtABD9HGPc4O
J6wT3W4V17XHw/V73wA74bQ9Wxjgb2pempJI+Dfn7wKdcpuAAT8Ff1iY5bTh3JDuwQyiIpqCEYyE
X1zXL15+HXH1HFz5KQmVPUID0li/edfjgllOSIvXQnzz3seU+gDG5OnxW5BhGO4NIcOcbVR9pwqV
Rb0GpuAngUPhj80nKFpCWXESzQ+ZwHi3lXzWoK0Q+bsZyiT89DwryExPNIxNmZjLksFVuStnCcF1
YeuDBgNyAoRHPvXv9V3p610PimhfM4Yd0t7eyO8zFCs7OMRjLJ4msOCEi2PzVpERN8iUsHl4k7oG
jmZOgQmTD5PN3EzW5jc7NSHlTgCQp75cfbPI/MtDMXsULQmY95rZFrjZb/yiJ4rSAQ4wCuIbiJmT
h+kWNszNaH3R/OpNTIGvhZtdHd4Lgdsj/rmsg+bNcMc+dPdHjwYdmp5jeEje/BxExtlg2VAJuN5j
u0pgFH7Apo4W6ZtKC/AIOgz/MnGm+Lp0SoafMqS46Ey2hdsblVQBcgcqCIqncexL0oFbeewB49b3
fA4BmabLTTUmHMiaLFPHBEORwCABeS4XsyrGQxgKiF5qyynmMVveV1rpoHHrrzt0Sjh2lORnfIn7
6Z5IcSDD9NBlQlKI8AQ6vRmNo2/9T6ng+sH59f43f+hhofU8tWQ9SIAg3QP4NgAlGY2D/WKE8dJf
H6aOl1BgQxfe22Kbz0kUv6CnKxBT4FrWSCFnwI7yjOLMBcjAMOKELCMu413ND+3huMdNWVjKmUsx
QY6lb4H+VFoKdI+vfPxjtGi+NLfGxZssE5wwwsXHmlUtRoIxnK7LsOj8AQU1sEP3evZSezsrhMhb
jH3Gng6chUNvjxOwrhHThBaLmfHyRSzFxoSCaZGxbgpKVy2nEJcSxdjN8befjY3GT34tQlKeV5aw
YPhbY659jKCMLvhhICQOdjWG7kOfQ9KfL68Ks4F5/0HXWQ/lfx55UfQ3P279thWCw8zBzQ7M3HeY
M6GrC/0PrvZPODHI/clAdI/LSi1ZaRVQDYumQXGcLpe+Gl1J18PUtEM5L9TCERx9sslIF264KqX3
efvYYWtHRE0x77cxRHN73DOy2GwjSwHa7ewlgQnYt/Uz1G3TRYaWbigFwGj9CFJTwfdhHtH7jc0e
BhERE6NgYIMQCxAJYhdwS1t6M4pfVSzpNQyIgZH8VaWXML/OVnSABBf5Y+9GjvQWlCxP0hf4dccy
oq7O2pXp4pd+zuZ3rHdZE8dHVsuvmocS8OB1hE7uKCR8/o8GXYL4/XZAr/pl3zQYbzs3mUH8oJCq
zmQWa5Sypav3dZj8+QWlSpYzKZ86H7SMtrnU+FDFENhEypTtm9OfOVPmhf5df7XoE/oWdjFDUI4F
k27Bi2/q9INNLqCeJPVDXxuxEFgi4zsZrMAwpyvyucEaUJt8HitaSIIj92asqCtg+NM1GiAz+ant
XmaBX4GBsD2zJnx7L2DryxYdYQIvSXj+CvIC2kwjvlyUHcscGWQB7ddqYS8FdE6n1L4lUmfgnscs
DK+cJATTDGQOI2aBHVE46EC1wllzHuZXKEZXygJ7L7q2J81jSuOyrvDXabcWZb8zbbyzrw7pqkCO
DIHKAJl7lKBQQgKQNFqhmfWrX9N3+vh+ifqkDfwUtq70GY4jEK6QBVKM6LSRWKWCIiF/x6FnQk21
Zur6vCyvPhxQVdaL5/T+rvjog8zpKDqz0O/m6gfFcYPEkhcezShR0nR3F+jroZ7CCg75R/RK14Mg
WhuR237dxYkZvgZCrok9yOB2qdkA/R7W4HPcByIVKPX8MzvzDzxRzz9/ihY3802hAa0yh06KLEE7
ifWvUfSfFAEiyxnI9gQCL1uHd0MdI71ifxXAS+BbEzd68OXgXGNfP/8+nhsr3TtM3Ry9lP5piDTW
skVOROvQZ4eFHEbkarcyX7i44eTwjg2TDzPI06oBTTwDIPcfRAhMglfBnyfzxPLdFnbOoCYt+zk/
Rx1lUA221Urrwc+tUgMm/I68hfMzLH2+hyICWpkacFT8lXdt7/E4Un4N/CzfEiYgQRIiaeLmErlZ
bqi+cTQd4z6Nm3pDC4IfpALtwGPYbvCo7ZkTP0XwH/ehlkVCYCpBX1KOrUkqxEqmo3vkCT+ft9yY
xbuYTAdjWxky0k4e8iLMCOLkTLfkcm66NqgNe4TManJk+wkNiXWrjSIKGi5jyHEYvEDTHmZ3ede2
f/lfnFFL1nTS5bLphp1PhJVpuCUZfVtZKgpSVJeLGrSeDf/KV1RxIAXGh8J+Xgj4CHOnJw4NLhMO
i8Qda7i0ocNHKZic0f3QbyhjbCstLy8wqvIVnqGEAaJgcKVry1LdgyfsTK1n65kCWlNUbhxDE5YN
5r5CmNjHA1m+4Tyim88L6liYDPl/QCbvlT0/xi29VthM4POI5k5IiZyEOZxfgmpKBwYmN2cG8VeO
FZltU/PasIXdG7BLzJDtNlQzcd4mILJWi5G4jlGVk0Hh7IqO4nFdhTcDcCMU8jaJwiBqtlCqPMsj
RySUEsTt94XQY70udMV2wnaK0hVQzEbpkrKVEJio2XnWBLyd2K621Ybg4/ZfHSI5TAoQyiw868Gz
Z0vPR0cksJPUjrnDwCk0HU6Ax8MnUsh0LJg8/tcuyVGkeMBFfkrEDafui/t/Bi1lvbsvlRogskO2
yYXVEkIANeUCjeTAl6muobFQItQY315yIYnSR7iAzzxTnJRpxXEfVmT5oVgjK85/bFSA6/BAEURq
/J4R3GiMnXsPqactsQRPEHxPUH4PTbqNryUzYQJLznKyC2njzMTGntOSETjgXhn9mf/aupV4bvkw
1kDFRNT3c2XrzIQkHzrhdbAmGaTfwHsV9//rSdKXnal2m6hAs8s4211IGjEiD+ZHWx72ebqM8fln
2hCCUAPO3T6i176+4pkjmRKFSdNX4/RzQBTVS+dRK8bEIEHChOe6L/KgVePFAhlXKhGoGAYAh5vp
A3zEoy9VOzamQ1XL++1937xNvQR7U0p4D79yYhOuqR3FsebWTs0P//DsRRuuuC9PhJanXm/zGmx0
9NII3gWDPVQikn/W1Gsb37pveRHOTP5dkC5Z72TS9RThwryZ4DwrfCHkBU6Nwy4qHNo/Y1iEHDrF
9OvVDfRYu91DNzL3nTNP9mMfo+Y04YXE0QYuWOmGnrhA2Hx1wdu9VPZW+X7fzJUnfmwNvJqJQywC
qKqDcQwZBWlIRXUlAsG1ZzCi9QHL4rNbedD2PaAuu4EAZcMufLnYWHooJaRPPZMNLg5mqosnU1yF
+uddh5N0di0TEh5JG5ED6MracfRjF+rqJYzT76/Mnv3iR6MaATsFWNXHJE/ui5NFYFvdiAuw9+BP
4UuHPn4tBWLt65XRNIyM+AFT8hUyH/EnQDVmpRahxMBF/AxR2FjnO5bjVD5ZUVEloRvdxFq8zmT/
0kYWNyh1q8nJQbiMrTxSCFP2+U36c8gjdt5PXTpiRPUf+UIjpSxJSVa8s8J2C/UvFHC0Zft0KyDF
qsYy2Snn/lY67G3BIPhG7/2plOpkPkwE/hLYpZ2n8xR2znMEKxyUomRyWJZRHqVuIkD0a2Iob222
rVaZNf35ZbhncLc/7A6dbmebSRAl2kOCCo7BxNFYzuG1HIKbPhruAg6V1Ow0/S9C0rv75Kqanz8L
ytpemkjkxW+cOKWXH3erA3du9nZER+yekFrLrUTfloCu+ENjbk/qDpgYCmGFF1f6m/r7Tp/6YXiN
09ijzk8G5sGOxT3z2ouehuk+hvpWvAJU/+aOo4vTeF9gN4F8f7IJHNow6lws07aT06r9CDSbgzL3
ZSgFj9tFXfbPso14cmk/ebdmaHO5FZE+sLkcjVe/LqQ10P7jYbonBY92phbclnUFYacqFYLmxMd8
XJ8QXeHb/aBJorQtIL73i1rumuWu3wGBgg8l8vNQ6mOi6Ydu6y7Lw9L0XxnOsR5s59GAgpfglJpK
FVpmy848xLsJFdPdDfwwcvkeylTc7geehRwscr35JLKQCko2LXjJW6tUSNfGh4B1CZIntSdTMibY
+OBoZD/HxtuaeQn1LowxLALfLbqfGf13IwEqRT17HJw8BsauNumeucNG8ddNUztvuCv292Udxoxj
5YQX3Up2VdpQeAuP/WKfTcd78zBcfBAt3CHPJ5wN5CntaZdLaAzR8o8ldQyMtePowa6EUAe9jpay
TYzycxggp8P+M9zwh2Xq5kHVM6pen3yCJPVQBA55tvTgqiYg4ztrKC0pqGf0Zkbh1WaDXnSY/O69
4JL6DBLgXIW3EyZrsPyeQEDbilKr3cUahCQaUMOsfLPShpoDIl4xmntzNkb6NChJ1/R3TGSS31sQ
j2kYoETXyds4ZbIHvoc/Ou0eCuK18T44dXNJmc9eDykQJrjjXn4z41J4Qhrb0fkAJUAKSfRRMn4N
GbMqcvPgqkNbxBncaYbfYsuxuYzbnO1nCNYagklha6apvwSgeIJLKirnNHRZYLwmJkGaFdfQ740D
jZsiQT6taFL3HNeA0E1/xaa47dlZhag9EmRf299b/gON8riS8m0Ke3Ihe7L+xOM/jom7b7ug8/RU
9uYgFrCB5iDa5+53W4FGYI2QpxR9OIVrLgedXJBjEhIGBjYqfLViG8eGs1j9Lu1PUFz0BaDxrbRc
EGupqHfVm0UNvX+q5TbvTDPwtOwcGOW6TFbmk2J1L1plk5hCEnPiXTfM68DviC3LOQrTjTn28XoL
iFboDCxizICvn1pD8kTX9zZZbNHHh8jr9nhUKNUXpZ12cFC6myuTf/xhHGvd5zDFHpw9NKfc6xZD
CJS8kDkmmtLWIGbRuZ87gZnXqfX68ZJhsetWz6z5keg8K+2oQm90UQAHpep32x/QIjHWXh9MXKzZ
I4iZazgRIrpcsBAjRnYp3d138qKv67kjRVefKDQvx0v8YQZO+2gIxiZ4EG60+i+BR0kiweIXJSOw
L6JSgPoWIhAOicHzgfSdLXnBD2vVTJLQjB03t++hXNhd6SdxfKXMFQvqOvIANfpoh4YvRU9J5ZnQ
s6QlwgokWHRT+1+jNANQFJECIRQtirMqHunoyJe1XrHGpt8fvmSD9AEHVdRq7FJ8fUYEMZFg5C+1
1Vr5CgtMaGExrZGnwhJfkoEdRF/u7BhuVcQUYFMFQPfDAGfZ7ZCZfmTFRzTKFmoMLCII8Q4uJr+n
08bsM7sIqKfdFV1wDsccUMmI2BWXrvnyoLO5vAea3XdaycwL/gigamZCV7aHfl+YJ6LmRDhAm6Be
BSD6vQj//rGoSYKrxvTBpTdScEpCioXjEKTpOU1AeEMp6n59r/ccWFQvT3TNEDf8pKMNPF+/P+wQ
cv0qG6x5ze8BxT0om4OiQb31S2OvL8EkJWbSEgKzsMmPy4mUviLM+UI7DrlcH23Hie29WzAtFPBd
bC+igc+Kna2nwqt7MxstTLB65XpwSB3MSJNRxfGj2M6mKW6U4lflghvcUnHghDs0DoYCWQAIJ0cy
d4jxWH9Tkswu9Xvp2O0IDgMrNfasRQ3juWXNGyXLeMb6oM+/ftm/zk6SuMz8olA/1e06KjlGUwu6
HuPvE/O9GfDDSJXZms9JOO/KKWNGL1s6nkcEIeh1CV5DbMffslcnn5GTOMygLbPVzE9GZ+evQhYA
WhXyaHXj3u1HqeAGu/1pbRQUHKTCC51gJ1Ifov7Pqjct2f5ERlV3ZT6BwsUVHJ2D3sPm+IwtA6z8
D7yfUxjxIYukSWtoFsgVCzRoq+rTGQytOwksKbEznWpV/K9ck8CECCsuoVMUuARZ/SSkWJweEgKB
xMhU9gBqGGy/eJ36QaNRmumdO2K4xOT7SZcljUy6N6UVlexlnAmcEINpOrUKpLQZTc7lgJzcx59n
2b5fQXcm/DHraavzjqve4WiANGQ7/wLXyuof1CCmgWDpqqFbmi73M628mYEh4lQsjj/CNUAd1SdI
HPjp8hikkuwAnr0e50+PYvoTzALQ7dV1pb0NjANW2MFFX300+jQKTOoRb0F8BAteSVuFp9Zfz5e8
mN4GHIn4l0fxWsnUWJnw48STUlzhmn40+Rr4vhzh3ToLfYkAJvtRwoZ+i7Oa2gttpN2LSwGfZYZn
8sgDjMN2GgI2+BhNuU6PxbHXK8tbHyjyMtml5N8oL1EFNM7jBT/7Jeh/1XR6YIDfNGjj9hgmENOh
W8AUaw8F7CHYXICXxSmWQhSvUR4UpoXWSRAgA0EnaHsECoDojZI7AfjVd/9Fqr/G0Fn6UNfJcJyA
npQvYJuaielbWz4TAjCi+wHazI0CB4echX1sN5pgQYJ/QRjathFkOFDoHAqkZF8QTiMEIeWcSLEt
bcNmxz5i5oh/I6uqlmdDo5X8EVIpiwcAg59+T2cIvKVwpfipF+PkGFewvxnUA5SwM3akTkr1X0AR
cwVz/JOpySFLyjzg0tvtqZBF4RAuNyLjxdOyBqfoDM+zxUiMe0rIBO7wKGBZG/kQLSWBRePOB1IV
7OtPgbaxCBsIBzjZ7s+x2H2T7PrW/1fdhH7+9CW7wBQvHEbW8CSHOK6uR+fra0j+2VbyZJpa5U4A
V2HUhQj7LrK6CgSTic/oNF/F9JZSNAmJ69f+bcUMm5cF4OIFzU1kJHLi40rVwreCUSRctm77fYeS
YafIexCdC7+0KP0RD/vfK2YQf1oiy74DenVRzE8PZyCc5bi6UIe/49dIpd5BnJCOSCRcaaqXAN4b
4JNqbQLlbLxn2SXYvKmV77KmHEGiLd/gsq4vAAv+ET66pURwRREUCgQEuEgovULcuvdc3OPhrqtA
Tm2ftwB2S/JQKxwC90Yck85pewTbC3MjE92eJg9A/jwzC9i3LISp8geQu8Uo3gvJXQlWGdH979Fo
NCWmLJp13O0lu6QDPFufIR6hYGJlyNLTwnbaLJNz0WClYfynklD8L7cKCP2GW4DwXYUW/O4u84sM
D79qqjpiHKQl5ZVI2NLsWxIIozIqXAby/nuw1u/t0jEAr+y/MaRMpNIN5Rirkb9EhI5XefZ+gT3J
FpfvswyEGOkX7scg4eELpBZp77f/GEHBv7wOZV/K3+ncNjEagoa1WkkeY0YGjczfwReHydkai8oB
XJ/pN1C1CMHLaQNdYBiofYGeufAxJ7GOrK8E/QN3HKXfO1js6GkyVxLz4U55vf97/i4vnrcO0LXK
/YdQwgFax0ffq5FUnGKk199YcXuACTogGMXJIBNGkgd1rL4hPPW8sjXjKYQ2L3Y5bvYCGN5PiEMF
98OTu7wJrVgLyw4tkUbbfy2DjgIliSAmNUpGgGGNZAvFdG9eOmt2xWKAn8hE28wKkbXCt6HHZXFH
ozmJe2S535O5go+497TGQXUsuBvY+xjB49+C0SZ1TepuLrYGXEuxpgU4rZhs9vCc2Ghq/yDmlrNe
eWpw14GZNiVSy3OXaywdOvy0oNsyQjq4EF/J+AdxybG/TGErsVQLMorzVAFZk+2tfwBFntgWvHE+
T15SYVSfOkhTajy/Ur9BZrsm7xRetybY49zzDfOPq7wJKi9wHM9x95rxCkWBamm7GwPjUacs+4jZ
NzBBDoApC/FkKliYuDx8sohS7MoOXC/hT4Tb8N0VYjJFlZL3ZexyF8r/oJPK9gT5CM9k0lpDj5Ea
Z8nFTH+aZbuVaGx5XyFuMQa9wBQvQs5SJaJgESMl4HPlCl9mUi16WHYiH2ET2T4qwo1YYjTFL/K9
/xu6UfmeOdKr4+T3ectP07wis6UIHYz4WzmMUv5tlHXayrbfe8vE8tJivMuQHYQTLdM9/NCkjcTQ
TGxKurDTZNhZ8V29TR7yC47frAHB1OzGXxd9NwNUydOS/ig4q9wKt06qwMCW0DVtqPmoU10gcSEO
rqxDPEyF4tVTJc5JBbrvXPpbeL8pOwrO/40WAlmBJSA6388MyS14g2bBgev71+Zd0gVM0rumhxar
JEox4BjeonAECzypHiwLsEjL8ZwFdfHk5SpinqLYDdtKvMk5rPad/uVzUF9YFbE+79yONM1UQ1ro
Y5h47Xvwm7em/vY46uEoAobaMrjje5Y3cRuPCVKVV+U2lg9yIHApjcFsJjBEmXcB6tD/atR0Px/+
WAkODTI59i/7VJS3HzC1LF1AXAxJu4nAN8VAk35hQu5CVZP1AFKJDoxOBCaghoeN7ZykVMPMyjrQ
2hS5rMmk9OknzEvxNUCdPEFS7PEnO5jaIWtyIPSwrQ8DwdkNHu+C/ei90KhgMelHHo3nTbebSLht
T6Sye6NFnEUzaKVAGoGFL2cOpTgC6WquxUK2GIRog7ClcRRkz6kSM6b19ooclbjav0xwvgTWgtOx
Jlgw6SmcTHbpstezAtE8fVTJGKWyjOhTmoalr9iC8YWAcrRnsoFBJKdKEiGWG2P43WmYaxkDF2sO
cbcl4F7IGjfr4N9i1UYehRbxawC79sQ92TGNmCvWSZjdTyW2UJAa9BnebSkIqJGZjaa4Hj3KuLKJ
A8Vj7zWWlWBBk+zdrGnG+FTV2D8rlmYbLI8CREYac5HV5Zl8WeEThTrwwUSv3Q3XAxbk6lzD8iJS
TDOmZNpRMX2qnAepyq3CbIRXdanqkIokNRlE+yqONAGY2RWyxZgbJFJ3ViOiwIXZ2BU5Nvppu3Xu
TpxdNpViFcD4Ku+VTKmqV2ZX2vZamG4IPCcZk4vYE+pUptWOoeoHiXoetpc+YlQzN+Vyk2PtdnwD
jkK7jd1hzltPJ6IopCuuIbyDufBDOH4SVQiSeMiG0UbX0b10AwfN2EOiYkKVFmW9K4gVWC/PXcwq
1xe5bLETbJ7A+5iRoFtIqS9fpImln50LvGZastfYWEi940WNw5gf/won5KMkeTSzftupbEtAEy9R
8vUEq4MrRmgSaSXLGHW5YmarbpF6npmP1gGvGM3GlWTxg6h0nuNs5vW6UvItDLaw0NS0kXD9glMS
hDworMaM9x9gt38LbS9ushwzR2AKXxikwyLbKlfH+KcUcND65tRg/BcqlNCmtQor85TnG+HIAWTo
mlMuKeRf7FJ97fgmyywla9l9FjDNb21C85YTetVLUFjVToQsBLHcvFcN4kIIn2XdRJM2JDBRO6Nm
A7ov+EcjGCIlSBZGXFrPjkdPSi0XQcMnOgRZwTS4V0BPTGRXQVVTwkppu86dWoOrmhaSegJTbyE0
lGDnly+f0mWyXuoVNXS12B/ExRqZK2MM37R8VEqswo0saa6bg8xqyWKxGY9ft8HmnOQ+ajUepjEV
Mq2JJWzkkz8PZYi1tRMywzxPYhxEW9djGaGa1T8SbVVls9FTERs4kQxK8sCHWg3yD3qgoT/tNX0G
FATSWU+nguKVDlqDwg/A9QE6dYnA4RiTvkslzJFHmSDDW2ZPJiespjP2i6ght8N3Ixi9eWA2Ojlj
DU/Lu33hushz+MBMsOpt7c5mWG8NC0AEntJE+sZGZLdLCl5H9mijvlk0f0fQvpxxh9iA+aFB4wSU
UPTbY39vuBG1OaU51TpSw7gmJzZI5yE4BlbB8jxkB5iOaDaDcI761c3gR+xnDNMvYd0X+lK60PJl
dDNmcx6LTviX3SfJm/edqzM0nUILPLDY3QbSfNLcFrCaIx6Vd9vFqK7DrEzbGKB9xm2ySzB7/MV3
GRFHD6tBs0wCjr2t0rTZV1fl3TNENvoP6D8RcLOPiLL9I1hZKwLRs4sNarhcBIOYreyMZEzqQjEZ
/3pFPmNiqhhARRrGjQCvsVBDNPlydFKYF2FffAafG9etj2CfkQ5aLAuHJ1tMC7N1A1IXBw4l5Xee
ePj0Zr/eGY6BFj/Yg/FTiQRq1DWgdG7jHKCH0YA9Z0rvq4srtJPSDfLe5IgX6MyUDlx9/A/rKW9G
mWJGYlImlbp4wxctHYyCpfbo4R0L6qI8FfMyT41yKyNQoExvPTnnI7seh1NjbTTytMM4FF/Yk9oE
x+Qi0d6Iu849JpmbtFPTzdMooDsHZMKtFTFUfiItkZ7Etw5Hcumfkee23w9evYKH6nR27dcs912+
DVHL4XDmTHZbAiv678DhKf4E+Yj/OjIP89oI3RqEj5yJb3BlF3FCReXTmj4zVQaFA0y9PLQwKP7Z
DsV8nJptLmV3aAZu9Eu1BrBKqmCz0W9vMfPjDI1qTSRYl1d0YKbytb7Wf7zRTcWk7H5InWTHKKR9
QyCXVdFjzMdMe61y23U3a56rQPMXFqwUfpduURfWjGF3Wju3orOJsXB0Lvmy6ZyJaS0uBPVHEzuG
aLugL8CLpJYlG2+/V3NGGIM5u64rmkocBfK6MLcnNDNV57Ewq3lWmH10KWYDj+WWCBF5FnXchXCg
QvXo5k9/xn3XQg+sw9/kvFWT8qozle2zCvvANO8aD/IZ9F282CMFLeVVtyQrTBiZNmGAJZvI4ttC
qkfW7B7y0KhF/4v6QEsgM94sKLQRVpwaeXT85gSNNL7GUQdJca4L2tlpKr4DGgNCHUgXGY6Q+8RN
xNsmBnFsgKqWX1utWHSHQzx3zLZ/16Dx+LdglhCh3D9c9egiSic4OUBT7SC/mDr7YfZw+hOj2Crd
HN2UFcQTAmpf1jJqyJg45+ZcM5DXzd2p+Z9vDfpVeieYPdjd96ZaudW82+upBthgXERoZ9RNY0hk
tvVHjws4i10wLZn4sqfOMAzPXDOwAJ0j6Qmcg6hR0y+FB3keLF0cwKRytAH6UNkTUVl+X0WCxwAt
WxrqdQeXTO6sIamnKOZC0UfqS9Jo5EaevKPi3qZVQGZctpdaRSYZ5347KEbVIbPZI6XFkumRH0QG
g64wwYD965oqD4LC5fo5VEkeqXnjI6BG/tK+d2FlrVbXsTPUgW3BZ/c5fCkvROMuUspHjBWS8zBN
SBXrF0jwRYgsP0eUFH7+281QRbjHmH2Ffpw5pQXoOAQe0cd8hynoR3RKmP9OOeaU/734wK94puj7
h+w2F9q+gDfBXejhdsPwYyMzgsQMc+TXYW4nBcUvB9jOa4wrQM2XD3NN3TjJdQqRIjMwqsHGWpjH
nTGfeyiIzrJGjW21WA0xM50FMVjwSomESMnLQvEOfskNzX7oQ9J++7WM+JUyDS8P20ouS0PjI7lq
903DIHlGFm1Jwr1WOdv1jRmMhlsHacyY3+2EFwh7lE0ckkYYtLoXqanYjvVDOPqMiQbIp0IsooIf
4U06hyE52HTGLTW8VvZL2jvXNpPWX3/1dH/4rFE+MXLb3CFPULol204BuJibv+rl8rnNDmhbFIha
He5gt3R+jqhxjtV9fEXGKHOw9iEE942y/e/2wOwF0gApgWIjH4AoXGAzEUXCJK15NzyxAAR6CzW4
tEvV0p/VkDrfyFtrGS+e6fY6pP1lH6VpLveWMlN4eaOixKhlv7cQCHWOpNkEfl0muruA6jhOo3Rr
nblfMod9bhQSBlFTGgBwiaNSgxVCNly6sGIQEE8zFg4/SIPdtQfzy9SMhnzXTT8slTHBsoU/1Qof
MY5oVuljWi3fLUIHR8ghNX7B3dFknFDxOmDXGQMe68G5X6ZlcNCm/+LJZFlTAwKyqzZ0nkccRw/g
LTLN8eBe1aafdQIpt69V3plMvZdNamzFH3XcEEvmeXvX+fFOd03Y3J1nVhzaEI5oPZ3DCT5Du4OA
zlEF/DNni7K0ZgSYosbGoww6pNZKL7astcovNO37jNt4S/3LGGaUhtQKiJj+iZOv13NGStJdMRLH
/PjWTPtlf3bm5MLWLDO0lSs1OiEhTNuYY4wd4kQSKRmQb+a007LCemb7hw88W76OOA/WScklU5Xc
OH0LsJJV+3U1Kb4DagQa2RSeTSMukaxo5O+vxQHqM204DTxjK3CeIwD2W7XpCzO7N9iRXL01ey5q
5scgk3TN7TcC0abekzBLbcGvEK9L5BkZ6P+GOYf6CbiDNNLGo7rnz3qVkdsifb4ag3sSjk+pdJCf
rx7sYSU4h2d1dB5eZo6xNnts4nmgC+PJl1yrVVy5YoDc1b8AFUE+BOP/+DhdIoMa/mGZiBUMyTLf
n4fH2CceBxDpDV23VScoRDp+edOVgsNCNIY2Bip99oMa7DTMiIoSGXT4bHORW7mCYkaZOR8ztSR/
KJkdQL511NeRJwCUn/y8+gobV2U3NaQxwDTI3mVfltSyPmyJb5kdKPOBBgjCagE9dqVOkey+1IRW
M4a/rTtQ289py8jFu/3UgHqCV434NJb1jFHr5zdNEsW0AxdjE0X0H1TBP1Bb9uboHSoIrGtgSyuq
gFmg4sOxbh9y2UNNAMfUa92Ae7Q/uI5U1BF67GbUjn2kTg0z1T/uZvIE2s3jGvtEyLX9wmY0d+4z
K8pzBs3CnxuSCHjO2AGRKWbbdxs1wPS+ZUHtx22rW14NLImh94sXIUhUAXiPZeaud6JDn4NEpXD/
bDH+YwkG0PbnAtxAtR7S+zQ8l8rhCTQNLOo9h/lVQA34I6EHEdLS4xgbs/1+y50rVszs1whdMYsK
BBfdguDpEhsSjYePeIQqgwZ4lXCPl9UzLu7KplNLjSwE4xVnlnwTWygIcNGLh/wAo3jtuhWJh79a
orOEeLOZZock6keyetF+h+acQ2GqWg0k9vqZa4Iau+A09PV7v1MgV2Q0o+SXIR5rItccY7ekhkqL
GTdJ0bZccH7sM6GqkoYMf4VJx6JQ9dY8lrdhZPNPXYzvgQxokxkQHNbqKHXbA4KoESSV6GmqOvFa
WErrzCbEngupWKdORTdy/BMEa2pOhNPQ+jHRxWoSG5WjTJnkvB7536CHUeOWH7c/GiWPc/ZlwLTH
ZTKeDeqtZuNzGIDL7l5JXez4fqCX+ipFn12uK2Z7eVuL/ssCqZCGQb7wYbX1Q898KlHE/WoSQBb0
3CPjlfJiT2OFe0hyaS0Ix8dIDXHC9C63l1joSk1c+VBfUbZzyjenMa+zqdqxSLtFw1QKyKbRmXFf
p4RIycZcNbZZOqhafpn6I2dwMr/d+V2YnjSdEMdOAJywOG+VOk4tMBjMhFHk2c8Vg3KfehLd0uRO
LUHCK6YPEaEf0xoaItG4sa10JAsGGaLb0nH+jSujEyYn2zQYW6yeOr60MAHff9Za8jdvVCh6DXQU
2b0mKJxXFQ9cJ+VRFOuaEwRmaZ6Vp7SY29B4AQQO3S+fqiy/oto50UIhZOitD2p71kYRM4fgHf4S
crn2iYGgbZCXLE112gUrd+f1TjI0VVJBzmZKbpb32SKW/HyEbqjtciGxbBN1A51AVX9/KAQN5FUk
hqSS+HLGTiprXfySiv5bAznsO1rBFao1SwoBFBd4oMvnPLL1vaHqp9lkV+e8yJ77jj0BLmEqLQQG
yKEBCgg6XipnPxRFDlgDCm7h/4uo0DsV0so3OA/E+CCUOgb6ze6o53kg32E2RA7PE+9rRA3E2ant
t9qkuCG4TW/Yk7s5C5r4HMtRuP4wusQYYrKCqWRudGDOXRCaj0UnGtoAM9zymitnj5JRSjQI0NBW
vtbETAMtGBXz1ENez9PnQMPXcnBWMKJoZpGi/RTeh1Gww7PebAERHQTtMWa1XulhYKzCttNTActt
/IrfFMn05yJUTIF3Yc0BCN7DHqal3CSHd/l5TYJXzGunkHPItuNWhcnPZi+8/l0mOnfzWuHtWg00
KErXv55aFEvZR80T+wl1R35qo/LvKWmIATq7cbYgB6boKmHIrLAHswOB/p2wCropBtpjR4cMr5T5
gppNz0ULloGmyPXv8MVIQ0BRAJ0e5KUdHNlJfD7yIFpzm5VzXREEVKt4wM6EO3D8PNauqwaQrRa1
7pepHdDmI/H4rqumhxa5mercEhbVnMR9AbGU+XizaF7CpCuKOMJxcWHmkW+DGvevkyOF0CrU0SeD
sRD38GfIKN6/scoX/2yr2xvCSKW4RVYWQAF+5/tfG9dEfM3jvSjSw8zxeNpi0U2pd+Zy1Z0f9Hyk
XgMBWeU+wJpx06FgGMrPwLq63ErLpsfs1PTO5y6RbAtCEuc8VNVLcE3GAkCMnIDk/HawSA8vW2eM
5MCFKpfl8kXamGfiKGeAhLpb0QwfHrH+8o4lk2unaWqiQ6NNZy+IH0hnkj6BJXjfjiCtFlZZlEqN
YfoBAhjYFnLQqZqsLYmtrlzOeLi8Uq9/M/rL0TJVEBxrDzGXRGs6gdPUA/O4WDm1a9kvlWRtQx5E
sSiai9tLcbh1yNfMzAlD0+w1z3+MO4Yi6svldnUt9nPnT2FlQa+3yDfKObb1i5ubiCm9RI+ku0wv
UCPjYJobqnMsVOJ1To90C5u3P2/v5wcLdccwn5VkbX3jdrx+4xjDAa+1MA8WZg4Q0C61lmvY0DzK
JuzU7SOdI6N5mdRm+pVu7NDh4Q55xTlZd4SdibW3ghiqTcg6ejSfdGjCooDEcjvcHJLDGh4CzRCF
VudW08zBxAHvUguGnDJy26qXCqXY1duhg8LjKDqPKk2zuN5EUHCAc4yjqLxzAjA/G/tmfdk30I9U
WAtDmGYChhFGdcaqprBgWsYqkgOQ6i6y5nE84Gspmi29tUpouy0sKAuty/z3yZuNBw5K5EUbqzta
szxUfrYr57Wwxlj3tTSLN3QFvOG9Ha4AgN+gW52UYA8dvTM0U9VjHEo08G7+I29jMACFdzS4Gnfm
mKWQ8QOAGVMLJ06Q/AL88mMf8V+dYDCQshCXYJG1UFjQ+UMrfUic9jc54psy3C5kNj8Myh4BpT0m
H4MNlmb45sWwtP5H/Af4H798roCA4Ss7p016+hSwGPKMzrnsRsLTIKg39kgVEz9Ft1L2TzHYlekN
XAEH1WSyAebC++pPPsFQo03LrOrIIcLZqskH15dSDqN8hM8Zx1BmAH+jCQev7M4TIzM/hKPgl/+l
7QCVe8pnWOtDLRWc3f485IYy2U1c60Al5bGq7AgNm/1hQdsqxrlVQfw46YEJgOUtFqA9Dn7yCUXj
S9PcWkAEPXhldiYSgYQc8HMBQzadDHrFRSDGkDsAozcB9KMdU/j4XkiQS4kfSJQg2Q3Wesltdqm8
gn36WPIQt8LVOLDF3P8BUHUs96VkJ+9wf7jHFAhxGbOI0NWia2CcfCuCOW2F/KEENrJDJDKnC5W9
8qWY/MUqsvQIwNsqZXwjLQA/0bOAFRYI/X6wgdu628XutPFeWn6OOWvjmt4lBddS9Uhjc/63Yxad
7WGPYyb4//opPnhUXZq67ZZ0rXJ/EM3WXwfCYWqbvv//EQQxWuRkB+hoEy3LaGmKcRZqjlH1FQDj
mRWeYxJKBZVJtxPmbTKdul73LxhGVksVb+n/fTnTJivs4U0Q9zrZ0YMmgrh3x1Y91QwL5ZhBDy5X
KQWM5AS2r3xi+ORoelAwymgzeCmFUL5coTTGVpgHvjQRtT4jBjsufmNeVfFagATaaw/hsa2Z2UVg
vzf/1PQ8b/KTBEhsBBhKGhNSEbJbGaxSG7KQNmvW7yCqH3vyfhlmYSU8vyq2zdKlJII1wjHkyM+9
QVE8PPs22H5qt45fKwkHHdJl6mYeMhmZXOtsXI4h6H3EYhvKmJnr4cu/SYteOfPC1OrLAIbhrC+s
D8+CM0O9IvNY3+fO4CpIXyuM4QETquWwIwthUJ3Jn7OLmK4o7NzoNx9mnbDFzA/26RLC41l0O/D1
tOvoP+FkxN2uGPdq7KVrZNri1z4lx9XzIZiLMI/azJMOPP3ESmoEqXU7cYG3ibAk9T/G+zVPeUVA
Vv4VeH8VvwYOaddffPq6IgKXd2N8vd4yCKkgYOMImMTCGTl8RuRvq//qIugmUmJOU8nEzf+HDSOD
6I6gTYvuTyk+9KJeLdQ6AsL8qFuGgdSFqUf3XV48Dv7ndk1CZbUoaZTmLvSJWY3WsZj4sWJAIEPM
6TU1hrVuw0rYsXT2aQHnLqBYWv5T47yNn6WB22WTx2HeUvAMs4qhGKXAOHfRRDeixDrHEfg/Hvfb
c+2MeF82o8q67TSPTFRWWFLQssrBzC/5vsBC6pG3CTIzUH5ki1kNo8dIe5r7eQhKOh7JCX4eIu2k
tllc0/ba7DqX4ECnt00ZM5ddt7pjyCKALNT2V0FheP+ANYvA6qJ1mEA/OPmAfYHkjZS5PlW8y318
AYzCjBYB+WJCxa8/SRU5AArRHRtNh31f4NpCHgf3KYcbgwnrwP7qjkcfjqSpXQoLxuM4TX15+KFf
IzLQHNbtNv5bn9VDBR6Y/1X9761TdwRibYmOLnOQSzxrV5A3okHmTZorDc2TCRfG5tOD3e0pcFqt
i1/MjoBNghetNBlvMU6cGit9v5942gQicM6MwXTO/qq8u/bVyvyomst6vxkFqhF67TGWWwEGEZQt
TCpc8U6mIF6yk1inXTqfgmGYdu1gyLlQtWRMWtvzVlHI4pNTYwi2rlX7HE7Ll5uPI9cwnWRYEYzT
gR90VWlmxjPWqtkDbnEsokVd77G0Vk/zmRJGufo259byYN0bwHqCjhZrsqvLICH1gwIsFScqPwtc
7E1DD05+l9NoWQ2YkDEyH7xwh+tqLvdtGRw0jKufR7DJreJE2TTN8JjQwpANPvsXLnTJJU3vYA26
8WOVyvbid5O15nPBz/2LY+SCiLdlUTJqob1j6jSUagBe9OhRLDeRMIce/gbgZ2sq9btu75QdpNKp
X9z75x8kSkZeRyJT41HN0j+pfLPfUH7oMxgS13L2Smhc5Vqc+W/aqZWNgICa73qF8ZrokH8bMA4l
uZVgTeWi+5y/HgRzmbD3SyMEaEKHSXu/YZMLRFWB2KKX+bldFN3FLL6A44PYh/GK7Rp0KmE+bGJz
J5p6J5RITCwdO1y9UZ5Pv3jFukvBmuKpyFhLPi4zjrACBHqxHe8CE9HkOCXiraYes1rq/KTFoit8
R7iyB5DMc/+Mti3Etdpoaciyvd2zCxeEvduXUSGNsqAgd54MCjByxVjDDwoy39AEG77JHA2044Qj
gnmWJb4CmMrk3QywsLm/wUjtCjxcV/8Vk0DQUHurdMeEnIbEaSDwlI8KygRygtbdQ9nN3sCZYhvN
8XDmL3j5qbxz5rwPDrKcwrm4lNh4/GmuXpS7DsbmUSZcxaVdgAAMItRwjKL+DPdTaqBe4+6GOwe8
ZYzEMoAkPd96QI5AadgcUPi1mxdJ3QLIbfWyAxkGUhimHAT0ezFylmMZDAwbxRnxrP+Mh9jpUbBj
q0di6inEXOosLmIkWIzzBPrt2Y/OI0rtmzWaLj84YFPmTmXhJdY3pG4E4L6mCUQV0hhGzSV1TD/u
5+pUTXMuJHy3qpMHLbJ9SNCn99yhCO9mQ0PxL24JIptMSxdUNTHkSVDMeBa7ScRFb9Su4G9GfmnO
34+gzefNI4HUx8k20EjntzR4DvExsgLLgiNv61pjXMiw1e7FWmK35eKPfm1rw1giXlJTq9/1opFY
5NhK3geZogfqK5jMwYW7iSSZWCmuSCX8bpFbiwDvtvaCGsNCSdQ140rJp5K4vMkNaQCrTp1vqzfP
aX+41YSx9A2Rru7NwKGJ6EztuQy9OH1u9IBJtzGb3CLGmDuII16hhlryjGqrqLKE24aHYyCxfUKf
/xhdelE80SJ8eTFUcfYnwdFcZDcuCMshjemf53nbTvyuVCdtW+oumsP+ize6ILRONgFTwKa8qpFv
Ga33wLrrWt0XT9osv1RyvjqwyQhAyleTtbsT1LHR73mEL1Tp5dOUop109wlydBsrggdCMcdka69l
Shw1e8dN7CkST2Ct3Hy+s+w7F09T0JeMAxOGilylAK8F2LS8LGguMhjQEv8BuP/2uuLl/0fOFA+o
3aicr3UB78R4AIYfe8q+2ZqLJ1WQeqneIqzjWM3a5DM1dIYueZhnrp9lxm0ZSxKn2I5F3UnxJxWL
1jK4PFFVbN6DPgyrTxEB/JUDCbn3Bm3uwDpiaWl8Tzdu9KMAg2UWn3AyyRLjYY0oK4os+BRQcU9K
+pn/ytbWPvN2y7HEBrwUeSnfiEhSKBwWAArCV7am5Y+dQt2x4wgSol4vukb1FlqtE5OpB/bKIlfJ
p6BQmS61FY0IfxOR9hvqQ22W3E/iO3K48t1OlGB0B4rBi91qgbXZ1A+gp1pWXnfKbDY5SDURk70a
I2nnFo9tw2yK10j5FesLnj2DYqIvksZw0Ym2egqlAR03q/aE4P7aW7F4ZC0911QTg6GrOnht9oZr
zOQsu0hr8qnH/HIG9PvmXLzxIJXNhhU+EWIPxB9/JfAa4mZfAye7Hdz7DpZU2Zg8PKKxfYpsJl1u
lNTn3LSpc9iku4i3LpDgYB8MsA+N+wPIaIl6QCxek9chcH2khN1OA7voC5WRDF79OHJb1VydHlh7
PBWOpqtFi+/3HxMRVs3FxJpC8K0fiZDbYXEw0wTP3aAEbu0rbdWlRRTAEn1ll+6LMGxi5D5yuYPU
vRhMumz/Cf4cWsvqtaaqCOtQBnBuSClPF/nfJPN4JI1Ao6fn2ToJ6ASBY7ukE3KMUKWCt52ygTJU
Qb8zyDTjriHbcCHL7ViNgN6YNBdb1n5QaT8M9Sy55V5J3kKGy0wlbz0E0HP5pebZZAw6PuCws3P7
KbQckUzcu2Jraq3AAh7+yGIu1oOE5Pcy9bXu3eAZCRsmzT5UuIuijPSrfdOEe5fo6ss+eUB98Mvh
UOBXcZ+6DfaGE+ekQO0W5qo8cXIlCGwDyn7ZrjzwO3cp2jcxcV9squYVrgOoI33c7EmYUkoO1L6N
9spXj3KpTstKUtV1Ylo1btyaOaC+obp3dilerEP5JnkJMHsoDIlTu5o8n8wx+sknUh5NasMZVjTL
VqAWPd3gb8fgq+lLRVO9KpJ6c263Lh8Wo4+quhYUElFU1sFYtfWMVDDk+sRpcuPjg7M/0OBcnzeK
fmDkzvjh2pBR2ut/9k1bb0A5UwUZcMWOj6S9qVR6tFB2a1snTbzYzP4dmTDVIkLKVu/9oOe+kDHB
1FsUJv27HPlvI8GPxm9NASHRJxBQDxO4qws5EoZsGJt/DGxNxKRA24Dx0BOuWSdj+YaKm4nOp72F
RyuzTqMSKQT1k0A5dKEQt0u83a9H9N7uPAXG0He5cy3DMl0exG5ynwFjegADJmdpr52U2P2sxW2i
wsBCZwqqqfdY8eNjtVbBKgraUcSnXdV7dUL71KX35f2zgJ16YcVOcrTrrlkjuBx0wsmi1S1T4DHV
u8ITKitnI38dKJSWq/MdjOTXt9k2sCMnzRP3f+gxhOyBeRFszMtV7JrcoWrHF1TYbL2q4gpuyJaG
664Nbtayp+qE8cOdhQ5Bfmx2Y7fY0hIXsFSI+9X6aIFMuFA5WVKuJn+3WGgsmgTAzeHNLnvyVu0K
ggfvcP6Kf69K738TdpiT1ISv+ix9rDanKX6HZsMhan+JrHRYSfOEmKO71zI0cS/esW+LbtI4TNK9
/txAE4yTa/NGhC1GQAJ46eHQDTJe6QIKnjqceS2Jhabtviwrao/fFJKRIf8n5+kyQTePvRLY7fyQ
XR9KOSyXx8nGlGItK9N/X23HeSjIFdqRCiNdM1X3kt3WP3WszPienjIsHAjfGNIu/hTcfG8fl4Sk
TeEoxkhXthLYlbv1bFyrbG8Zsi4WqRmqb9xw9mNdUhtOPcfUuBauC+vHxmgGo5YqwaoJ28YX4W95
5ZIQSPWFKAYtA8MyMl1I3aij+SL+OFDPLSHD9IMRqBO03lKgrjgTVFiA2d2N526NN0rYXRXY+ILB
dKLO4LKLtBubwX+JbbcljxlCwxQxY31dda7C8haBqkCcumAvRHBA+xjYQJXf0+9zD6A+KKjuuEJI
7AcfVEUermQWSw4JPVAhyabzgxv518iMz+Yssswj7t9MbxJ+lmfQsDKC50GfZBUrCbP0hFpMFPg1
7JzNHGjgh1rpbDyrb62Y6D20ym1yBSDCQ1MEESI4bJmOMs9NoMU0C8TRqgNfB7Te/dZvN2cE0RyC
UEbGO70iHFHeRMjBcA3JO0ZrD8KFdLsNnIAtaBG434jpb1u5smmUrey7VIWunu4NfRrCrFOOPwCr
8s3Jr0mFb+ow3xZ5aAd9l9/bQsIvPodaIWOMm+8jUVuGW9s3Jh2lYRfiVvNmOXaJ2/bUDw/+4lwW
TXpxuxjieULLsv5g/QiRwjrErd6kThKtiEPRWx99pVXFzIcxTsVTgQw9RdtX+6532f/VQrRpOdIV
oXPfpK1DG1EmkVBlzOXKkxk3xRW9K0NYUQ72kcBNmekV/3Ifuws5U5EycRX5WdT51htlklm7bJ2P
plgdcd5Zw9xitPSCC8SBoCeNVoFBuOMX8eUCKdvDMj8nWgdK6guVt1RBJm1TWHuDGAi7ihEYr3cc
K5Mr65RPMkV/vCPoa40aKgv/eJQhn7n8uUlZ4P1uChKNgvPEzvlFNr7Hc2jLTXl7lXY62hes2snf
Ixn/Po6nHlTNngAH1NqmvQF16Nef1epmp7Oe/0xKEhfp1ZIfclAyxdkydePeoKZ/KhO0yiS6pxQ5
YjCnGVpASBUlDaWSi8/ESTil17t75KAj3ThcpQ7r5SdNgubYG1+hWuf2Iwe9mfXd7mj8ppW7xyVl
P8kJ0ofIUOLbWS0iSfrcgrQdMdlHJFnLN4e6ZKpB5MFQk+6n0QMjhnTkJwvfbV4zizYqTqlkQlUN
jDFUeIJz9FuzafGRoJtlf2j0o2VERGxHIVxjD2axJ84IdXM3pAOiVca/xalsA4iCJh9PRWQ65EMl
oljZE+0IfeDZeSrslwQ7AexymVCrI3FlF2Vfw0qTIkvhct91Xi3B4qs20DAgM1sK4xjfMCWM6Ten
aDe0fnpXNtzUhnJX3lXs6/iCEGlgv0Ssgrar41XNvH4nOqNx+VXLCtRRE/mrzuIHlDDO/+mxi4Vj
Hy+XqClWNfut5h6wemX0N56b6fEfnMrVnDxbuRg/hIV2oLfTrn0mX2OW+Ke6o4JDdcTn5qrCQcb7
kMWI77lZc+ZoyRPL3Yk36L04pWD8Slo7qkKTqM33jtZTZvV1WXCHcREP7OLuKM+wodiJRjTDEjrJ
FK1yVMe7EZsy61wqmaIYq4unRvdqdYwjoJnvCIY5Q8c3gtJ+q00B0OqbHQRKMH06k27ODSPOZSqL
Nc95e25gQuFohGkG1HrWI05ZogbV0PkseUxJ6h+aPNjujt9dCDTV3Qikyl5FYOujWi8oqUZoKp15
zgDC7i8rbe2Qx8N8MpZesA1pFIAv7Y/NtohOak33ATKf6Qd5DztwYVj8z+NAjU7HKdi4FEGUvxwj
BnO0ehJksK8mk2J5HHlFNZgHN+mzYD7gM+TxMwNFTloja3+hb/mlyvCy2cQsmePCeeIOHRrM8Ey0
Anw2wawKvtS0OvjOzvaV3z5h6SDkSK5csZD7dnA4YMFkbX+jfC5TdgSSwHdIERXfT+O/EoqwjhLa
7hLiDUFiQw9C47YkClZXQI6/9vqJblYneKd/MAuc+4fIJAVWYrZlSdeewT1jalI/rhbvaPDNB+PU
uCSUdMOxb0jn8kK66Tda9KpdTc1EWcoVVl/km1iwvpvWh1FRiomqOvup8KF83oh2EfWHrSQG+0P+
v/rL3qNtx9gF6LwS4HwECpMqX1RgG52rR7m3u11LjGUmaB4Wvo6u6eftPikChHyDE/XBuBU3zWXY
l2vZCBCCLeDxGEeAux/VVvJ832Y99J3JvZWZnWZiHGG2Siqz3gJklwoWVvZcukVVKcFreIFE5+kF
ZQeZ9txHga4dm/cb4Giwtdr9W/CgwQA5LjToKBYj7sPtpFRfFoUggHmeg2ZC06x7WEQ5Od8aUuzd
di3qY1St/HnckkirOi+3WAGNaRHBa5Fwrf+pzV7XWkli0+CBwgy5rL6amcKgUmNREEdfbTyPTveY
BJD/uiMa58ScImJAoMKNVXydV3C3F82KqG8qOkaed0Sc5rrnevXzoj1yvkkZ/5bPA85ilDaFGz6G
cIR+tX66LJEcJhWuHMoDyshNfi0kQ8WgKdya0DS4WG6Px/Px9iOAgfPvMIlFk4B7EwtXo8tCdWfT
H8UvWuKxr89Mibiu7dJBFS+Eq7HTXXswfjT3FNuZ/EHqu0fu29mL1Q4K3ck+RI/AAO1rgnuxoAEQ
kITBjdps4ZjyfLV3D0ixWf/bwbfmDyU/RSqTO4e/5iuc87hlfSuKOWk4zbP/ynPWFcCUUPobKWYb
T2Pt1roCNsFx8VJ6tsZxQqzluLwroIgbgH01o1saGfyh4eAqeGpMQlicTfcuEnf+Gbn7gY9SRcOR
wUOsqQNdMntfJG0NB7UZmqLofwaH+b5RcKAKO4Ni4bS0rMoADw1OnZ/d9e4PnCpbe+xPCB5RS9+m
XWasFUPzGR2emylZxAyDPvtLYN/wNwGu9IoFsMydssDWz2RkXFbM7dYH7rVyeMGXrpIr0AchqW12
5wZnVFvvLu6C1SjKBzRoAl/Krr3l9ZLCDft1Tune8l/CpwG8LWk4AMaZwgQqHqrTjJCuzB5lJtC9
nUHWSj8PrrhvZgLiEPmxVhUzsnXjBiFS3phMbkbDP7QbqibUQq1txGMn3Ztm+x7icAwYMra34Uei
s5ZLG/i5JgnMdN2gqPwxmGpvD7IDTBNS8QIBo8shpuwb69Nkq1cdeGK2mevnLBVyHOwM7Gr7oGxP
QIhYfTtG5xskuMCTB+hJVqDZYYNRe1lfYMyRTpfPHq1u4zGPYm9pjWBD/m9pQUr+X9uUn8fEqkhd
yXa8GMZGQJZotb5e5bx4/Z/e/3XN3rUeYow0VB+RjHVNJ34wjSpLrWFP62wqinbrnAwphvm5aN9X
j9V8S0t7eIfdWD8yOSSbnUrx8/5XfOZ0rWWLX7m7f0IlNKCC5i0G72iPvaWGTuTEITgo5GAeXIgT
X2cUld/m/irEaCoBSyBQTlagV4MgPjdSgTRFzhJoNb0HF5uJv3SNXRdNa1GlC84VAPG9iPo1lEAj
/GLdu5OwJtSO3/HqXzzMlgYMcG0R151ElRZbekJk5+rLIubQzrs+JuSdyJFqPEhl34R0eUiktnjl
SpfW8aRIjrh9SuRUXRYwqIFC6Ss0M4ZhQ7b5b8MFcfqFteSa1Ev7pQb47N2iTwblu0+HXPsJQ82d
k2E6fpbL+38/a6MUS7wfW9cviMR6e5Sa5Bx+f1iQiNK6Q/zB6YIoWWiPhh66xE0lcV9Ohihkt9M3
tsZILCc6qxk6sCzMhISg8VDPy6xrzl8otaWYOdkk9pbyeskayNByJwXm8zURhVu3USmtlIS7m9yE
beeHsOVCeOLxZYqTEWlJ3oTBb3yY5RfgTtUc9WPEh31ZXTpAhlqpN4h40/SDEqT8XIPWya9hlyvB
Qxayh8+d3A/jJuxfbN1wybGkQMpbKqlxXkNbGN5PaVQdk4qfzmd+PJzx48HTAyXjrkX9wmh4rrL0
xMmuMenRSKFLL3Z/DBdYhYCGQjYPFoKGkTpvGMZDT80H4Ks/dG+HeiUsxYr0Zsu7AWTbceYA8xeW
Tp7V0La3tv4xnENVet4qelQzZNGJxX314/E5O3JiuKpYd7Fe0eZjsAQeO3NlKePaNjSlKu30NRG/
DdClLR6iW3wLqFDRsPwjVQz1nTdzV9qF2Dav4S8EtcE6AaxZ1RveW8J7NGxv6eF0e4QbD6Ac8zr2
RmTMvrqPEc+zjvTMFKwW6WU5EfNW9OA1FBOzPXXH4AY397TJxuzhDDAJPgYnm1zXkGrWbTZu+wYp
ljVYwF/nYJg6VENG0XI0QjKNl+AEQQiL410Hd6hCHVyhizIWPY/9Yqr8XBD7G4lKydmSu8yCXj69
wuHyHLaiZpfx4F+Wsbv1vDPgyc/irrUs2DAg6UJzCIahiFWJ9yKV/UFCUeybHmLBbN331KCIfN4Q
L6aRW+1vLPcBpF6Opuphg9nIDCr9aVEgDfT+ZY6VhNYrsLuL7JCqtnBeqMmZMCXQyFiHrVsGeTZt
VFF6n5N1t8c922ju/T4cJGYjFfjCAedBhlIy98ltXl9rGlnekv64H/5+ajjYXYRnIZ826hP+ij02
QJ5FZrcYVLo+YSdwiO4SbqAX7iJEUbRELiNnQDgs0NhX/h6ExdjWsnzB9sxbgyOL7MOf8KxF7G3A
hGuN5GhNYKIc4lU79JIeYP82S4CplV8pLSudQm2SkJ6xKuHNKrOMy0sHBLnDRjJLpE/pTB12zwrl
dW/7bahn082mMUBH2DdxaUVqF7s1kxGGE3SvATBaa8QDuds9ogyWk/ROJ9m3W9rQfnAHCzdasIxI
Iie6HfYM2kfzRRfOXH7vHAVEfcMW42eLI5BHqg941jmvQCSw3WaM0B0HThJmLG5Jcywc94TNpcx0
Yv5fOq+BiW2ZbLj3BS3LxGw9diCqeeOZA3awNSSQAdQdca5oVWhi9r5hLHAugakKHIWrB+Sgdiao
SB3rzLPFKr3TuT1C98vxXEIrDrTv3LV3r/liiVcixXN8epUWAVBW8ImXxl63ktzWG31CkOMgCmOz
0IXFwIFgvotO6WnfetX5yu1vwo/R5dr67EZ0M4hRqC7ku58c2eWux/OpPfImd6Hk7gXqd1Xpm8t6
Rxf8gEPpdCHVr7grgfP4kz7oQaUWP7KzBQs0PGkcfh2brUNDkJ9Bzb67rcvSRh0pc6PeK3ILJn3D
M/sWZcJ8uf/U0O3G11CX/O0LZkwJ6LLOh3Ki17Kb6w8/pm+IKiyc03iikX861yO4LAdJL86QJtfD
L6AfM3ZRcfhQXAAte8ZmN0p3qba46rLJy8bl9rgQyfnVLvU3cxc0s1iEWQ49umnjKO92J3Kp8xNX
wN1fR0N8pG/namTQk4bfPnBcYSyK3+BKN8jniM8PWIhQFNovKBv6G7oOXw14sHM4Jr/+CwAvCSgd
KdCfNOiZpuoYsBWeAN8cwStyruC7dVKXlcdVVbUlENQxUnnvJAorEzbJTehJX9wmDfndWQUKO/dn
BvfxQM0QUBgA1i4AoQWrxMirAsBsx8s8G1joq6tgq33GyVBmRvxl8ZMmUJ6aVPhRDOsVJzsRbx9S
XYO/XrfHf+YARqwuQr5hKGSK6Uxcp1OwjHhnTi4G9BA8yIcIkkh55oxc9R+K6HMFm73eyGDz1kN6
4JkKEdb4EDYQWVbejeDeTqrdQD29VCXAgQ9ZtzFhd6kBbAP28ts8F+G9oHGD6eQt9UhsRUhKHWy7
UASFSAbtZZFKI0+o5Z8Z3VYHeVNIsWwGAahb5C6yfCq4zN94Py7nRWrtRiADYmJenww00WUoGjUW
ft2Zygr+I41GlezL9Ke4V3A5/16aOFsQJp/7+xWxa6YZ8Mg1ux51PvC/mPaqp3PGU85DFXee+7fr
OwDgNa5fnBBNuqlTOyFwMkaTRj61WmnYVIeluO0Qa1cOD8/ZAsIhcImjF+i8cnl4hNT57pYs3jIp
TvVvcorjYilOHx1ECWUc895UPnBmvJmfKwbZbYGPCE5mdxuYpoVtWI5J+rsaJM65iOdWLG5F3JYy
BGPS0CfUT6eDgXtgvRyFkQtAj4h6g/kN4ZdPFH88ideibJapqzOzblbaBq1wZ3Z7do3+xY0XfCoy
njJjicnBBjCptTM09uOjrGlgE246oA7eHeCwOzK8/KrzQtZ9l+sj4NN8PJc7Ddbv5YwfSoJ0nBCF
9F9vPo6tZWuxC9T7Oyq0T1tx4BswfhE6inekYA32wGJvYrKKSE9a83cSt2DTYi0pCjt66Dn5t0jG
GjLR+GWNJ1DCBe993mDecBnnnUeozqZz9wkQE4LnknUyrW8SErZ6lBNUJ9YRn040XvlzRlbw29AR
T8YW3Lb+TSnVJvH0WyQLUiUsdOG7pFj/wSvazD5Dn8mSyTaQRn3O7+JkAlsm2mEsMG1vyZQfHMWN
hWOsJWuYAITnOCudslvcbWR672GyqZYp29LTy+CvQprxC6jDTbOjavSqO+Z0jede288XhU/neUUs
adCqCxvPjb4WmjHfWkPka/4zX0VYIniAbgETG1jc2J1QtrJhr+MlBrJiX4dgiqaUiMoW9ePzXdxM
D1kJlpXvOqjoztcoRWeOJB8+gm9W5DQ9aJe4musf4svOJqSmcZkED3GZmmdpVIhCmyBpzE/NlEpU
haGJ6P/E6eGyjk5FtnknM98NQ9sHgAW5m65sjaq4DH8wbXYVVKQ7VGrDLEvtHfXN06AezLfHEgXj
Q1nBKAl9z/4HnqWK+8jrnwks9IPvCsQybrdQpahf37F8G0VfoI8gEDFTWLoz3ix1b0EjyeEBp632
/ejAKvy/455R8Kt33/I/UB4o7c4IDwedJ8kdXwgZfE1H/KBuKGn/v/F2l9SzICzDBeJ8qKK5yt+V
R4xN040aJsqrY8kECGzoTU9QrVCAqcoZEcFt44eURs7jUiMhEUTfG5tXFELhaLJSYUeMxrVSrRJQ
YSxUzqIgav/YYp1xP9gs5BFOVOyMW6LqjulKuQedkutlu9ib8Lsrdjxg6cZ7vJd8oCThQKXXwNUn
0xiUoF81l6bvbei4kbdlpTxH1IPTUz9CHlXsBFJzoLDwwMUEOe8AZ4hySooQb1M/OvPTMNZB7Wg0
13qiW/rbYLUEN83M+rUgwJF6NlOIQE29HYUE2ptSeAu8vqQhwUWiemUj0iPACXWvIqMxG8zR153X
6iSNu0pDY6PnDvwc1qoun7e2F4uyXOvu7XnGPaTs/291ei0YrD8fefQmOMW4XYGzTs7SMH6PdXVt
GRfzGg4ZP2onqY37NFKkLuCi9SpSfpKzbIVR1mcbP2nNA5UE9oQtkfgGqjgsovJQaTO/rg2Eh8DY
YJODRJIgFEy4WSDo9/D26x5rojA4Q+7RmVvJuf/LQz4gIWj8eDrYikZqOvf0I69g1sU93iFyg2pi
XNOceVWPMrr3q79k36d8FI56NUVxzPFdg9umsxDwoPezYZ+7kslx+0zYNI/daYidHdJHRQpYfOIm
eJ7T6xegSBlthCzEIwyqpMLVaK9AFAtRU8clTx6r4wU+17V/7V48mPcWvoSlXgp9AgZU5bqprw2O
4nUoEoIUQ0QDG7q+17WhY+0j4EbFJGQ6PpsVA2VMmreAmnBBWLBuhW0tb3+qM+RX6Hd2eGEug01B
YqOxSP9E4W9llB8OYlJQqFetWBeC/9SVxvP5/HkWaWFBO1gBBjVC1zOdhlZVp0B0X9BSekNZleu8
Sjb5RW3bwCDIiLfQ6uMEehk5DbRakZqpeBFMU2z3TvInjg5gpkY3jA/hvzyMpelz1MaVkhXGqcVa
CjwoFriEdbiOC5I9g6KGgRI9m9MfLRRJNMFuneSFpxv64ftVywam3DkIW8MZfXKXZ2xJsyNijRnv
mQhSOEH7tw0ucVZulU+OSwcwllgrddLDq9gdqeCYmusJX8ZrEPeU/zC6kMUclTA/s3BQacULnI5O
GIQh8WgY8Gn7qMfcP7k9ZDnUHwJLOWLL32QaafsWBbQcOJr7SgotQ6AlDkAq/en2I+IKtDsh5RRG
F4znG6S/erBVMFjYH/xFQjemzNcvNPDN5HG3twtDIpv1HBoez2LkNtcW3riYkWPiYL2e2aeJkarn
qNRz+AZIoTbMPy6i9txqPoBt7yYBkUE4AQDtYhn1QTBxXYqFVL1m54xqHP+eKWjZ0djJaZBhoRm9
xJ55Qw2o0DNmXCNuPBvG5LoVekCuXh9xlIxFLJAYoQqKSnQiR8kdyl9dJdIwSLgDw6fADhGcAb9w
SKgDV+c2twGXnrFVsF+wHIiWBw1P1c49rlKL7ZOgUrPnAiEXBpsYhKkxnypxtn7ZHanZQffdm/Q8
i5KAEn/NKzdnWg7QKl+zak+jY37YPMYu2leVe4klhDsx8cAhQa1x4Z98Yb8E0TXgij7evOK44lNc
Mxf7RVX9PrKE2+WDX93E4wNqV4UmVcvmNH5E7F4lcJO5oqoBL7piHq+5FmLgV0zKVPvGTqYXz9bd
WhVythDk1fpWT1De+tyamVsU6phpYM698nhy8UWu7m7gSQEuOrb+zO9oJPdDtZtRbf3NzvumCDMP
PS8cZCBfol7LpAmOKGOQvjD1UQVt6q1Ln8VL5O34Im4I3WkxiCHAYFlBX4hFi6qLCMQ0xeTziOjw
TYg5TVChlcPzEt9jS1I8K/PCEFu3k8wo/LpJ98nmMM0aYObYBOkQRu7rIuLnwMi7k03GTK/S5gNI
r6MQmnMz9h+MV82Wi7d5on84fsMecyo/nC2yMJ5yQykqej0u03mNuBKiDA8lTfJ13CH+sC7gPn0x
xEujEO/+S1cN2poPfzj6L4Re+aUr06kS1I2AoBgLrdO8BnwA+JjBJSYujBKmE9cw06/kMT8L6P+7
DiGAl28kiTXLsGaC1OMch040G8XT/ODwdyFE+e2Vwiq0sPPy8+ozSlKA9+Ws4vcnQmew9XWsdjSj
YGob5kIksh6K1EmLHSz/WnCI5xyInOp8oPdxGQjuH0Y8eZoomeHfAnNi1jQwFDZcb9o3PRDqQxLI
RM1gw5Yz0Bd0w+O8Ch1Blxyaud/7liHv3Cco0Cgm5Mn8rVQkc+/RJPtFaImBvJy+rzQFicJanC6q
xqYFCmOXe7d/+pQ0bAjFuztVkTL0O/IHri5gNtyDYWEZnKUwh2fNF07aF7t7n3wvrY1NyMbSKdUw
YGY2GJemQbc/lM/LpiNE31G2Jy70m3BxZv/aR/XaCFPp+Ngst6FrGHu+8RWvNdQhWzwERd7BTkw4
Lwwk4Vhl/Dr1EQ/Td06GQvJu3buidMsrLQLg98nzYHSTE6UbjLdK+TBj+2sxPxe35QtVfCAk9oVd
bxIXNvJc/gQBRg+oyzWdo9x+6Zr8jQRBvHaKn+OOoNZ+mCLPTqqst4WkkFx+R23C5tA28z1i8/Qg
1znQ0uzRG1uHm2qCpS8a880umpH9Dsqi34DAbPscQkDzRW4ul2o8GrSTrlmlpKNycE7kcbGJXyuQ
+QUduX9P/PB16HaVUwTYS+/+lspST/Ll5c3nshimNlfk1f4KWrPLfQvsZjueuP9kc//KpujBZ91M
gKJQpxw4a1FDsCUZDmYiAC8qyhAml0nOUbl4f6B9826it9yXXHq7SIBCVzYxB6e1WD35yxdntuJw
FQy9EsWKn7MY0hdR2n/EZOhOj8wkREYqafW0DvGeQOO7qmXVzHCIL/T5H2UnEE07aSy4PcH9l9qq
OtN9rXG2x3okpjretxNktqtitnefJklhq8Ff0NPant1n7Kk8FoEfmVe15Xp8N/Ip5i1GfohBQEkG
ouLi5wz0N3GS8AScGo4pK0LUlXLOehQhhkyqih3bWaqZAQ6HpQCeBLIabE2FyCtKxkdrba4M23Uj
e5IJ9mpFSuGv3QOCYrtcFGH0TiSy0i5SzOKzoJLaXXRKoPxwIbjkRRW8Img9pvRsCDFa0He+E/KX
00+Ymf6w3+P1HCl+viSDn2SY09pX4Qbx6Vil71XxRmZAn6gj62rGDFX9R1S+tO/792n5+0Y4n+qb
vEpOszA67qdlRMji5oTLdApgslSj3kbrLEn2k/KJxFlOFy1eyIcpjDfiRrKwzbHbMwedYFQ3kvvZ
hVZVUMwIfh5Lo9Th88amPq8ida0HN4/8WaOgfmEn7t3vZIxdc4SG2MleHBGVdjAuJ7cLgvgyMsyb
wZ7sCKNZkKm2IL1LslGlZLs4PWhG+sUy1Cgk2H6LF+9+vEIDsxYSr7OH+VErCoqNi8HAeVvxv1iy
uPbegSCRcQueLS2Jz2Fo1tOmyI4/Qm++Oc4ThmBHIEYrQbbbNlR1FQc0E9tASJ9FuOA9HiI/FTJb
MqVg1Q2QNoN802369zVgoegfkPGAvGGfc/FNtAMgEIySVuPypa8p5+Jr0g9tHp5dQ61/IA6dmsjG
NP1ST+GaNOsZMOlHrFF8A73sx72FcFpoVffVlhBQ/u/Q927rC0s4n6vQxEJgD1Gz529k2kHXyB+s
tOEqllOXE/nOTZXL26H6AJEGcKC9yB+FiuyUPq01r3uYcFp3fqJ6FNws2mSqJmKDcenUAqzp3zei
L0mvQ1Jx/TViIg9tqI7vvElhhM/wUz9VWnVCdSogG5wF4+/omXtRxnfX1RYrAFv7Km3C3QWzeemt
7o/4WVxy2R6P1ukQt9D8FZ4/LD9eBav1gIOGlbZbDktjcrSSeEFBvHoyyCFuahDTlUdUo38lxP4N
C+axT3GIWjpoQMIIL05pNFl9C7USZN4OmXNPU718S+M9E26NCCVaTv+o085CjZ8lyBN7QTuLsWK+
9acbQqrBiDkxdnD58Neg0kabUrA7rakGN5N9weo/oh3mik7utIf1svejWeOYVIsdLq+w2hBlSq3v
IwU7EtGFKypezMhJNzFgkmWxXKcRuufj9ew3zAJ8bLTMgydOqS91cfHCupA5HUprm5jyfuxvJpwk
rMF2l1hHW5ntwAdInIS8CR/gLpO/X3jroEctaQrAMdG6f5sGOi7muXrUoTj5pRPCpJjtYpQK6bzG
tLC/f+aWhb/B/vzRqxKPE+fVmkVoXegCMN5rOoHgn0UHPxu+73dK5TcehVc+1Bm9Oau8Wk8mrNQX
bfx0MC/Ot9iUoZbokj5U8/LDs3NZdleMQd8xokes7UDFkh7EGzxfTL+IgKIbmZbY1i+LaaGHkq6O
Tjfwh4eTXqzfsrzJOstxgqh9YK4IezmZfpLQNbmKSAe8CYwrdowc8HA4gQe2+shxn2JLKCWHvMAX
ZMbVyc2KrqmuZLDZcDMt7W6PFfcvZjZcK8DRDq1c3ErsFffe+IEHBRxhvz19mIr+Y/oFf9FzVfsz
0whWR5eOLOwkaDrYsPqvYYsnbU/Pa2QPONaSFeMZiZp/uD2k/U/HBe1U8zh9DsDXkl5im42/tZ1P
nRZjrde2CpWuTCEg1xPkx4Aa6j39lqeRkKFARaMxI0GXUFSaw8ocBAOKDyPbvS18ev6CHCmCTgl1
AXnWdPN5yPMFoBFA8aw6S0WW1tYahRiyDasAQj91kyUM6ANbMnozkavWJHauaUbLdMkEGaFAxB1d
43JfEJWQFQ88immARMVuG49i+9mrpDVWFC+3Dg0ikUlhPPJCVlW9oJXmGyxlyVBJrjVfvrVo8pRX
D/Bu1+OJWYEkqV2rJcsdtXsKbwjWZKfdgCxZChdbdGLdD8TthIWGGvrh9ljt+PSc8s28jbFaaYMU
J9OQWUIQkbg5uor9M+0mr0ZmvfRhLfC7DNwxqkpaf0RhS8XllcUZ2gTEY3G/hO59wnUMNF+giV2i
jg+xmfSRn0f3gyrFZubpIUh6Zqs3ZCIofvith8GCAPhdJsqUjT2ScyaBRqH1SgtIM0++B8qpprxn
XiAVcOfjN2C1XTibv0VlMOHf2hxL3LxP7bsPM4EhT12kEhJM/Jh+bJ43R218HWLYQEDKHPSfQare
LVF7AtG5K4xCRzL3aoeGZOMhAXaz1oDd8FuroRtu7EChqoesdJXanAsNm4e6v58rhyJHpY/59Mwn
d2TF1vZBwwVitzc7YumKFMrdkzY1y2k7428+3HAS4v+N2cB1BAbtMAVAg0Zlp3lss0fcBdAKfcM/
M5F4WK06kg6RccSzZ9fKyLOA3E2AWXl1ah1Jvt0WH3A00BQzkSgykGl2uz22kE2Sr09gcrpBDC5n
5/Gjv2N3BE6FquM9k7mii06cTAbpoXzPiAW4VYu+C2/rDvDmvcZwO5NdxnjSHL44Rvx/syZ1ROQM
rxoZTyIzZknEPg0CGQoymzNYVpKIrYaQHg9LgfygU29+iCrsN1bdD4AEEx4UNIt+O83vHahJHe1L
gdLDcCu5y8kt0VzmpjsbHYPkO6hxNiQ5/b+/vgWcW2UwGUEg2H60JEjFWr8T98WfF00wwPaWm1vO
md5j0DDcunHGjRakNKbaQ39PIywEQPXQ0TZ2POsRxadJnBNKexCo++XnW9Jk+048jhCPFrF7YhAJ
tpas8rLb1RyEPmiVuJgiO0df3WNt6ANPrOweDZI8wDZyinH0FJ5ha2kD04NI8pwo6B41CqylTZQs
SfOsrOW5AXwsBznSkQeO40m3fBhr/R6GW6woDsbgBwTKL54KKuBGfd7A8jd8svvm2cpmuB2u4ivI
lPNzScl5z43E9AIlQEEI7V1q2qlqsDrYjB9DzkWTi8djRdfwkITq6Tivd0Z3czQ7RemgnqeM6Ump
6q0bB2yGfBzdTa8VHub73/KdxHjhlKz+A3PmBGhk2N5G5+QPybioFJ6X5Hq08mBSEd5MJhl9ba+G
qtIjRXKrf9NC5IPKlAHQQw65MgY7EYibTDz2SK8ILI8jJuDsk/41JzaAGEvAdRqM9igFnKO4r8Fn
kBwSr9lpGaHTCcBCQKjOlAZEFT6feosKoyFN5fl9x9LOpMuU4ZJTgUjS2Y7zaOFVHmKsbWzbij4Y
UT7Ftb31VjYhGY31hugKtrORwUeKqgy/ma72vOZ5JQyBX0DjXa04pJv5JwYt58YqCD1uMFTXYzlI
QTWpSsepDouX/hcHruuGrzLLu/OZHkLni6MbYqblXOx94j6pctxCc6/Ykiq/8+sjhKIQ9g9anxIX
P/W31Boixl10EatJfnZlztOyfAzD+kYJrDqiwZtcsXP0pvlTNAU5fJnwhcNaxdO/uXgFoTdYDs6U
wTyjvwdUgkBe3z5ib4ZwO3etWHyst7X70z5mgiaVDfBqBzgUh37vVt/mEzYL+++3achcS7OTl+gp
sKb+KwoooX60f1yoe154Gd8SbnJvD5G7TyrwxjUA3W0l34ZppYLGj3s0LCcVVRgK1EDTsYF90iKH
xHn48g4kHCWADmqBDgwLfvlW26vZA14AVnGEQ5ANUdNQl88AyE2Mc+M1hbYeEibDKiBeOAlMmNu6
8/kb4tIr51a2NjqK/+ji6AYXIki7chzgsgen/0boBscCObRfXCCDnnKVrrOwoQZ6gsnchM23q0MQ
IQY00cUuyfxRgpFJKazk617wJcACmNFZ75XoIk2lbo7r2iLY0CtUWqMIrcK81LMmNfrnqPm1NF9O
KVH+BuJCs7zwlIZuxrC2UvHK/8Q8eyyWjPR5Tjf7ChASaYNCai2bNNeA+HTIz31Lgn7M3Or7gkid
/nxivDZrK/0sYV6UsFnGeF2P+x8mPeuqFtJ8UVNtIyXMJ18HcKrXPRpQ0VF7Fg+qA4J1l42DlO2i
VUWHp6V6HN6rC+CH/pqWXj9BH+CDP0qlBPKwDPJqWnD3AUGrNsm4fhmMf0vVHqXMvqbUWfm7q9Sf
eI8FSXXjFR0EWU85xXcU6iCLvRJTNHrjdMgjfyWlYpq/3rmsb7BbN5KnMdsEGjhIqTpyddeJeSgI
DJUu4fEj73Lmq4zp1sKiVqwPYXgbBnM2BCr0xyPNar38G6v2UbDlrdbb3iozKGPglTPeZ8uPsbNR
pOvNEyFw1PEAd1OS6guOFhaR810pDTb9nHiUAzus0sla/DxKVnYyxBccnn/0duLwR90Z9jdUjwb9
T2H/Z/gHBTl94ejQKMENFgoV8QY4L5oYA9wcLVIdnMR47LARXCkZAzoKaWPeTI9bmlmwUjakqjEu
Cf9PBXdyt28PtbYjx+yN6Ph4bWv6qpfEs/8i/GegLLrrUv8MRnGxQ1u3Q+xZQT53YfFRuakvW0Vw
CgRT5ZFHZIwN4pGvVQ0Kc3jUO03ZYLqGaJSMimGO+60LWd+lAbdx/kMMuByhEsQT9EtfcmOCugW9
dMVTRUpnPHbkGX5jtoKmseqIBbxLEVBhow9qCcbjuR+OOgjdGWlLi+NAN59788xEkHD3/YB/RuQD
QOQv4T3mlZ+pKUytF1REkKTFaz5IqIy6vMs3+OZnsT926rOjFgAE5PQG35sUqlxC7q2Lm3V8ckPx
Y3azZwYZNyFlI/RJGcF1XPku2CNMPMutaHEyTNP5RgYEMX3e4yPEjvymrKSl00Dzm/Z5GQvP5lIy
7h7czG2f8fz5MufZDoCIO6Di0Hns8M1Pnt0GudAKEucOnyAalBz3OvL4XrCIYfeaIwZ5axVP9npF
tuhTIZ2SYsZj68votfYz96YWHCglAv8WR8gmWmmawTw7K99TjqCP3g3ywY+zVdtmuGV44YD0ZBxc
foLNwdfiBkAmP4uaAPvNTDhZjNHOyGSoCQnqq7OkHvkDw+0JDbUFfTw9haSEZttSwORQK0z4XdkT
KNPW5sdmvnednZ1oiRYP3gnq6kJ/ZbepgOH1TpwFXN0f1up96fo9pxLgdAXfJ6eFP718tQmW5jjO
EUzMDBTFDKYGmLXdCEJpKYB329FbgZHOuvlI1wPVXiQ2q4iHA8fTuBMhlKmxkthr1C5ag+4A7qzZ
py9YriE/J4lTebmJX6PFsu4mjZFc62XMkcG8JQgCUV3unwr3SUOb8Iz6P33AvJoDLa7ge1a/jywA
Y+2MVuntX33/J2I6epfjsQt5XKS56ww2vdDmFPToPiJSgRvvj14uZyqrtER27YCcj/qhOEnwSaVv
lGoXFjEO/MPuPCY3oVWfngO9YYvTffvKxGrw+/M4gjXOPXrvKH07zNNVlWTejOHoV++zdlDdLObU
J4lcXTzb4GkTcEe6DXhwjRkmPZd7qnor5PUBvvKQOwpKDsuOMqaE+l1HlP6smGXV0hb/pFC1CGy5
1BHPl40H4Xnzy/acXi+KU0Yd3HDWrfOHvXyXtzW3lTuK+ZJHPZ83CDF/l6WV8+ESsRNqH/dx+J1N
1cX+N0Bdex7Jl96RDyBgv2zi+UvTtvxFT5g30QXjAbxkmIVL9Bnz7+S4cc7NHTGcSoXFMj1vvM0K
4K+LC/8z2dpSegD4pxr+h6igVpy35g+hIXNLDmPEd5xKhhFWEhn9LV4TpijIaElZVrfVJiAOBh43
GcaXVwoke32HPyy7aXdSNTrrWN+dPqzQ8FO/NRa28oEjBoUjMcmq8DQWeWswJ4mNg8S+4jZVAXTs
vqOw+nhNzeUmdkiwXn5gqTwrME+b7ATYTcrP4bnLoaB/V0sEldLlK8W7ttGzWMdPDlWnTN1NcBqb
y96NY61gsbf6Tgx3h1Q8/VvXehixSGkdZ+dEliQGG5DnRqHhwk3sXKJZNm1VERJWn92xwCt688fR
itr+t5QGGKAk+1a2pyhCfnNmTq9qWY+ZfBbd8raSXFaj0Gwu0ITbhfT1bis4LMKjPdkkOfm0MQIL
AKQY8qUAxNdmxlBXBNItQIsXCb74uDxT5oj2VIMCoqPEq7jOXsn930TMSutRHlHymkaAZCmKyVwT
C3OQcd/Z8rf6Y1tbeU3LQYJ2uAsEvXCI2gF0P9Sdc5O7pZlCXiiCyrYS264dqxKfFjSzztr3ko4u
eqvjHqLzplsejbS4xa+Y9eiAbvV8AmoIuI0yObWLS8mQd5aLZi59RbPDetni3YxQIECum8YpL2Yf
NVoDSPfIB1GFEl192HAPh+mbqYCe1vlSXatcBbR/vwkAFiiR+aefae646z4KQOhdolscTppf5Igl
9GQY9nmNz1G7HJXkvlQCTncjydXOF8bY8/2dxT4evb8f57cKfbxHI4nFPicDHAAAhvdsWq6of25M
Rpwx6x6Tg0Wj3/ZMiTzyLX5TJyOLesx4W7gFpYxPdKDzY0El3Sm7JBoLm1akX+jjQ4xHKrlyDpnf
r8AvCLm/wz2eUkpr+7aKxiMGbUm3t7ZdatQLz6YxyeEUmOV00TNA/ptyNP2+Vmr9n/j5cgqrFwT+
sNzQ3Y+xM+2n4Cdko1iV1UaFh1jALYKfSyth8YV9/WJ3VgebS+D5l5RpP2Gjz2nophfUK4UNJQBm
2g3ASgi2mpbH08u850eODtewRso30xcZMg0WanVNjfz9Ms97AoiOXoyb7IiZZquH63V/6HdTte8a
btraMvTf/TEEMJ8PVPcOxbZila6/j/zNs6C7aOiy9QuWpTxJZgTgLk47u6Nd4TKX3iY3hOHHARcQ
Yh3majM/fXHa70SUEcWnaO9ejPjIhAzwcEK1GxTuh17J4A28ZV6vIpJDOQS6FHTgBCR5oW1YBj2z
b8mixxFCWRotZ01R4+i2a2107Wqp+f2pobSolgCD4GBkAbn7Dh6u+BNPwmtQc1hviUrtxqSLz6d4
DY32c3qkbJha4AF+AZoA6caTNokPeryNyd5L+9ljrxCn+JuX6xxy058oiiPAXA+vgKSetTj98WXj
fPYBaTut6X+Oxe41XVsbw7xW2IZXu2ImV9vguIB3lf6Cr7QfOlXVtpOY+g9Sa0HmIjDR9Tqm1iLZ
jDudAx27P2BXzzclOMhAx9qToOIwYJD4NKh+AueO5eGzVu6yocZheZcOYcGkY4oPa2rSzi1qvw6G
Q4XusIEUdsYJnF/xmpwCIpqaJJ3DWWzzkq+xqivSEYWZv94mCDk/CyoiVrauOcc3Ax51v85ZciW3
KM5WbLAVIrSUnmA95cyRin6NzBzCT/aLD176xqwpBJzbtkoFoTOOlfJxKJ88iwNbpJ8DYw3lmSUz
VMlZ1pHzi/kKL8O07eSDCz3KTTYYS3C0Ker0D4/IfOaKdeZE0Oxw/GMX/bSGPuwKnyemsrkYSCE7
M6GNeYGZJkr93nNxmVLhfyxkG3hWkXYWAjXAXp58nxUoOmyxVByUPOErD8e6L5YfQ+4GWJVheECL
p8qsQ3qCt2xBXlQ/0BkJJ+prTdTeANgpn8O5pvcRwZPRzx2nvyxDlIdrfYWafbKyXdYULRoh0IgX
ozMgUJVeZBwaJAPykyZjodJEb+5LIqpgeV9HJZmO35PuIWUxoNqXRe8pWLCzQRytg/+3zfzM60iC
0iSauNRPGx0/jyzxA+dCL2yrNjZ04N2x3uOcMMJqZN0SuGmuSoNEITk/ufIRle4lK6Q891RGl9av
QBTXLs48rzq2LYfdNXpzMMcZC5GVLtH9aPqYptH1ftgy9w48ywogsBj/dHW1sIsMVAcBhp1hIwVf
GVnlXiVIYyUCoarcLF5aesv8054C7ItR8wRSbclRAR6K6luaocxm1w5cE9B155NUcRSIclYzUZeI
GdFA6SF1PgWrzo2SNjMDR03UgCso/8yMcfZMLTH1nro3xfnHT+of15UY/2zlc/Wl97YN4Ip3XjAD
dhmSRNiuQG/xZwHvIcHh+p0mn+Ahkg9d/riMHhNuSzA/dWgInZwnYNCXqtfZSk56xA7UDdfi/rFe
lPLOAq7mbSGXf21hrv++6QBO7K5imdnx6QRZsiflTpiq3NyCYqAPjE+17qUmGEZ0QksWNYWo1jDy
YWWrEqh/o27Px9XEl9cRWwCWSAnZiv9ojCBuw4hBSqb4Azw7yaihrdcGr/NxLqrBr+UfTJD+Z9HR
jO3faVPFgju4WTSKIL54ONkFrE4Wt/IjTLvI+INhzLAgP49jCxmzGQVBZNyK4B12s/kd+dPwHDhz
6YIXLeR2aRX92oI+1ObKNhmeFdoT1z3RIDNNs1wcDDUEUNccz4bZ1G3qqEc5Ji7jalrLgJjsKJ7Z
V/cSigODn+FCVYfAqtx03G2cQzPNTar4P/1tp2RfzkWZtCSTYHT9O35O2rYnQwPfv1bBpHDZy9BP
Pm4+3KhxUTeLWw6N+K2MQA3C+LtWt9Nw1bYtcbsE276KEAI8GKc+1Iv+2yNPtvDL4iEB9sSDcXCc
905+6zaypKCYo0nefeTsKoIALovhTQPy5B5j1OpDoD64nvw9ZFcpv8l/mCndko1cvr6pMTfBTGhs
voS0XswpcCRMEMws31mO6xS6Oplfk4puaEt7M7oj4DeFuAzhiMA6mtad6upqPDq3i/1H5ckIk38Q
RQbUv64egg1O2oiaqMuAYsTyhtIwWVRHfM1w8edpbz2NIHeGNhSihYzDiE07Ic1Yk8zCSmxgcfQK
SbAQxY6c+Y3Ni4rKRG30lYLYRraO6hWXkF5pfkBCghGdvALbLCUctlHk0EK+NC8dOlW6iuCRfIE9
VND7dXQZRSfiVP3Pq6SfLIAhulBE52zyTbRuvpppMQVd/5btonPLVZvT8WuaIVL/tL4aokAAXp3T
vw4qu/5AzI6AXXB1w6aioe02gOqy/x3N5hEzAijacOqAXwd8lOhoYVn9NxFAb+YlUV25eYBmZR+r
DVvvHR6FFmT+1MKp79/S/FHYVJsOHRNADxu91x+31jpOkXRWzESxboWGRhjYmmVe4XhI7eO+Qecg
Wl+a+U4WQ9BnFj4R+/HrowDGXnjjh0qqT9MQ8F8+WAEk8TtkciLXIKcn1dvg+gU4SFGBuGuF8R7V
yZgXVbiXVYyUagZNEUU9MjP36/+gw4pOyKAAp69ImjkLG7kYJHCfmIJKCUpKa/87F6IiLEH7SaGD
h73mJR6Sd+hNaOMm8qKko64sQXdak4CBjxGzmgLm8oKhSAzqIZqi6bZnjgUrI7o86cQTjf9u6FGF
Pla9QGvhAT6Dji38gAza5bbAuKbi/y/6srSXaqDlaL+E420WX3TLtPaBSS0Hg6RtqJjTcZOgiaqm
TkZDB9jCCnnRW7KT1C2HIWLQFNiP16WaBsSqWWzeOKoFIEkYvFaNQqSyVEBoVl+AigPADEA0CCla
X6ib+VaDykKtMC9//8N+tTR56lMq+u9l0FpIFv8s6Y/0X3ZVvo0pgLB7YiNp8YeLhZgU4mQghBMh
BD3I5G75OMEEESbjSL218GUcYwPx2Y+AmfAy05r0+UDWiV5mS/oxrmuRqKdiy9whu04BwiYQsnbe
bZe3voGpRHbWHa1flyx8dKF7tgv6v8z80ajvJUQb6+u31qyLnf8goMC8xXdoB6Tg240MNnp5oORK
mzu9+lWkC72ook9GSPMPiXu4dP6BpJOxRVdm5nBxWKpV2c1oPmrzCAXCrgkSoQEgAyDsgb6f4yhz
yzmExbbq2mwIjskqLZosKHWTEf+0tNCYxx+4UzGdA0KMnsVRtP5Jmn0ogCddZ9WkBXTOBdkQFiYL
GKv3D6XbmedMutu8FIAvHis7ENNuNe9xlo2zFsLAvXQcW93QdriZi02zyaiaZlM+ABp5q/FaKXQg
4intt/hXQKzrlkQU+bg4Gb5VbZ4a4OmeYoMdglBgvLX6vN5fkT11pQ9Kox1PpK37Xdwf+isHOl/V
N120ul+M7MyFCNgpjFcD0lGIcWCXHVpDGReKMBf1zsyi1NVE5zo7j16+l6VmafTMK3mOfHnD0QRS
z94a9W6yGXXCkd+UEG1gC047x7YywZPZ7nEFFyJ4a3mdLKTwJaNtA3OgtFhPt/BjgDnarA0g6ZCb
38BeOOdpjQLEzXGzZIs0U2XckLC9YJU0R0KyT7oLeDJHsoc3xbMdZbjpi9SHndK1ymmWObtYAlqY
Z2nDGcYczebhgY1j5HNpOQ90IFkPbdQuNVTnFSTp5Xm7WxCA16V3WJO6O8ZShJcyllRERA/TdmJ5
Pg02v2IJsU+wWnTZIVmK57ROCXkIpFVxjUVPUuSeLiaJknhc9HpkO8UWP03tEw/jsLPQuQAyqpss
z0zdyX/R5GdRP67eee0i0vuf/Tvp63xxcTPoH/jrDVPhRv6VmQhQNy0KATG+EKPkJhsCkxKAU3WJ
XI21g1XPNq1y3sgnbNNDg/CjmOh7vfd92nIpnfi35a+FBCzCXBVhlavzrEm+w0N1Sb+JA9QpppEJ
cHnxg24lllVQ+GfzF0JLMckbssh6QGxGa+Cv0AxShQsoiyorvwZha3+sHiOCihpwBXFe7QCuxJ4L
hXr8VzkpkiYOsT5NwZa+lFcwfWOZz+2kcq0j+CwPMpoeYkm9Pz8Me6IIhcF3mVils6g4dZyvk/DT
YsnieJUQ1EV85g0rXYSIMrMZr8LnF4ZLRN0QRmD34E+HrDXNVGpyLU0m13grg41jxnBWjSQcaoKA
/kY5DF2n6qsKhoRSx0cVRfLwW095Fww5XmbeUmX26WRzlEW61qQd2xc5G/Z3nHEWUgkUgb7nMfNc
PAr+v58fniUUA6bouTHS66IKeysjtzM+GBLKI2VrcjToKjR+NPt4rCSgTJtVwP8ak6DDHSznPFrO
tcaV04ytAdT6UKuJFwbLfNdkvNmY6A6dietjbJXK13GskkYk1Y+cvMnmoSUzuUvHidbOoP1pisIG
gHeAqukPVvza17Vpvtj/uMD8uPHaBJNMjE/kx0WPqYL7A16CvgHgvuGHsv+doPWSIW4XvBue7EU+
MCnakqoml5ok/akdJbiHgPU18tjqKyJh9oOuQn1rqAZw5taVKD83SCpPFcypP1pnpO2AjLzLNW28
3v/XQDm8os/cLgKQgqgSu+sLOmVATzvRtrvpk/rgT102EcWnk/6i7Rityad6A0JcZKbhoUb6MHGi
GjgT3DkEYdNjhyjQ5bdOv2wd44UdZSQ8+asQTQUF+IOHMuUhnfHlYXtHHLb/36px+TIPa8Zpdw87
XmbqpY6FmD+nfJi0JwLutfXKF+26VR0GXptJ8InjA/BL1ZqK8WOhTM73IYXLOICoHnZtUzXnK4h3
wgbqA4hZqRUgMTwky8qfJZAscoqwKaDmP8WMxWtE/GEmuH+3i1UeW/lerQtsoG+7r6fVBeb2Erj7
ZfNL+6DUcD39PsN3N/b29P4Y3wAqljUdI0tDt/eangKDH9ZToT4ple7JTo2PeDiYdfVH58parBRh
74MA3ggzpq8MGk/evQdwwZEzZ2FB7Bfqh1BRtIfS0Mmx44X/wwc/9ch4OeCc7bBWuEGCjNqL/7C+
O+S2K+LRciXB8xgNpA/rwN3cWbT7l1PNZsfHHXKCw+vSDpkUEJsz0l8XPv3avhzEtjxBErtVrk39
7WyDuaPRo1Hf0a5nxy725vCAeEC/HcyiJfuIn3G3AmS0vnVEhJk+STryQ74S8IWOE4bZx20vTg1F
WzsF5TP5MbqsaQzVHfXLBl/REdIc2fA/zKtOqhPo8MSbh0c8k9OhyoRgw7G7j/dpKT9lj19ptfkD
+AAeVYz/fwT6JfxE+KVti2JgUH/6M5aPZWgI4PAjNNge4n0W4s7I2PwfKuDzpvozmwL6jP6fKg+h
cE+yAZ/vTjnSs1E4iBG2ISqxmxsgnW07Nvg7hCQsxjKDssFw6Pb2VfsTk/5lOlvMuv4JSSiaBF6X
fQKbGLs4tNuoQwxAIbN35FN5ycSA+COTpu4c/dd4zwcT8tqn3kJJIn79iv8VoMsuUdoxdVBKlLKi
gljfX+xJVQ+oJEv3VYEL2P7Ogi7uvK3IstUwhVaEejKqKrL3jjJq7kVsHW0OdJO47UmY9SAjA5aW
MUCH2/XUZKtuiYrNRzJlozvfCCYYfC2hlSGzHE3nEIWWNaTrakt36a+NfsDMQgqbjpiCJf4qSb0+
900rloukOXQGVYzoDkUIMc1vrw5tMPrKxTXwnhCOVpMNdZc2zQGGvmzCArTuMuc/JgxSsukDpgma
YxXgTNeH3oKi/6TLkJE7hW3SFQjxghjB2ajgqit2wxyVNa4SJtCYOZE32agYpsAi8vVMtBw5QRLo
J4cNd3gPbLtFA03+kmOQnLc719CYaW1AopmwKzEs3tr0+aKZGPIkXb7gSogpTPMwJ0qNsKHX0eco
9pwiR8X6LZLxAU8zJYOdJJOi+PggGFxyz5aVqldfo6Evf7PYDA5ktiqybCd9Aak0f3R7GbJxC5GZ
L4RjWxDnS3cEXkO3AUueOe87Bz7cpSmE88KAAM2P6C6UsEnEAqnZmdDmQ9kTCQTqThaBgIyMSSeH
X5NZlZLPm2SWXhuyX37UEEmpQyml8BTyMbclewT1jTiEWmpgY0fI7VNyLoIwLqa/9ZB5RYou77OA
dse5eROI2v3JntGqZ3sA95cX6R1mTCOBALjzD/JkAZZsuuzR/ctfQfMLQvraZySE7BeIVMdIhRzg
t7JIKObzyjwlmZV84PbiG0TSGQ98VXp5YOc9kZ3SKq2bcpYKpJd/Qsyd092SNviy8QlMOlRYP+jo
mgg0ggZ3XtjI7BWRuGbUzSu6TyUauNWzp+rB6OV3KZHzYRsqInWxlBlB65rSMvtQJTX3RyH/1Ecy
SN3WjsrnNJk/B9PsWQlMfJtt4G6qOi54/wZF55dYMBqMDXlQPq4RXGKB9+euzVgxgDkpkWYzSK4Q
Bv0GcFyvL44JUPDwrtBJ6lNVMvxrSqrD6FZ6FWJ+F/9VEn32BCOszuxksudYXExcfCVHv8HzulWo
R/2aZB2fo8ya6Zci5OlLWYVOpkaV26C5ZctL0gfjwp0KK8uMBwS25f1NMbg9AKgH2DqylVt/EQ+n
S+V4comTYYyGhWmWDxzjgZHcRIkOH21MuQ6SPy3zh1nqsROqz+speMAxpZnQxF6UINil27plxiL3
XicutEnfEK1kTm+U1wgs1ZgW4tPbs1AcufYD/x2aZK7fSqXVbrnyhdGPLkVjNrJ4LcP4KQUrQj5g
RtaTOE1NxzjHwge5V/SIRuka53KFROuUTq3xkM6CE5o+5FuclO7241lB2uv9tsRl0dt++1p5aobD
GdEVshoADf7F3/BdTLHkm/QekJcEwC+byujyizQvcyel00Am0XTXeLPzVsmcq7jdBeDXYIDBj+I2
kYdGVNwJpr6itoz3u+gTn7nqK633O4LvKlLBFib0hWDwbejlN/5n14OsmYNijari3Drq9hdWzXnd
rEdRcSQGjqMBbPliqx8BvIxqn0L+jO10YkXGwpQDBgXIZRwKtznImPmTIngwReq9gbxFhAjnmQ2q
+x63DJyF8kY/q1YvzF6yoMRhYzOH7p6J/Urwx0TJHh2uThwhO52PoBH2631g/PZpgyoXdj5spkSo
LqtAh45FrCP6RVo1ICfPOiDVQNfIHu0QVDqMv3UNQ8YapL5yF+Lj3yNItcFFThg0OmdvtMX/GSLp
lW5dTpjB/kGQAnGQFY/a77+Mp5esgl5hnM190/+YT/AapWFlT/qzTlnU5ut5Yet9zL14ym7GtT65
HnyEOaNs0p2vSCYf3A/7a5jjsYwZnmUHD8dQRt83hcBfb9ho4FKCa4wLyop4Y5NW7UiqPB6WNgMJ
6yNgTqwc5cOneD1NJm3SslFoOwqrcrFSVLYyuCICvksS6rEFQLumDnQVoeOAXixmDeAJA4KbiHkF
tOzCxi/tOenkGrHXNVtSPsjrRzb2fVk1rTQZspMpI1jGA45LyyvYkMX+z7k8CsRIqxG1nFL8Tx1Y
qjEp97ldLmOhsr0A/6vy3k4fjrfXbHrzvZlSzRtMhNWch3TOxrC6ZSVIFKYqySTMC4Xjy5ZFc7dd
TYSc7+r7f+N7TIfLHO1PxeWY52OU3VqSMRE5fwrxeW2sSBeAN5mYvDxilqHSSQLXHKdLCYJuSUHY
tRbgpAmTbxIqKDPpBIxEBAlEmyIMWnEUJbqVhGqJTEvM7iRlVlJO43LkEFFHtzcNsEJdfUYTMb7J
NXr1Uq9IcyKsFMDLUyatEpCeDYVBVpTBeR1GqTpP2kvTl9vtZ32JWpPS1yzcES5C3uvr/Siiv4yn
9DeHtayShflnlhvEIKqLAJBqeIENBHuhN4le4Vet/ZdyrdO9GXqiH7UyNQzUcBP5hq4zWqfbouJD
jsl+YDepkPVEv+ja2WzRd9p0+Upk/BXAukuI3FKhOPMQHPcTHZnPy0EZJ+cpjCQ1cEJsLaukrvRs
2mx942I2ykUyHZV/Dn4XwMcbGS45LJBouyDNrVbN5jTcUZCSWR/dW84wusl4PNSUty/Kjhtx9zAk
TFCm3TBL0HBUG6KptRAVCnmomxEvPs9rTn6+IthwPOwUMGV3JM0WDXtHyOr+qz+pKaoZQWnuHkzM
gtnkw0A7opNMISsRSfJ4sqGH5LtMrRb3j71MYJ8I1LtkPqyFq7sMocy0DLvMwBLx34lT6DQoe3TR
6dvBGIIjstBQgDzNKFi/vBRJKAFm3E94tXRA+kc6WEvfcMTi5yfiaSF+p1gSM4dSt5Fsb+AkiTM1
6rgSCGduslKiwP4c/fpJdwL5EecRBjP102fr2sQR7CjGnzjRz4iJXnfy4ZHJCHSfRzE62mqskwCW
lkDeh1MFNd3a10/coXNtL3IaDxR4+6kU9tzCnjO+/dqdy95ljJh//o6VCz9IvyUjXEQTjpL7yEOS
QOIyWmjl6tDB3MXZPwz9POslPpRZEZAz9xPkduIG9JpqYggANTFXbcrQY40bgvmc1rauOX4c4mzJ
f7vgHFRpL+OnPsTIcCNvgRIwjP08ZVTSeRmdExCaaIu0t1uUMaqWPuVOQt3osRkCyKZvPtXzwCvW
w3B8vbggfN90ofzji9W+uh10oIEzluAfuP/pgEBGAzaTX1vzP14A11MaogrxyFh8HRut8/258JF7
k0HWRrCVrLlQ5oyDsE6EUaF2EcmK2aNpW4ma3iA9O4l7gyFLy7hdh04gV49iKrLasCFxHO+TMc9M
CwR+grhC8/RmYN6tkWTWk3wc+9q7b3+Fh8hEz9DobKAV7dOeiQC4v8sSxRjBLd/7fhA3yRvrcjMz
U8prWfiHxRhXbS/OeIYeYos/tMjL8VUVmAW0ho3B9LBG/ijUE4bRuFn8+YR49oJnGOnLHtX9/W8w
E9DIYXYmq8VLHwDqDzc+ChgfxhgtIPn2G5fS3kq4TFjs0Jf/PKGBdVpSKMW8/TgSQOp6pCGR3KP5
hL48SXFA1IL5CYjnaTM6bWIrqDUM//1kTFlvfmANN8u9glo40PEd9rzamXPsIQ6m1g8uhgx3lIfO
Fy6Sq2WIh5Hr5e1jprTvw9XrpeCh8Tqm0C6qYOl2aoH7TDdNjS9Jtrq/Pe3VZjUEHFldF78pwDxx
GMKcnh7QKaHgU+dFr0rRKcWJ7Ocj4K10pJTJPjK7SOSTV4lvtFVTQBKzG+qD7UFvbr+k8yP9uMcy
eLUwDgye9NyAXEywK9HrP5AM4wSzuy7QK7CC0pkhQUCAptlPGC52Vl7OkTxv6nDvEPFIXHCQqBL+
eKzp+xEzCX4V7z2JJ9nCJDhffE1POgX4IJMinWMHk/qtYoW8rWzcuIUslvEosM7LLqfOY5+48jFP
LqUBdqORmfiyN3A4ygITkQ0Bh80c6gsqf1vxIlqYifKOXEgPH6sG/LKJUw7axeCJMRzsq24cF93u
Q9l2UL7CyMyvEhLuqDrArq9utsuaAEkXTVM//9nPYRa52Mfxpp/gw+mBqnkzcmCxVH5rRtI8mXL/
OgWVDzLJ2V1tVidCnFbFFIhYHWscIMh2pCpVPoUTqLBy7W420D987u3B/mkH+N6EGKjaUg1JSkh/
Z/IIxEtetyNoXbt2jkr1TS9/Z83EuV5m2GhDJOeGqLTjUB+UOMQCOANZThs4YdVldxdqdrJIdIUz
2K3S8US186SMEh6Xatk/5QmK9P805PsTCOEr3hu90vkAi+c9L7ZXDSfwxQDOtXMBeuNviTuN1zI3
veBSpVJXDRxwNSZ/yxHGxbLf6EhsA9a2CYoFAtIbZpkdpjw8h7oUpbXk2cPTYf3h4KS2PTY/FsvO
h/wBEPBR0Ln6mcl6UO6sRoTBGzhUW7gtn2m7aFiveCDzoPCzlOmdh/Ssb7rWCpQFhZKtav83LAlB
mz6Elnf69NBripWuL6CTqFpMw0hgRTOEhEmGLXGUgI8LNRKGwAc4uvA7tfvwduv9KVlGaVo/92yf
Vz5WPB6sj+YMRFTA5CGSEShmMQksIAj5bs1zFrwZF9zRjIHIzd5VmUaDrd1eBu1NY79gV4ZX44lO
+8+Wvalt4eCKzXE9JiRhhQLRqFTMrxvuRZvK4zhblDb2iXkpM2wIuqZ46TU2rndyQ0FaXhu71QSq
yamma8IDMBtXqcidLf51gsJzyl/CcLgwiNHzvRaLDIjibtIaCjTQMrCVwfpQ3cxf4PwOOmBcKSsw
5IGX8moZ6JMKGEFZxy3IXMvH3kU2JdYZJl0N5j6NKQUpQam9KiaJCpJJFWIpUGtZmWFuQICLwCh6
uHUjWe7FMV+l9IloJkvBinNA2G59lNR/vDGVwkbYicfNzD8i9vrgzZhOSZi9vwiGm3jdbA/dtnlb
WRxsAahI85NSg1hnR46kJy5BNqvoLm6gvOONV6Tz1lnzHDvjfa9EuBqXwi7igZF4TXElZCZrp9Bl
xBQuKth43XM1s/fmdjtQlKDgpwkOMRQFKU/Bdrzla2ItNa43d1ns+Yrsebb+HuwOhj3Js6gRdBbc
ChSsIDCnlde4Lwj6FQED/K9hm0XtKXT3eMXp7Pd6JprLWpB12Aub1f7yTn+Z6+0/Ade37r9ZooLV
wlRo60qfaRukg8kmIMqnDwCCLFb6oxUEWB3k4hu0djkJvX6gnMYFVejhlSFsfoX8X5lWSsUmLsyS
PKbQZIgOZ5Ovff7bQUa3/ruN3fazitrvmI03+1dswC5r+M+8KQ0IcMdfjuqR+ITM0ndZApcGAPx1
PvoSfRnuUAZwlhNSTsgvFye3DjA4nu3jvWXu+Tp6Obv/uQouECpFxNT1dfgFzjo6IaiVWdtH3mY2
O/A9Dsurtf/JmT6Zi1F0P6xsO0gFq9zHS26nVy+IfVp0YG86fklwARYHKQdlQHnw5/F62xWCD3Y7
gk84a5X3RVSg7TF//fP6QTBUSEUUiGfQ61JHai5d9rMoyc0oMACgREelreX1/ao6iqUDN+pjpFPn
HpQDghX2m/gIyXtowsREZCfjVHcyBpzNruziPuBvU9Apaus+ChG+JXSpjEDQsX0gr+Jke5VSrDjp
zetkatAkjGL2bzSTTPtozh0GFBLBTe8elhvMA6jcflmPgIcTTd/KFAbX6HRl/dF3jFyMQzKgWWuF
ZVeTIIMm2muLWNNpD/RKof7lLIZxsMjfo3CfcCOQqa0mmbJzcmftjy2Kr/8UI6YkPRiwVJQIiB0K
o32f1tzN0w/EwO2mBWU626l1idHT4tx5cHkMIff+gJeQJ3LH4pJgWVw/FpfYkanPXAna3EMUcgdb
n/nDdBMuyixmUMbea9MG6g5hKt7DRj0cYIepgEDh5J0IhxXrsMHjL63Z5UuIsceGFM6ARqt8B8EI
XKYewLeNLzCSLjC4OcEcjA+fWFA9cD1HvGLLl8LWvkaXeyxAQKkSEMFP9rSP1ipHWeoNlOwR7c7S
R2xJcfTHkagSutjCscxtjr+x8cy6xOn7G5YpZ+mHJxZ9pp8rYu0QgwHaB3n6bpv0i57+IPk9gEMr
6ePYXIch6QSBoTSp6vTRDzYVHrE/TLXr3mdA+78Uf8+RPiue/5oZwxvQfIyJfxeCZTKRGGIDwYnb
IL1TlZDX5XG4B/HwXgT0loiHjFC7/42lWQIht09skRpyr/aV2aYS35FH1mkw3EghptQQX3Qi0evz
bGNFYKd13WM9T+hRkTbZKNpOdaU7uSS0g6yIxMyd/z8ggnUYC557/vV88KtqHJspjtpKVDcUWaGI
1/dhpcC8LDWblaJYA/ZoHlz/W+Udo3nK3k9xPOEgZI7IW8ncY4uyFJVbEUM4sDH42eiibftf9fe7
3+OStz3YT5ODdZyIb5pvBfgtE8XFQ9o3GRZv2GJScs6AG6Mh0HKarn5gQ8VBhjnFYxAknlkSTVlD
ZVXmxS0vaIam/i579F6/NQ/5cahY68WETDXkpb3TDzUyPFQn12HgG8bUsfB3IkYx0h6Rkj4qncze
ZOiRudRoktqUqrTfmwOIR0waOoust6F1gB1HqOQXvlJe8jkUWTPYh+ML2MZCBaIdiE68wX7T9gCd
pDUSi++SNi6Mq0gVCFNQKWHNqOpz0cdkkZTsRXYjh9o4/mikAy3kL3PjuIpmP/MqKdA8P4zSKRxU
s2F8vT+8crZTgYHuSi10LBCAk9/nghPV3p+OTvXniGBQ1A6Onb3lhSre6FcmiHGHLrk0KrrkDioQ
7slY2l/a1IDe4PCVywN/R+EXePjwHOx3UIcDg7NlSxNf9vjQOnGq158cYAU9s9N1kx/pFudEukzQ
ie+Gy1572G6oZtHflgiajZ1GhdnhFLuUR/WDxrXbFDhfH8DLQsO8wCFg4ywUDIN6A6Q7mJbU+2cI
ttQbg7xCdtQsQjN8KHTGMXan7zSNlN44BwfZqjdOqFpO1RwAai3S3A+7LVCUzSEy9KjM5eGrj/Jv
zPlNImfRAsFhG9rHsL0aaDUn3TPoYfUx6oXB38jQx8+qSpCYMA6ffJBClEIdLRh4iUZYAuWszK07
7A8CHLbL3vgow3S8IqZA6x26cbk6UP2a2gTt4bHvMZkgyLXYsJThH5/t2OxvxgPWREzERSeCjhYY
UZW5lLRv9ZDAl1M7l1cFDBlxqyvlDA7OgjVH7LUuNH0RqZuq+fidtWattmTQGcwAZFGx4n1dNzW/
WyGp5Cg9RMmQRRuqiOcMp+IRRAarHLDDc0n0yzGZkFgSvoCJXzuTHyz11btSUNUj68VxQUGDGxMe
GfZfP2baO19kSjskXA4badO58RtlGJ2ey5ZTYYolaepBBAdIRHDLRXiXDKombjmFOih0C3mDd+xS
BqbOqse4OY6TWvcxuQHMzbRViILGe/OKcHXOyd9bhBlhtX8bHSu7JF8p4Sy22sEa7zljZwArd2YO
numydbJlBmY1sj+wVKdhPVVeyREqE7OgJiM1t5RrcG+2hLJAeOa6Zu+8qb8IUp9+V/BgKEzUbbvq
0TgZAYT6kY4MPDHGQPHcN898KH9O/uR/QlziclZDK+SCNmfj5czl1eadqQgIJXfZfWrm0yD1PPhY
lmFL1bJxCv0OybV6Gg+hAoAFnUNbJ3HvjorxqNujvLPe7ntJsGi3irh3OiB0SWRy8kyakxc9trBS
BwDnwAhUSV6naBlWnyeS0F+BLSMEZum1a+yMwdnKQrUzmtxAONqCNRM1zHBjbH/pF6LuuaaLkcW1
sip1Sypy5b6Dn0bqfKnvP2S0UybbSGeHIZtFKMGwvgRLiNDBmQO3MfD7XIjGsn9cw69jHyQV+mmM
8Tf3zPM8TfhpK8ElbR8UXve9e239S26QM7529i4mNLqjZeOJzuEiYomcIKwZlWSlTn4gMYUDU2F6
rlbOQ+LSyvcLFaG315tUEHK8VVn92vomKWvsK0z3SqYB2Z3+/8lhzAwjnVQqz9P6cqdMuPtpfXeS
TfhJRIA/MQXRZBCV46jvqZoBfdix8zab966QzSgNKdLcKSmRkYjdWrWoN1Z6N3iDMSWSken4WTbO
LVu1xrYfRMayyHsw0JMXQ3yZg+8dxYXmaa1H91BD5XmbsUq6lbFxeX66RFBa329d7SWnqn/GsJKE
aVF6LaRDWX6Xa0jTY6FS3+wkJfbFy4/mzbE9jPgi5ZKSZB4NqCEECaYChaYVRSBpplJSW+pXFJm2
BF34+XRDeAy7YeTbtFYARbSYtl2Feizku1T/4+cKVnzsWdbcM3PCgczCeKHXW4X2QCwIMPVAzLEV
EQSKGWKDh4KEEq0DntgLbflp1wOPsBmGn3aolgJ4ztEE2fE5Rm7FbZ9tUCIznR1CMnenurJu8Ibh
ZWv9gJK+bgSCLgZ8dL7Gki5P7O596mWwKPTBAUT3tpxP1nDpPIFKegPJ09yE2rpGC79SrwNk8fPX
RJZocB7ZTOBXiqrjpc19RQy20v7LairsEZm5DhsbNhtN/zofsaewlkirCczgD4xrWZG0CxBgBj78
+w4Fc1w++xPz7AJ/bGdKtHBg+mjoug2kXAZFfcZAxXTKaTMxSVvM0wzVza83hMpLtPKOj0F1g9Y7
nU5aUP9IpwlTTeXPXrNp4WM1085l39DPIWI5ObPdJ77uU7u+YGuUp2fMcFIz81+oUr246WTqoMc1
QnazaKl/1K6A5kqihvsm4fRJapqUSkxxuZrvK26YGo6dWl/hkd7wE9ixSDNS41jmvz24NmlPoPvP
3BPdUdyB04FqjUYnOuRIFwOmai9UvnDxAKeT0z+z/xmpUySE9jemo+uNlOwp1id4MQjcm4DcW2Td
1vM+POFy144f5cozC9bLrFk+PxjnmU+ULQ+7ben9nAQQRrLLgG4ATZ1/1Ag3yPZFejfLvfgBF8c5
EHWwUyxzEizd6d7c1euDCIuJ8x1LzcmCDxY35QPlVFC916B2pNdASRgM/Xnl9TKXEYBPnwr3WAP8
6aIKmDGpI7DsjvSNzpwslOWnaQ6PW1hP2Ra75n3v9CjKdGCXILy/xTsPk5XVU68w6j9h11gEa2m4
xBdMfldYbML4UasoK6WP+DBWahJSgWIhZDVkWpqY5euJ/7R3Nd+xN44iiWUWJUplBDrt+Vs70lCM
gYsgabDcYNMcBFlImQAmuAPORqkXnlnMmQ2K8CUWZ6UEUxq8EpuygfNcetr1nQ7m1eFj3yOtbLJQ
JMkd9BZouEIzgueJg9Yb1x4xc1+XMzo1hBeXjVI9pKPuPJs1VResoblI7tCE0JgHNh5txhjP4e74
kAZOANoqiV6Em8KpYSnGMwAs9OVCR6agzAnl61a5WPPdydiATBUlhYLM5oknu2415U41ymLLnT89
sUp6s/NcJsjLxQPlg8BrDRNC/4xTG55avq9beXIoELHnlMI48r9mcQv/SmVrz7odkRgSbv7dou4q
c8j+8e2c6lenDTt5IyGieJdeJxx9jmzAkBCC+iD3w8GG9DtfTDvvz7yU0ZEuQ8mdUdbKNbVgv0Pl
amLc3s9/QZgH92lDhpLHqnk71p73TIovOk5EvQ1gJfwzcnTMkRzugSEg0Br4ktMcVlhQ4UMkJXKN
tYGbOR5lH2KadaAUrnQQpcjgEtVRl4nQtf5qkHbjL1kWYerYxZb/ooWG+kggTGRFRl6648Vpo2gM
sEA5CEw+OM+bGL1owT9wdniF3v2iKwQw0j6Lx1rskcV+jGjIe1Guy9zYN4PP8vb6SZizXZk/ETZ4
NSKO/f6eJpb3MQ5cI/lb1+7KUohkeMvXuvzoWii+gUnkrQz664NSJx5JVUBs9Ae1KuZQG7DVscEt
q5HvvJMAwC5bnp8ZrBfSctRizkMPF/rkwuthJ9qMYqlEZGvmC2677zEhC5/ughU1L1gzZkw/H+w6
psl3KNzdUT6gIXN+05RZOQ4meW/gqu8j9a748XqE9EekojCWf98TVgbji9Keh6ZZlL+YM2/Ysiuy
fUxcDZYRMDzCXAzgV6gaYJ7Ap348dZmqcmlsRANNrokxGOEpfMmF3g878m+cMlEAnnPOOkEwKtCh
8h4DwzFbknXiMdF0VwPFhFGU0IbGw5XWLWcju2a8g0XeEfH08GXW/I5212USpYZURvEKxiOjmGq7
wh0vkCbqsRmgehZr4VHUspOlh7zZhX4POaITD6Km+gz/f9pxoJpyk01FpSBx84Chav9g20sgQWZB
dML8vVZ2ERfUI0dfW7TJWGEdW4+dRFdM4UOeRM1YpPjJNnp129nNmv7BR6vHMw6BqlDHaBBkDhlO
rzMNMCX8UXed+/BoSDqDTjTFakjkcZYt4SPXa/clHGJJvNMtTda3Ahd50lZ3iKYguJtXR2/8hfXj
ZfN2knzoZEouEsKcfJRUqIEOlcDsya8EP4sLqf3cqEQ01tCr3XZxqzW7yqvueMEtBsn/wcONUfih
GTYg7W3WpjJH1LkBUJ4inGm5pH8w9ZgOEIu4u/FmWL7jXPY0vXdF6oXHjzY6/hMknS3wOgm5du7m
qek7jIEC6Oo/4JKXJ2pQBur3qFXgd9R2w9EN9GySc0ssxZBXD4V69Lk64BkS7IfcVcXcV1NA9+nc
IC3IPmrFVyffKOEcsMgDhuCA6hZDKt7kA+78hMU1RmrlH4M9l6M4ELKvuPh91UB0KnRPLn5ujz14
AqXSxiJfsa1vBEs7Mjym+gyAbi9jGbBd/mbpQcMn/KAM+d9oDSTmO0eMGuJmjz+Oypq4407qxWSK
nmnZAZjsKoYBgUCG0wAZLwdxlDKjp9L0lojIjFreMsOo9EQ7X8riuOueap8rqHor2SZxd/tckmJ8
3OtI04ys8lgtPzBlJe3KNPT/Ezf7k3FCuaOerw5GQJQ0oQmwujt+bMRvUe5eoCwcP/M1om2Hc9Gk
U0QDKjTGCOgy/Lmcf1gPVgaUhMLakNXJc8F+1zK3eFYd7GdE0jDHLVDppFeY2qDAs+mhRsuqgqQx
CShGpMHHwamETYhnUZS61TojaznCUx9eUrTe/F+WykehiyVx8B6xCK3R0xWzNDkaykg2e+Ue43AD
196XxuPYGRx95pdVUukQMcNlupXn2u5iQ0mWkLHVOL+oNrr9hM0QJjPZwfmS4hGc3hXFYtNzD52/
cT0fxTxADt1SqHCTWE9ou3qCUzanOHMd1iXwEOlC1BBXunSBiBLzUvu6FKKj2yD5KJbnJvMQF3cg
n36AnGIjN07CztvjyLSQ6XDlq15pzZT0COTgiHadrLqLKa0pzJqB+vHoFbzLRPIzJ63I/yp7xCi0
pX22/afS97o2KmATG0H8b91G8d88Vw9SkCbIFEHGr9aNqCq42CO2dRgvzYl0ebQF8sXokFBveWrz
9QX/LyzMS1Laakd50z5Yi9G8EC/Yh0bGwayQ8NOQURURvzpjl0fp8FgAKOOMOGpmO/E1as9tkqKo
yhAPcYJshLjc0QQ4+Ql5AS6jSWbE/DhomaSctEkfHlCGJXovWdKXC9IBreMasNcbG9EOgfqklZs+
wFtQNhRlIQUwKJAVt1BeFmyLm7A2dplW6KdiwLq9vVeqojgInN28P2L8OzdMM/kDgnRSuYmd4RQH
e7hCYzZEl9iViMn8871iHBbMW5vNlALzBarOz1mMk7+/8WSgFcb1xoPePcBAwz86eoYMqzPmOQUr
3Ro8zSF6LpUA+TM/kNTVvLUExlMqtniL8mr+peyro5CB6uASqiuz5T1qnOqMJEtc6Xfv0w0PXOgG
3Uhv35XsoraFXn3suunOc+ZHA0p7f5I0ncCu7lBDF1sBtLscOwRw+3ZmC49P/5S0Ip7UuepxfI5x
UmlXm0P0Xc35zXLDubdZV9uyGLY/YD4UlzfmIPn/jz4ZKXeIMHj6BgOs3s+/c4/aVQh3/+3FdhkN
Ai7JhJxbD3yl/z3hu7ivnhmoThqGy28QByzaOA144ys+CTTVg3yI7zuYuO2hmsS5G1d6gt/AdJsC
RnsflORZifIn6uChDbW3J7/GrRvSerI9pfEL1P9nfbkSQN8gAOnPQG+d5aZq3iXlufPlus4F75dt
JV8ydCJaaJBYJ6xg5dI3G1ocB45OBbF/q1ph7IlyDt9+VmwgR4dSnhL9ivMY9ocWzrE4Zq6mjRgd
NfnhzxBXI+ERD4SJrVCbmaehoCXZLNYMqMsrrpGNeb7bXCCZV4FDP6fpmme56NzupUVF1uDPGqyJ
8HVaq/eLu7uhAdkP1mv1Qq62maICc2guzoBuNcyaRLeuv696D3OYm/SbAz0miNu6yYZhpsh2cFk2
2osoheOpz278X6OOgGr/mdLHLdhTgLpPQC6RotdXWznyvzVyNFg/57hC30Rm+EqtMGr5LiWviuJx
cos70YU32ONPYfV1oRAwgcb3j44cQaFQaAbfH7y/Kx/GQZH0EHnD8fSTNaJOKJoYqteSwXZuhp8P
CBSkudqVKAV+beKW32Y7bSNahO73HjdZkFQ8HPnivcDtm63L4rZ1qAC6mbHV3Os6RFbvq0AMi6ce
oePdMrXs8/+2yW3cAfAhTK43JnJvag6zOCw3/lqTiLpMt9nygqpN68rYtysRyspmtkuXjC+JJ3t8
C1GBUarGffhcOvsiOUuiqk4asbmvH81OTJPwk+NI2RTpM5bV0h6tLbUJe0U1csgFKVY4uRw9UTnO
17n2NV+0Ms7xjmLwCLzksJPScTK2rTTm3bsl/+IrvctY+R4IFeSJ5V1BzH/zEq3DT+6D2E7szT8t
aaOpYB6IJ2zB5tOp04OACWCshw5wcwBkFWQjV1tim2L5BIwiLIgEmKHhOO45TDNC1z5ay+kQvO/9
PMorDs9ST6USRjeql4ud0O9LiptnS31mJ93jiJhBTpur9K2YbQ2BBe5IxTZ1AbwAMco32NYOg7Mt
xpMPZNChQ9u/+UN4VF2Y5+/Gywn5CP0Z6uj7woNXQWfXaOYlT2N+EFDeKJ3sUpNe9Zib7HjfRe8J
CLK2sqMtaGiqiBuTWp8Z4Jp0Q93OwO8aL2CloD2tSxRara+R2MszymuLSf3yXTXpJ5Xd9IYbIYnQ
TjsyykM2qNyYh7bBTKiZoloXZTFmE6hPlSTjD/+4s+GIKwL1HrVmE05mlJ0dJ0TFyNMWD6GpjfO6
p+OICYjbyahnZrXHJTPbWMa58qlGuFHo6TysJUucTHnoZWa1RLQ3iMdWmx3o+rIFhqEd5lWgSaWP
j3u/bNk/PcTG07/aJm4LZC0/Gh3gXs2snE1otYW+P6aN69pdFQrYUKoJIPDC7naCImjH2AXKZrQ+
AEKbSbZQIHT56m+elfCAVj32bFwLinIMi3TQrS2xkTMCCbdrqqZlRNiYNyQHeKq1RJYoG8N5eUhc
Jtcg7g4IZJTQcdh6VPovr/lXP+5M8J937ZPofWGxymuQxnG7/ugHm085ipYA8lCGaLmoMj06Y8r2
KmneH+0aXTOoDNg9zWNyLalcRi71dH8K8z/RyewdKkxdItOMJN3uKingFiz8TtduZdi8nQhjFAnz
R+4p4PmEst6L4PWeto4la/M/jUrv2Ckb7iCntr3X/kmqg2NikRj1ilyDc/BsIU7XO9hQbdrD3AiU
/Qnv+9QShAOScipSmSTLMhal+w3+N3nQS2QkYNP9s3eD68NfDpmLEFf0eYiYg0UExy42mOm78Mgy
LZP61xb2G7CpG/R8Otds+2vAWRSTTesrvUR/XQinMGKGaV65+Vly0xbASZpyueBY+tx07w3VYL22
m+yrkykOfZx17i+q0ptgE43rJ9p2IgxZT7LFOmcSOHOYKMUG/coblA0kIIQ8cGBkyFA0xN2s2Wxd
HDQ3KQDmQYFdiFZbTTrKtVw6TDxP0RjrB6Lh7CSjMymtB/UFZfXWECycGtab7VtyqWRAmviMe2Ts
aaZ5jmRNMu1EyPabNzVNrMCLhRhR63Ui7xGetei7aKy0tfJBzIf8UUwqTiPhnbn3Go/6QLDvpQDm
QDQMUStaXDtd0DhtJIC7suXTOmxdgg6q69TeT02eyzChDaJm5efcCSKx6yFxtOKEjLnR44RPtHDQ
uynGzfY6TE589O6U3rkYzw7jm5iJkMHUFu3OWZ9MjgB2j+17e05DCuEALcYdCwJARamvCTIKrNYM
P5mJD7bAhlxqECH/R1avV6Wjyqhhzz9UDXXJXL16k4x00MKewub9zvCS2ELa2hdZ9UMoWcK9Dqp6
DBpKrYH1qNlTpcIxnX+bRsUwNKKuhsgxUZqZbrCiqSHN4SizQEPAlIvT54mCORH6LFT44o9eCv4C
+ziOL/SsWntJD0UEuNCDemrQhVkSlOPyGhWVH24r0eA1dwZrHv/Tq/OTLpf4yVfBMDr9A/wcaBV9
7fSqCfMC041ryXNYB1IOJo3P1t9Taq4laJFbZnOSTqQwu38Lv/U/DtXyP+u024n6h6xTarebYDoT
XMQfxslUNBKu/S3qsDObYzuXnuD2pqbqflGAVnxqnRA0XkpxI6HhMdMA76DaDTsqVF/GFh0XgNxh
U7o7Ib86YFex6vKud3+Lu0khntD9UISYYEZ0qm3j/TgFuzVqy1Z8GAAekxgLVXPVpNDV+DrZsYId
BsGlkg0Vr/5ln3jqv2hZy6/tW/ilo/6Kk5BjSDisg8E7IfjH40uiV59Fv19ngESjC1xYSpPO8/j0
raPSVbMl6tAwy9y9BjaYspYHqxtQpBD0X2tARW2bZACrjLm8W3iWzIrUuQxRHi4wX8YeRNIhs5BB
muE/tETq/hI3QBzQLh0UekXbhBMmJhGXKXRJ/1p+cYLw0TyVQVUZUY371NNyPrJo2CY85Wd+ZGk9
uBxWLQyjZsFXfFcpO6fnnm7UHOgsg10I9PWZGZpkw6ldG5Jm5HQJuDf2DoFskyHYTlhToDO+h+I6
lr9dbDq3PAkTL3wdRmLg+UkoyNFfT+7DIzuJBrZuIJh3ZUMU7AHcxpy40BomY+7V9ppVkDUfzDNp
XmXzBXUTT0N5faFShsPyaUwj98NMfbmVjPRzJNk+4tm7HDr8ydF/lKyFUsluzB/lR93aLCs7wtyY
RY+I0WhEm0u/4E0DDfdlX/9mIZNuH/QjRlivWm5LKYqME5MAyYAiwUpEKMJvwHOLr9+fkQGVeGsj
WoMwlLops20SoPpx3KaE6QL+O+qYpTRXEh7T/ZwnUUrXgIWWYzGmtwEl8nO4M2nrmiFD+W+2SeFx
ieBMgPymksv19urzG/20utv0+N1+DeA8RP4DQfmw7GIa4UsWdI7zMYi2HmtoRawr4Z/K23xpdnCz
thwhvu8Jkdg6hlR1Tt+VKX1tXfRuljtlwhqG7LdyZYasp4iDcoxzhTT0nDYgsi1ScnW/y103tGcg
ue7cw48EeJc3qdoCTtCdx41BbQD0/Nr0ul84nd1a8g5Vn8VACBao10ESAQLWRLMvXvZIQFEAl2bi
fTWxQoC8TCKgKXoQGBmt5W6FYMQ8ZBApzGvdXy+rfW5aNYEaRjJSDrDWZzDu2d+rrz7VIcXETDFV
ML3s05uzAnII/VTX29I70l9gpV3KQHhA81kpmKPlBPApEywJMoPhfmdQX1qgPpJh5qIQcV53rVF8
SiJe3/jJjExGBmkLq4tiP1uFdPhBRLWyy0wgsfDF5331jPsspXabrNGuhDEHHknQ+2MtY9kxqEXq
h/RUbuQCEuzfF1G8Hyy0vy2s1bQWzAQix5YatIrEDtRxb9R98ZO6MeVIt3Py3JG0Acc6lrPh3QKp
HYT3JFzpMN+PP9E/s8bBUMxV5R41OnXogNNBDxDV619U2OvmINofUl8wRTdQLsqkNUt80eL8yMN/
2GOjqveCQcjFECJUPR3oFCQv86mixbrOtZmpv1pO/OeYxwrB6ISbC24tNaj0Vz8Gx5+rMa690BdF
270L66pCuqAKBlVdtskOUmuGpKV9fuvYae6VCSi5rf5Bw4/fi1ljyDIRDX8tB1137nAJlSKMZZXb
bzsbgWRBBSIOU+kBB/4ixTZTzpxKojwrb4KzZjbHDdiFJJvYzSDpPIW+hd5Nie+B0Xxu60EkKRfw
dSmePN1DETWbO0jnZCKEM8V8pwAh7geJOM0t3h9Zs9qEqMPdYVjYgMbB6+Tp9lCCEkYjD0aGsUK4
hMR5ZXoAqi5+l1NdYG2hreeEBDO2l45xaDGcvQf96QNoViHlgvVb1oU5i+2wBQfN+D27+wnQPJ5f
dHiuDFRSfQSZK70cPWzYsptWeJmfSfkIQVZAAGynOvMxA2wh9At+n6WpOb0SNp+TN8fbUiGjSDQx
hpSXRi51xzdC0GFdbAj3l4Dvs3AqmVKL1XCg7qYnUTxIK2wRmCLHS1E4YGl1IyomHBNnTF3N2/Jz
UYtNA8sdNU48LrJzjUvU+jNrZxskGBtoaoZUIV8lvanp8TxPUf36LFkCwR41uZfUbmlvMduq9Nxm
qe4nyCk8D+bpJwTHcSQNT3ugcJ1UaDsp51vtwWu7b2/iA5h6M+oDAI073boh1XUbxfdyajm8N9NZ
H3Lvp3gihpk+TK3bRzKbKXdM0iXFkAJ3JhiB3GrDoRlV/ts0seOxUnWFva93Uceb1f591z7CJAcd
0hzehpOZgSSYKMWZqnpNN+bPDAsXOI/jS6zjZysA+W8jHbbVrul2AW9Vmz2SUjsUDR3rR7Axzxt9
cXxqA3zm2l+q5JUiO2UnantMLX62rg8ybYkS0cERNQaru1p4ys2sAGIj8nGI63KCYxdgp99eBtw8
sTo7wfMqhzqh5uoPC9hsJpZ7wVd2RXrbxZ/BpyBWVRr9EBbtniPzbdggPIIPzmGx/8hfMAOOYsNr
PNGTXVLv85dlRbchy4UO8s//AN20G97+g42rDKZ9Am1Pfnp1X4jTqAk93ONGzdd9U++Wx5XiGgy6
gDHcThoRTrFA3OShZIMTUtlLZKOBLZosjwPD8xreZsi5YYpgJkn7FVmkDm/SK2MBeLmJWwF6wdcr
dcoT+2PRxsdKLaMdm38j2fG+Z2iycjShnOsEa9TtY0dNBbqZUm6gRw6jVop+1NrCN00S/UekGq13
KvrNWOf1fx3tVZsxtftfGBNdJQAm3LHMPn55KzVFCxfWnbbnTSgfOVJ0pyRUDgpmfkCZ81vcWV05
tpCfXPiLyfkdRBGYFGnbFB0NJtqyIhRBBtjVfe1I8GzUghG9zyi+TSSldCyeEQ16+hvur3cdlVNU
6H2XFSe9dI9b72pSz+vuL8mQD5tQEgLT0ynV0Ki1/LWUvrqSU0aRM9LM9ndKzp24Z5hyIay9wIsx
LGDpcqLqWy63yzz1IZhH0zHhdsT4j6JKWV56bn2k/2Ane/JT6R6osodPoipagTDSRyBw/9RKVCGt
9IaXRRydR7UgUPZFxdXR3KraO143ebK40E8c1DPqPJ0leYWuLGJWJMfO8p0nOyWk0/gyzN5z2zCp
DSV4vjjMHcNyw42s2I99zQgbTTqYdgIdA/6fPII+WeDPcCJRfrHkzafGnrTWfM/BpsTNy+PZ37vQ
FV703Y4jh/7FBl/Lnn4vx+LvQQ9DuH6diuUm+9wLFF2a7YBSvYb2+jQgCIYiGP6VuxBiblHvUy/x
3R2e/SEcLqDT6+Vyb60LGXwHzBNaViqFl3Trcyabqegkgbu1GfywXfg2SKvFOw+IKdo7eq62F73U
ND7BrCx4DVlPxW2fB4FufSD4ZDFVmMDF20/B9qxBwEOZQmMa+Lq5GAOvYboQmUzeqKWG2JwU2XtQ
9V2wYIEaWwxXldoEd/vbpDGS/0nyRrVTfrQPYMF3KkYMC0tuWzxNQhhDqzO6k1pcSddtYkWRAtej
2WOgwQ/QljsJ1w3W/o+hawkjoJ2Vx59kf1nOxvSxq7Lp4pTHePkDqbJOyvhGDcjE7/qkMBjcKHxo
7qDLYvRuYRdYgFOG+jUUbT+LKezVLe/IZoA3UIG+oVJ8miaf/6q03QCOqV5OuY3y4voOsGEDl4Q6
IXp4AsLZnj33Wlc5xfhzBbEy1HMmtlqqooxgOpi4XbjqQzUI0b0i2q8aEPP9AUSB0gbH77WIz48F
CLXfN+NHvASvJ/6Frh1qUyWuKs7bZNqdHQfWNXov1JHypbZQu9or6gCY2A84VVTWkTo251tpOzmY
JFCxZSN4Ji4Z1xQqmxDxqpa5mPh6Ju7xD2zsNjB+foK8WDD4cGiCdcLQrIqgachyQxnktegOHmEB
+XupeH/opcEw0PMwqKRSCVHCheNwl5E6oKYrqE/tY99P3DyDWLj1qLEj9T/RYid1EtzmUpOcH3qC
rcsrbloAzII6dLWnLm2QJvsTHhfrmg7ITZIz+XTvDcVsK8f8qDgrvhmq6eu8xxAxbG/I9zxuUFmR
dM3idE46SnWc3H1AB2AT/zKsa3lXpTlUkk9DGvPzkHOfbsWlH3GqFNSKf9xw0f4890nR7P4LIbiE
EwkyB76waaIz0lXSxYQBYWPQBRjcXCRreD2jHWWc2M7DZRZEGZkRgLUbHhzUmuew9+z+fV7axvzd
yYIlR4hmG4+e+47Ak1DkJtRofykp3JlOoKwaU909TvLK6y2/vLmPMyGBHTQk0YhSeZc9TGwFhwbv
wIY9cqyJasoL0ag6OFv1B5SUWa4onUd29zcByGeLVKDgBhuSpDhI/ZM/it55pdVUn5EdbdZgMJyd
zs4WYJogJCr+Fe8BmF7eq5VhTfAX621FqIHjOP/1ceAkAuaCdaJiyIUinORsyBxZkpFkPaQdUFd7
qIIVrfAYjUg1/zIuivfpPif+x6qs2l3qiuOZeWooWB6k4KRJGHD6IaKRwwAQCm2KzGkpoTpOcP/H
nI+Z2vZzvkXJM7alEIsbscpIDTnlO8tEjdwLyenpjukMcTd8wgqD0TGkpUB/h5qts9Ov3xurJZqi
/nrWhnNFQ+5NwKI7W0bcIUYHy4uHhTcwuo2t4Y6LhKq1VJF5s/JO/sJYlY+zqANsze5QkhmWGxIt
Dh9ExA4R7ArrappPMu4VRRH8nm36OAeyODfa0J1gTDdRhIrNhayw+pAteWDZ6kEFeJVLKnIvfgZe
rGE/i/RvoDdiS32yN2r30VglIdLsQI4bd8VsKepq5y1E7h+EATBBtTJjHbPAjp1v/occCk0RtNlT
KsI397/N4MkG1jS6btTj6FgNHlKhROtMWmRQphaDnb1T0n0sTZk3uESnBmjnz+3i+Fe8GAQH4A4H
hPmWXdyUjun+iyAreSFslo2+Vq9WnLhhoXFSWBFYRA2E7dypDeLjXQTDHsBHCuDk6jcSE1ts8qUS
QyIRlULQB/e/Cr28EntD/0Lcr29m5+OG5t4DXMTOKtxUUCr4BVZbmn70Ept+Yu66S/LQkFwsvvR+
uPyuaHTNUb/c6NSSuVoymM2lhCgRuGW7zAp2qIwBAy1cnmqSMEll/LiOrDdbMXYbBDcy3YSwjs79
500g0yMmHdSqWQvxaGSqu2hiafOI84g+cNw9kTW8Af59EnF9OsFxRl2MjrRaVaY9m2RamcSfWdTf
qEj1d8ql5Sx7LA8Wn8TSfcu1pNGu23tEjcN8cjnwS9ZBY/6nwm62aqvPN5WSndOUnsMErdIswBcN
88MZp5F6RimxhIokzrYaiW9XET8XZxFPQusgKgh5UtccWzjTUcSBPFcpLt2T7Gnl3snsHPd7W5Hc
q11lOq609dN5K/ltUA1WDBjhH5NlCkmQV5EUJIU74ck2b3gU1NfWnxvxGjagiFS9hRemzkb7LjBs
VaQw/f/o+zXsYTPPZDKwBeRwTPg7821Eh/QT2JigotviqSBtEinzvje+2U2mex37bECOMlOZgC2S
KAf2PHZzspZ+prkB5lGGw79hWJmcNoYVv82ht6FaFVXSguoO6Zf+gjXojvmSq3HAsL/TybSU+FrN
4Gaj9bOzbWAnwndY2hfBsd8gfhiooVTsKX5RHl39nxtZJNkKZUVJ4OGtM5wNVznnBHI82T3QV2gW
tLRUslju0ZdOwHpQ1VStjo7uOYztppPqkBieMh6LBwiU84Dlt2oPPwbOAKrYaKWUvIWLfv/PO0x3
L0jD26aHz5Rkv2uQoioRMDZHsMeoYggSdvycXF7dHWFB+djuwUPcstBvIiKzrv8l3bjQAcMTgwWq
u7r5goTA3WFuNCuYGZkqg1GOgoxu7MaljlVwxaGaSRz3VCTjdMU2sZxo1mNqmYzZNsFgVxpppfnv
K43utRnaERnaqhZe3dC3FIr4d+vd7M7MkGQW/4VFonmjsbuLKPM7feW3PH8UcAP7lOyOvLiVupa8
MJCWf4E0LLYugXgGG7pvp8yJpnxnswehGJAQFpqV20rXcv5B318bn9bN+EC4OXKvJBJjVyVE2z3c
seBS3HGUT0ubSMSF2qvxqdWm95Yw4PJTywetPcoMrMsIisJiIkPR5nUrY6S5ZLBC2lRToTWI6Pe2
vFfPRXsz4cQlVILtK9J0HEOUAlWKu+UI5LF87aKwED9yOibU6wZ1eJO0QvE72qrd3xIGv4hKNF6z
sQJFX2oV1J3+8Z/dZ70RH27agx0zddGDZuJRJff4zJiHr/MDeRuRuDAfQMGPWqEtc4Qx/IeiTC3j
87It7vCq3RlYcXcUo0nSVZIIh8ci49VOn3ZutJ12Ajrv4T9reKdZ3Zzg1XSItzS/EP5rkTwLd/b5
UPrTh8vxM46m35khKd/SuKLG3d7Uj9l/CXSob/kK6CETWkYMlTnymWLMlrHjWyAY/FCcegyvD32K
cGAobgSazdKRctqbazByMfOEp6lfOT107V+kSKuif9mbavD6J5ED/Y43/HS7Mikx3U8v0GFXGvFP
NabA5xNYGfFMn18q8sicxVqeEKxc1AxZ/UTMRGs7qa2G+GWgruTXl9Xf23NXY7w4AOGKjq+wHvV6
MD0XWvT8gW4us5SpVyeh4JEerrQqGF+PERR9GBlI6RdroI3OqKPVBX8E3bS77g+lvFS0kGCurQke
VePvYaMwPbmg9MX6rx2duZ5uvCjOBjpkQJ/6JA+U8i1RBAB7KJIMh7JP4Ycw3JpGnoUYddi6g+Az
7MUwjBynWraatBANabRofPXRBRQY5efl12ts5nlK1Fq3xBV4KgXWjP8TpgIhSR0l7Uci50233yz+
58pCCBhkr7TpxJxuEwDIIhnwT0pybvr3R8PtynsiJvK2JadCtfxHPrLH1eND92XgSTFhKXgloYHp
FSvndWFTXfmuTxbukwKg+EmN2EteFp221RQvYg3Y7Sm0R4R/mhG26+SMOEgzuzK2E9SKpE/P+VPI
Achnc61dPvN+7/OgMAoXBuvwAwTaXDFEv3if5TWnXTr5CtODzLZoK4ErUk1NA7SuJNvK9wWPyomJ
PxymT/ZG/sJfR2IxtDUfG6ndYDsPljffJJnSrieRzZ7dPNZpm8dgmTmvMXqd7un/CKkPCQLd+8ss
MGYP05ijervpIeMkrSdZY4vXKi5xpnZOU7cToCZWteafu3LGRy6kx/A87eD8jTuS8Uo4PhlNsFlw
KDjEBkcBSl1PHrI+PdVm/n1vQCh3m1Ayeg0Hp4mQz8fx4kdc5zYAtM5y/wjxe2PlGqWuRGGBK9n+
pj8UeLxoyWHZw/dOT+nRNZ6b5fvTB/MxcCqBXGJVoWvJzzCHHaNcT3FhlbYHz8Z/VJanYShr5ivL
/7PiZKKC+P1hvDzgbo6dO6EtQc9zc1UilPQInP6IXh0p3/nOcL7/LKsb0xoMAyAYaRxc004TgDbZ
42aNcfOxGAQABQcj9RhaMMcYdKjChdgV3dgin9nsvbtz/9Q02u/bxDrcLnB2x+26wrJZinkT0zi+
hBiy99PQjeo+bIoqbonydt11gjAtOy+909gWlmjKs32YI0gbhuPWZr7T06+64m+1Oo30FGdjwFBF
lk6dLq70OT6Hxg7CySFVa7ugnnAd6juimR5RNi8rAvWHz/Ye5WdX92WI8tk9eK1DiwxL8Cfo3kSr
JMtkHnIHSsoNOZ78nFy84IGnU/QubcORvVRwBQy9/ofRlZWLe2LLSrbIcZPfu1ERdSLiamEElIT/
qT1EjYBMpsMWtdcXCCDvrI/umkPtyNAUxy+R2ML/l/hUTxTFlLt+DfTmNIUnHOs6BBEitjf68Qgn
8UJA3pW8s57ZXT7hRQGMdf0TW52YAS+tJr5OldCp6kuhXcEbiZQkpPysqp3OO88IaqLffVqkt182
a4/XxWf/dN8pPfcghIhqT1aoztcQe+OxK3RzHqDdokL1vb14A17yMfvuJ05+ht4DyVoABCsx6ek1
QICHwHeGrtw84bDtNYKP7H/Qy525+3fsiIapIaVxskHWX1Uk/F9OH0on1J0ERR8TWCZJiC/C0NH4
XlCHT3OZABtm93KUj1hy23pDyK/+YJIgBctcpaRrlSb+IjldfYSv7RJFm6t97/0XflWzbJpdz/CA
LZzRG2Oc2HJs85wM4H24lFCO5XFqG9wWInyfgPMOd0ut9aPhAKBD/lKztA5gVvKwh3uI2XhGm9Fm
p+9CTXZenXzsLyqPQpUW9TvFIq9q4aGVZM2o0VbqEFEvNy4wBzOB2bhqAILSRQn7A0eXJd4shk82
sdFtUO2PF2rkHpQttEjgj342cXRXSicrcs9ZUwFFwSzeIew1QS9OmEwHJTC0xhhmYnQ15zbpGtz4
SF1fqwWjTBElr64Nl9F9Lr/bJVs0F+FyZc4wmAYa0AqnrJnks6NLK1wEOpkZg4U9DA5Xnbjgl1HG
7bPOe+rF4Wy84dkoKTPXHITG01N4x711gp9XZZ+jBg/1k9Evn/FBr6ixRZLW2q87dDfxD1ZfRjXL
7Jsw7UeNrUeruk/I4q+0Nqdf7jsoRJ82Q9IziWtsKCpNjryFeC3eVPji8la3/QOtnrnSNVgQD1NA
qPcLs8mGgRE2UZ75M88fNj2+i/fkT1mBG+KGX0a+rOVQ5QSxLkn/rm+8iBP+xV788mMURsGd8oIQ
CO4rHIBH8+mUzoFnzJNMiZ3G6afIEomd4d1NMocp0Yex0ARbXRNAHMJSKbYg0RB2fA8qhHqfmf1i
IqEDbS+Jkw8FYWmC1qEQI6MTVyBocrvNB4EQHW6vUtQuUxWBtYb62MTEBpWz6vHFfEC83X6laAAY
RVBzEtqqCn9wfUeI9W1c1Hv45brd9AuiwiPj4+PaPSOynDgYnRxWxsrbLngXmQdFe+Csg4GdV4i0
wJGv4ivk+gnMaWCdJyWWlIOc5oRqK7sTSZTG4zKaUR6/KoqOStF2XZWHixnP80AyvS7sBufh/PUU
Pp3CqAllVRr/9iuRcRL1Q4s3FW3lYtcfspJuk7ChC+O97ogPNZxCYtxVmQkgjWPvEzF9TeZHHtT9
PWh7/asQI22+Pl+bjdD4NQ592v9nwTPjLuRzD6BmaGhcC1D4T8gX2dWrPDjfbyMSOyYjkp4QEEgg
ywAGI0YptCzcHiukemYmLPNaQjmFa61RaynJ3SQctBH246fb0YwJ3SvtMDK9MQ15eCxfD/XfZaPm
sue79XZWuPwZJA8fS5NsgoMs04/Q5oZ3ym73nogSJU+Ojy1HGB17BtVnlVNiP8lh5Uh9u0verevt
q+V1It47UyNFpzEQh5eOTu48UgGqTxOFBC8CXo9HXWXiVlE2dVxSfS7ckaZS7ysns1Ll+nUqaZqI
3DSc1IFVs1OhcK8k8SrzkWIOIK9uXeh4NMYOubTX3J6JkZhu15v99JVTNXaiz9Zet9qhrPYRm7IB
nDEX3b1pNc7eQWjNHs8PKfbTZsGWyE4CEO77lREn4vnofiOx64PFMAxwkuWlurvYVkFf0T5mcyUS
EXroqsrDSNljdB8+wi0nhlBGNVFjIEh2iBzwA1MAqdlhYF8Ckot4AnGWxDFMqf3DNlyHfbEKPoDV
jXJA5f+t8ytaUJoRmL+HkT2jlsK4QXxU4h1YJcoL30z4btBTJyVvDCF2QjxtyG57nzy5/YG1ibG+
0gYWfrCTDJMoJJX8MtxFCuLfqhvGgBoXfUcAovHYuHbcevdu2c8PCPIT44Gpy+bWwfqeXloq2IA2
OsQJmTqRA8ud5+Lpz/0DpPnZI+UVojeBAYFChMlqz1gTAdiL76ERl7F2J/lhlZNeZWkJ2seEvikX
+qLFUxkCvgfRyyiKpb++5E92gnUe3CIoy71TcHG5H6LDN4hhQyLpDpe2/+MLLJEfpWRneXEau66u
DtAJhL347Dd/tEMY9ao2bI12YD9bzh0StNUwmy6H8MyXn+a1GO4X2P+m2QZY5PjMEjf5ALimxsIq
sXUaI4LzbcH6sBRcDI7T8Bo9VEhJlWTXChlYxVVRL9HizIOMn2CBGTIm5rwcyrQomlAlVtJGaaFU
gVs8s7szuNYCDT+tn9A97hSvW7HEwH/oG7io2MNIcJy7/frUr4QPQGs0FV807cNhmFBZOe7c8fOU
VQwmw5NBRGp/cenF4nZkfymmwTtnL4763teDFmmGMLrEW3QauUoEJxgr4MhV0u+1TBPHsRvYuHEt
GLNOipRzI2gTDEYEYe809y/ygl2HhfeSyv1pqQtbJc/t6g0Oo5bnNjEMRlE3Zv9Qc09n4RLIHNRm
EHxieASxV34z32K2LoLTulRJfBsRzEIZW1KRuFmfLYKlUNEqnn+djYqnkMnvEwy/rdWg5cWqevb/
GyS4UgrE/FRc6BT0xGNtByigZln74++0zHEfYk1G3JggD9dNzVocZ8CAGPUlyl6KzEHB2Gnrc2fc
VKQDWTCd9ShSReFipL+dTPtnNLsR2+PnZDqakIJTnduRm8Owbkf9mUe9/n/NaNyp0d1f24lrE/zN
urFy/+SoQrQ45k0s7VEeQOxtv11YGuWGSsut2pwi4UA/muy018rbeFzwfpTXoSVAzS04+1sp5YT0
TBhD0rfBS391TJHSKFcGRmZp/q9cHS01mcu603Z24eRQvSmzW80CL2lFWhRKXXFZAp5qgno3cGCJ
OWa7Nnhi/pFF8sEYqFdFDY1gb8AqmxL+gPyiV3Tc9Tejm2hppGw1HMjSGTAR3P/sF9wT4A8iGc2g
SPCocPf4pPM7tuiKpZSxzVwSFPuB1aEd1tUNJOuGJHDhVe3++zF4GE+ekm70c9KFY9pjsvMYE5Jy
JFvctY/Z3q0reDQM41x4haWQwiJDaWy4LokGQgkc0cjqL9gNqzIif0SV64kximOtIbGM3LVT15VD
0WJqbMwUaDA1CqBHAhoWz/KRaIMMP5Z50/uH5lbCl8/AEti/mkBAnjDXpR12Zo1Yno29L/PSZg1H
umtl259QQE4BqFyIL+SMYXGQorjwspTERjUzrv1EJtLFiLB4YKXPVQeadfObRajPhkkWS/0YWpP9
6yvdh4kaGtrrEgZaBaoLoGZScYDpstU/wEQM4m2eTwdfrvFGbO5kc3K+6VEktjFwUO/MZgXpj2aW
s72ldb9pUz94b42jh8Exq4Ax+tTT1WqwnlfRjwZhAfK88Dx2swJUP2PYG90XcRtK9QWdKVubq+cH
uVhTQGywblb1Y2j94f5e0MtqpfaRloXBYIqKZFqIuVQdIe/If9E+HDY2pOnZGsJKprwiBYTdrWTG
dTfd14fGPYfLOCevYgjrGJcB2TNT3KSe3nJOUJrj4U3JLLiJ+4aTGVSSCweFA3RGruyLT2bFWVaI
6y7Bch6oe1M3K2v43nfvcAr792cZn2onFA8CkWdoogsIDjF3YzVasMezoeA3FBwKgycRyqOJpqX1
XCjlYUyfsyhkFpLtuORxtvjbhCt37rzdZbWpFPkgQcX6vyi7VlWVIVSXu0DdYYBJEcRdwFnj1aEq
aRIHEvbBpJ2j9LDSN4qBx7PdTE6bw0vBZI7w+0r0m1pQ5oEjQP1GBc0fmOofJNWCqoTZGoOmm6j7
+18udRW1XSKtH5s2CV/4GVVnEUx7hIhY0FI7M/qqVRXjyIVA8NKjpTuqspUZSqf7QrfmC6X0qwA5
vjludQVDXWvdeqL/E4vtdfE21IVHsYZ9qOmZ3ve+MzlDGbs0pOIM9LqKKAnFQtO9HMJUoWlnPX5U
IgLWff08iE7FuMuE9BEOQfI85F/BpGwSZ0EgL8agsGid/Uzc4sNrCECccUtorbGAx6DkAiqSsIRy
nJg4kBORe3DJm86nggYBSAN2WHi4nmjnnZTImKGzFGkz/KWtiOR1O91FLi2bbWfVh5GTcLNYLEYU
N344NzWKS8ZbOC/BW8xy3vgZQVxpxY1n2FEXXB/9h/l+Uc1wBgDY74emnF/L9ZzquJDzunxxEiZK
1w4Cqn9I8jqRm3jOx2yUFoytQerMtMQVJ1U+fCBmaGqK5ZfDGqFRUsEzA0CD6yinrwYwdIpntNqL
3qR2EN+Mqr+lUsIW+xelAuViILBdfncTXszIXl5x2FCmXXPe5OukODRohNJkCGd20yMSSElYpwk4
5F+/849DtlJ6TnHItcPrj9ZfkOaCCI0mro0a6c/K4siwJhnrhX54WsRf8fibHc8BfuJzbWDxbiXh
5Y/kvGj//TvvgrxDoxATB7wd/E/wXcLqbycUK/ddmKmANYfIqErLQY3FTnPoGBkiORGCVtY8kCop
cAcn11iCW8qhWkKfQUBN1W6HA+nj464fVagGuc31qBzHl9JrhqSbX+DBiJiPwm6lVnB4oiRkDYNh
kbPFBVzJBFqOKYQDRXddGHJk+n/FCPfr7dUwS5a+Ny+PeneLZ5admGGFQBOJgfizA+P2340aHn3N
QDFPpbgdomwgZVZEmikXSuYlnccY9fQo0N0c3PpCKnGvuAcA3gAdTIBw4FNJSiR6LNQ4QibfFvn8
vh8pcLw8QzW5aqxyFWrkRZV8wV0CH/ck91eNAeAxeFh8eFDvnIZrnExgbev55y6/w4StNqP0Q4/K
74P8cbrv+NjrdXSYLiTp0a/OLZHNX5EL3IF3/wYH6nIetjvDcrcUp5nJs+Nt+NlLeuuwuykHF/Q5
MK+P4iskgxhEXjcMr3XTQue4JFIpsKlIWA3Xw/KfYYh4RKqaRge+srbuMk6R+WLu7em9LUglbWL0
lOS9BNxYrZVeT3dozZ5TQdAEA7ZKombvD5trJod22m+R6zZHewP/RkK6AnBWpaUlKVXOLQDVmY3t
6HsWaeMKMaopKR5tPjJJjWTcwDn2uczSaQ+TZJrnPxBUnSy9yPrnPe/HWMjQMHu9aHVqHmFZ4R3X
LMOUz3fpLD7h4Ot7228YXt18lodEtkLShqRcM1RrUNQNXONQpB/sJy+iyOSHkD4nUbl9hSxxr4nK
M0IIrTYPL9dJ6HPdgruF0AvmiB5YjlYalYP16eSx2rURSGMsgvqSa0vRyFVpeOnEvto7oftKt0bS
cmX+2E/yMB3yya1ArybV/OtGWl3XB9efUr5E5vaIB+r28xiayjBYy6vm2zr+fEYQgknTigYG5m5B
9xXpggB3/giseKuwyVaYutkmmD0edSrJp+qmFpZyavcJ1nAfDcV7eSDXWdr6rjj8KfwmCaijDQ69
vbUnI3LhrSK/4qyCN1E8Hvl/QgEefu6OrXeXxnoYDZRzOk63Adc87G//QfEe0uu6N5kaiofYYKOz
JxJ217VYSQgvnJpQY37VRRolLeZ5sYrvaj5HvfJ75GaVeeSY5IevpTA6DNtYAoJCsOdi5BWEd3Vt
K4b55GI7vSBHyboU4Vq2kE04sE+fYVOxt0JlBb3lSt450nMG/ok+T++mvM7D6oqbCDaqa8aklCcQ
JxOMDcK8uWlvpb2sGsBto/95DJ5HwretSb/0isUF38qrueiepjS6jy/7mY7aM38PyLgObzTJApTA
ezrZ8J0S7GDBk9yuL3E1E8+OlxHQoLGFZwBpGykQSzMMyJLdGVr+w8cu77ZIEv1TjB6E/prSuHEh
iwuwNpC8sFJRaxZe8c9MuEga4t+FG/3ymG3b0zpy0MkHKZbPyQxWVemVkta4NEU8fpIIM6q+FZel
1tfRnBAaG5cX5XvzXBszTSc6D6Nlp42ULJRRHC6/NijlGiC9dcaPGQ/nNwEkj6B3qriDuv0VAvmI
n9grDxAnBQbnDsut9JQV0n6Qo3VxJgLQvhjUZlfwDR1sFnZ7HxokJp85QSprvMd+pEdgTVvROTIO
epi3HegcuO8bn8b8okq/ayNgsZ/3gFe5VsMTClniInATOW992HhDH2k/XMlOcCV3KLowG5gyqxdc
vNt29sq7le5snK/zCATgKpfv9pPM3WdNbqxZPcdQJAYzL0iJvFnqv4sUJb4uOfZE8xgeakjj51tU
hOXVtAECDnO9zkww/DDnE60POWLF6lKfS6fw5oCDGs0lYTWrAyMaoXzIn5aJWHteqK1b9X1Nylkm
wTA25SUnO4btQPCHcTUn0AfH6EkffEyeX90CA762jbLhwIdz+7lrSIQf5ACo0EnNXPvApA6T1ir0
ZFSQwkYRE7vG5/v6pXdXpylxy3a6o+SDfCfNrXTzDLqF5Hi8Xl68i5qnrdMsHWqsbnXVDfpH32BT
u4wzHjxcnzeUsTRGCJ1qSkqa/6Eqvzns47mKhVanmpTRgbA0JSD1Tnu6rBqvIApJZC++2cVYge/i
cTq+CQ1MmLBbVhe74rMEo7XooHXV/+t7gvwmzUNadyHUsn58+Wn9J3fGOHyCTezdnWnQ/UU7Fnu/
EKtfJjB6/RPJVApHtCH/6BZxTQFEUNDawD6mhZTxMyaC7GSJAHaSNr7WpwOOOU6goSFEk+IujeHl
MIXKMSbU4/FJw9uLZCltYCO8SOjbLmg5wP7bzmaoYMtvUdujvbHjqzGWVz6oPD60advrixE4kdYb
ZxHkWyqxnvmGwkAcrEFLpAoiQAvRYGK4fLiGN4QcH0ZvoDPHkOXWp1MyZHGBUTOtYD7gW5HZpZVU
o+No5eSK1pY7emd7g6Sgo+OVCB7kKkDGsIWQzLepTHkaxo2Hqd4jFYZfmkVAhXzmbuqACLqgNQgG
97uDtHFB/F2w41D4lGFTXwehvgb8MOfg8WHQFN+zRt3pWDtHXZ7GXnUCirC08+npI0ozP+XNensX
1wOOelNA1vAt8IOjGn89Z13xWQNoWWMfWTNnYQpJGSx2R02tSHIhOtn44idICw7FG34upGzygw0K
ywvMYNDNlwRgq8IrW6TH4wTPisJB+hdTrAylpSfFq2imXwV7dEIZvVZwHn7POYLV8PwaNccPy/Lh
1eTu0jTjgt5472zyFH8EERlEhBDHUGIxIo10KVG8rvvAtiV3ffreoYUQh4jH1eU9UyoEJlkb4o/Y
H52wc1yW94iZQTgEMgjfoH938KHIMxN8FVkrYthju/8WLeCo5MXckndK3aAAeRgE0z1oy4oEJceJ
zxqANCEGsHE0dj3r3gPo72F0HvIRmJhZQoP/nfmIZPnr9Kn76bHba1wgvF9Vj2Gxa+nzpApvhqbi
Ct5Zjob3qaTuRa9jQy/Q8DWrGydgQZ44tDuTtEZO6tDBiwmp0w9UQT2yFwJhxNfuiSQhonjn5Tbf
8tN9i8Al2vsVWI3OTDQjQRFACKiodyFT8JwZKwvCEFNhdjHbOWpNSHy2EKFvJOElvulZj9SPAoRD
T7+f5wMgDmWxubNZbesaEXt8IuutnA5wnmc5JlIh+28iFWFIfD834zElckgvPWhsHOKY5Xifwm3X
W4U2W6BDodQ/ZTiT4tb+V8tfcy/GG6NQVFQw465fM0bdKMv2dgpjpnGJXhfOnjyLQLgfOt4tbx8R
1eXcXpjsouAcjJL5+fNa+DjTGYdfqzbdIHMIHqHZLfDPZlRD58OWXWEmRzdIg15BcS8tJVMidvqQ
yQAJfqHRHlXWHnuLWOfFpTJg+CZiBskYo7wLSJx3fE3aJZGARm646AEXEYXmF5ABRFLBJgAsiid8
Q1bkRkhsMFatACO5O2eVgBp/5Ow5tTV+q5fUp/ySScXB2gneZmr17Pe5hdzMIy7a2UDIZJlBZtdr
2y3fScVGEsx0JZOkCU/yPA4SmHOAVbrFY8AOPNBc/IakvkPta/WrXm4h9S0JXzwTFb0I/eCPgbTB
bYXIUpKWR9p/2QGVAQOop/+LW4SzP9yZeWPAuGGD4r3lb1mLxZ19HvNo+eKv/CPWnZQ7z1xemFV/
pnCIHvDr3MiOz4JQH3IlwYkPOTi3QL7XolbzpF1oCYGNyZAD+zMTEJHRi6Xjl4/he4RQlPAti46Q
0SBoaiNcdi300ju17LGoyJgUtEAMU31ZHFV2hcgrQyCSo/1i6ggVYVnrbIv14s5pJsSEwitrq81z
zuf17mDgM9V1sCwmf/KS43ydkoDWzWj6HNayFMY9HzCPetzIkIj9CAcy18brJt05Sl5hvSJa8LGq
HJYfTXU9XMHfYJ21yPPpkRpoUNwbZ8Fpien26a0VxvgX3zTeFoUWtjjzNXC1u4VrigPBbvhePzrz
hzh0Gyzb+1tvxlQY1eBQeqgT/t+3ZT3NQpHgVrALELcV93LigjC8BEUYXsB9PIy6cc8Pun0qDPx/
wziENbr3M5hCYLXX0CMeXEqwRZ0gI2Eqb8Xbg4tx1fk66Tkwzhc5kpVtdifyfO61hgZrLQNLsS3P
dYxBCF4ixsKsObPV/nDcAXqa130lQY7CSxbe/5+Z3QMa3AS07wwZG3L1CFuxsoVmfG7nwYEwyCxn
0DIO4kLmrh11KmINqffUSXyAzmmXguGuIS9l/5VYitWC3buvk821ImjhMGZ2DGtiIZfK+V4K0cwM
QHdL1TeTls7LwRob/D4ySQbi95iHnmhxD0vZ15UXr4cODmQPNMCioBld+6RQPakIQ8Z/YT7SWMYM
q2+rMoV0MU6Pz1mGuwh+RlAaQDMxwGRoWkG3g8MQ4Bb7nUZPXw7I4SYI7tFsRd/5WDorcF07QOPd
P0sIO/LLTOfWjUJqNmOKoMvMh3MTofp3QWywLnH3rNjy/i71UVwHY/p7U0ZbAaeXbZFFhPi2+/H7
QWb5m7IyEcUBGbzTrye6D1XYFIZznid/zYTlKIQlHR5ljvnevWYhOG++3DcTtDxVXK6syj7EqCRT
enqA2VOtMPNKxqe99WRx1Pr9yfgzeJpTTyygP2Lx5WVDrEBV6gTkNUZzaMOzKE70oQhW9cFGb8t0
xyaRIVFU9jYnk+s7/arnE7X+mjUsqE8yIxYTi43cHcGRJeKl813Q7dn/rhBgqJcmN/qZh0oNRN8t
dcw5kGXOGHiv85q+aZw3S73TNCofw0TZx/pWkWC7EiE/78IvhzR8hITr5nweIWfl7e1+usGPC4P/
1kCA8ADwP9VI+9hQl1eMJNTQbuMUQ8Z8Fm5tYI+UvTjnmAxFYfxkEvDezwWfMOcZngl6HblTUfg0
SE/EPCuSQiU3Bx01fmZ1+fxFdM23+OETe2Wjte6lfFCPb0ZFcJRb9PXgW1b5Y9HLRoJODMj6dT51
t5NRi8pdsdpC47mSJyY5zquIaaBE6xtb9DIvQjdyl3GU1CNb0uCoChmsCldolIz1WY+ePJAZpbGq
UfPPMOD2Sc4jH+Ko/pJtA//+VfGxbzvqytZ/N99DUIOFsdp9W7Bm66OYUYtnQ/9rZqm1we59X8vf
/7owaWE8oKHmLzXlZZXplR7X9+Gp/QrBSUso9OpXBOyWkeDYuzUzTHkcf3HUNimQqr8BwIVNL7lE
Yh4KEjL8KI9+dsZrEkqzhn1kqfI+YGBPoWJEdVdA9QeLWQW+BtPV+Giq0TtACTdx/fODHqMWdNF6
rjK25OB1Dkx47b8LVu33DuqoxpC1tXfwxmzjxDpVKY3/YYk0JWfNCR0v1AUr9Qo8u4emsq5tuBp9
Q6+Zzu2UB13lZuhzrN+o6sVKm3zOIs83KjCz+zMXGlh5Mh7nzAtRx2IfX80B1i5WaG+TCBriaJyu
PfxLRq62lh8dgbH0SuOgZYO2VOCz2Vjdp18+sF+ZaDeRlt2Lvc/hdQJGUpzN73i8My4+MBJMU3GT
2VKyB/cZp/TvNfkpuOFNuVEGHCJfjw4KvETeMqzPqHyF0re5DtY5YlKdFlN93lt5DoDzvJV9ImNo
NmIi48HvrxfbrlYH3S+eOjFcnbu2UM3yGc9xCh1kLWvLb30yUuywGM/cMmmaw4+BIZkG3fbFI9lp
pjMRhKEmoWyf3YOqanMO+nH3lroQsHTqb5+l6nf0Ylhn+d0CTQaKv6rRCCs9F8f8TUgn3gUmLgo8
t2qN/fLzy8xw9swD/kt3n8Wj5I/yNSPdrxXqxg7PFy5l+rwjH5u/CUvpnUOwFTtnirDIYNRbIrSL
v+bRXbYzkoJbcBG+pA63qTqQ4NCeyQ0234pAXbBx8qfrB0pPlf74cqtf+i5iyTwbLcSDcywp27bk
eHbLKpb9D/LJumh0b0IVbEiuvuSFZpyMQdBTE2RI4HXkBXy3p7dzMnBK7RNVG4ZiYC9bgyHD6vz8
qcUsonv3qSK1ofVANsPIoCvK7F4lAAlmliuzRpCLjIhH7dKf/WRVd/cqrE3A7UnuKQfisPNYHYZJ
t50BvVKYrgUBW/DQHOb+s8P0f+zSY8/XOj70ng8EntPFgbfSGYIsXei/xGMLZgTceaR+vTJyJrqO
872EgzMtYtxlI+77JghzSI+zsBAtcw8Xr3ctjvWI8gHB0ggmdB1fzVtfSUK+adp+QbEme0owyuJZ
T5SxyB2uLP5MOFa4c2mMBm6mDMk4+3ZDWrNqv0DWgq7lVZLWL0JQpL7cnTdRcgKW/7xWPsgiXODe
5fuQDSmng9TcezUhbdchgj5ZhPHt9m6HoY0FNQy3dOogYyAbL3rKF+ZOQNeXcRINmFtTlGNLnDvk
pVlMKvx9wQcNW/dnU4jm2U3LCQ/v2uraS+yVryyenRO//lDqdJYcWtjzfapK2Y7L2Z9W7wrmej5n
iFVmbhnl4vWY32ADAxsgJ4r/gbKCXfk3Nb7Guq9Dz3cVP2BvawQJ3K/oTBpsZ3U5E0KZ/g9YPaDu
br4OH3PlQaNm1RAUdSknz6WHihTciA4N1q5HEbJAVfVxqWeLaDyVqtB11rye3uO4O/fMyYeesj3j
f9yNJoTtqVdtL3CdJglLKEa5yqOQIa/cFb2jmG1v96wQv8DLh3NRx3FQflpuGPcbcYhg3NSXcD0o
bcmDrusfHsX/Nwjq3gylPzDmXNBstjYczSzVkFtj+maSt0YOIXxLRZ0J0kZy+JPww8sJll7X40G3
YIDTVn1h80avBzGlVHZkPYccjOnxt/o6xhZrSmHfOyJDL4l/WzE0sgp/Vz/mRdJzD1Nz8l2PPyk+
WCOYyIvl9SQkAC1VDsmyX2eIkJk1s6ouJhbMAtEUVnHzckUemMaIMqwKLIvz9TdmY11m5P77KAJb
higPk97r0j1tOdXxifHr+ra9+GpyZtOhr/WkMsuXFfa+e3K28rJWRC1pd6RgxTU27E1hqM+++GxU
0M2XF7Rf88u/C9JfRuktPdxTL9+0//X833rxoFKXmIWZ/zy2Et2ACyg/Z8ShfKmr7WZ1dZFkF72n
mBFneYKi6SNactETCKzXTNHQoyBGnWKmMblktyX+FpPKUI1j5w/VMlAbD0Wnrhiggi+T2JYJlokS
MF8A/daNgO5Rli/opRf8dEOXL/S18v4ok0F2fWBGTjpeWaXoHo6PbSi6UR4WCBmZSUnWpag4RX0i
446EOisaEhdIgKA0JAlQlSiGr7SpCwMgHS/9LQIUIsrF92/mxtlUgWv9oEhsdQ9meSsyGAMpuiGV
H06je862TxEUavRHuPxqW72uNfRxGErPCnKwRXAW6fuDIruimobkNhxAbjIp7m2xWA9T1VvfRNAz
UYHCP+i22Jp9lpWQ9ZV7M2Y0QAmURoHH4A4FRhxzAWlO5pw9E33+3k8ZTWNw/wfGIj8uy3AOaNq8
9nXBMagY3RvTrCLXZsz32dowZQSJvnQByLl0MUFtzLbDSrC2NglPJGhySAJxCL/Rk3W95+tmrzQ8
k3vwSDTpAqW0p0iAaU/OsaMnGxBgigy0PmPyrfx6f40bvlBwslAd1I4lnPqIu/lwIJvWpKuzcZJY
MfjBiaIxIy7qkdiCwXbOS5RoskIX/tTEWDG5Fwy3FYZYaKvbKlV72beEAUoxS87b26FMr5DMDItp
seTZsO6dX4cE4FvhgFneVhMT2rmdKGmHjuv+UrCqiuwVpy7HK+TJI36Vq+nl54+PQghDzOJNDABF
wbANqhoVaCLRXznvTxD/SsSN6NFWf4z67MF6htj4Vs54OLeZi1DDZbEvdPa6hPMa9vdVwz86oLH3
vZxMJv2vu/rjs0hD1ta1N+BPpQGuRryUJyVd6lBiC7+Kbcm0sRzzymqbkWt+zxFNbhQ33kUYKCmI
GhmTMM+wZEGy02oYpHUan/yX7++k6Je2wkoMwMplsT9rarhp8W4sueg4H0g/cIGWw6Vl/F7dDoQb
TwWPRs3eLpbiylNwB8Kg2fUWgxa4toz8L4sjiqW6/vC+7x6J02x/K3jaALtqeUfxO+l1WilfS2fH
URPZRtoW1BJDdarxNbQ7gHrg8vsoTyQZiaL/oZgBYVRbi0d22+7RmsSnLWJQEjGayrT2gjwdKqZV
0oraV35buFG9EhdARWEKpag/8lYJUuvPA0EVxBUw9//0e8BoE+z5rXXjt9NRWYlL6NYLF7ICsGVN
shCuDp91eqtAhrX/48MHKhykn49JOLIl1fNvYjZKP0jK+gxFQYLSA7y5TdfTyxD3g5XIkkPQbpjF
+T9zira6T49dZwoJlgdWh4inXd/TuLx0WRD+Ljgs9pd6jogGQYhHc3gYN0JCGOAFW78hBs4cQwn+
/PcV1UAUeO+zDUXNUpWIAz0cmnH38DYy8nlA8m1m/vzwcFmNukEy19OeVca35qQS8lAVcNtz0sym
+P5rEqvb7aYPKDCYRyFKdqYJb4O/shoEkq2fxjfPhUCwpx8Jr57Yao9EGfV50BVTS2zYz5WdxD8f
/BY86sFyRTyd3TFkdniksswHMxKyRLAu4Mc8wwKW7021MZ6c82GW/63lztqJSV3hiKKzJ0/Wom9/
xZIDGcnNWrvtkg4UcSsJNinL87o+7XyGN+oezqndGkimHm9dC2GiYy1cVFBoJdDIWojXjtQe/7lo
X7kjgoYtHyfd3x8ztXgx9UuI/vP6ILK0GfEtwjHL6U2oka1wpeyxEC15KpJTKYeBOC+rrgYlQoNr
Y9St9Bz0EKD7zlkbxCN22LKfVtXFl/Xne+lGnHPnD1tyevmCVBspNJsTXYL+e9WixQ9i1KNXuj82
hCA9WylDcSIr3+69Te2Tit+NjngBucchmDjlY6ExNxZDiG03194i1IBtQYlWigogegFI67CV/UgA
jtjmwqJr2wBHE4L9TgwF6GPM3+aihjS/jIFxzeEa5E2wCTOZzC9+joYsJO0qZzogymXUiOxN2zgK
iVHzBVMbi33p/1Yr0Kj9gTH6p0WqUS+WcXglYAU7Y4QnA26S+e3XtMaV0c7AkI9baDo1w1J+ijow
fbfr12C0BwABetpmgvVP1qJAB41vSxHrWA6uTGSefGnUKSiUvU3pirVtHfMU5Fu1O/lwndiyW0BE
YCSexWPs0Z5Cdcniq6MW6DmI5+bNPKvLUbusNXv3D6HE8Qt69n0eBL8X730G0HkN6WeDxmfcXXkN
h4LDgnBecbzBMrj9urO9V8lyS8ptzHzPGSiMMdsp3dBoYEW3I/CtTSDNsvXu6ySIl/OO3RTsPLGe
OpWlLLMuNyv9cUDVd6rgEk4ut4BSZBqEeCuE8re4n3CCubq/HCn6MBxgSLfniIQzXEh6zzOgVwih
W0q4hCLYRKCPoziwMnjUomwELecCjPGB33sTx4iYBU1yPOIYcx3LXkb0gR8DV3YusYU3cBMWrniG
jy+MzNKgOCl9N94rQBTh3RK7XayJiAZWdmFBg3LQu2gCfa2UbmdgSniqGd+Z1k72haRDcYDFmygo
EM7KAwzObB2qeTQc0setP0t1GX9FL1DA1TEACyniiUpogYzrkR1FSxvE4XqfOwxUBQfAMceSquiE
Y/i9wTj6zOetoocGmZ8D62M3FC+AE1Ul+u6jxBaseK2VGKwTwHr69b90h2pgLDQsHbIgHkNvEDn0
VankGJlghrqwFH/94ZmoxU1As7y53VlVN/Q7qRWoyyCW6FWbyUFFU7UzN3CcfajwAm0iAaIRKfNH
iCma7KNQdJ1ohPvwGCb7QH/x2wt/Ny9KMU6WX1p5/MBRTpXe37nrv6e+ox5rCPmgEu1SbsqlC/m8
ANVaXnoTyjJNJA5Hl+TKp0qdQ16ci5viJagci5cq+jPuNR332D+CCeWh5LqB0RFRuLtjfm2tVZgi
RaeKomHG4blhfvRIauRdCJksyH9bFL60XDYmp5yXuUh3NjiXjlOYw8V+Ob744AWu9x4CsxEhTHYa
BQHeaY1DtlCoDEag2A6WqrmQ/fBxOQArXtnysN162ozOBrZhog6nbT/ecUUYWXUsFTfhBwBCZpWG
c5Kr1zBrY5a+NT9iMNToNegSBdRRsPFT8cvg6hZqdWKTk2IvvY//VypfrbWCf3fpui5yqy5GsStw
W7Fmyn5vW6um2gnsCRs4dYviVAuqAn+7B8CHbvl0ifEV/TtRVcUIuk5UaSE+t7zSmmpJ4mfxjwZx
REDq0uad2tx3QeYeTXeO/Wxiy/0/52husjeDAI6Yqf7T9KcCYvEKBRHQrILI7Rh0acCW9Nauq7Gm
old8nSBhJTlulineo0egzLeauvGBLih7ypBSa+5OqzUPUwVU8nGMhtboBRK7OC29DN4VXcvMMK8c
4t2kktRAczqlmh4favdTraDRLHHf4WjTdnTDNr9BInJxvbDX3grSZzPMl6I1ixqyPQM0KMSQM/mH
iOzksI3cMD9NOrNv+4vH48sswPw5GMu7ZGVhhTiZj2u3VySSlfsZNcFCRSdodhC9ooqaoS4Q04Yw
sXok3b6h9zkLGiQO4MZUSzFteh/InzZ/Ay8OQdLPziURtWsgI33NvHfO2iYGVMy79pGdvGW0Z9U7
d2jqMD8Ia6ORvAY86nihJJ1pIdSeft8wUeRF9HJqDZsflfbsVVUQ3LyzYml4B/MmrLqCTh1W67NE
Vpb7hC7XPVf24Cb7N2orugJ6TZnvIlL6vJeyp2F9cKTU/QYnXjVBFKdPj+jcpyrivyQ8LDUZiqGU
Tova8dkkZZpXaX8IIb6QYfSM6K5XLalZhKwYtX+Ycv7wZcMP6BLM3+GKQ/0Gs1CeKCw2QAAPnA65
8v0aRrQaFNbqGCjnlaCRiBqtort79HZnGngNLzR4mAi7DLZaZYMO4JbOAoBiup+rmT0tfOq5tQMc
ofGmFOeK3Xvo7YERPfhgk+/Pad85oyobw6AYI0KUyCmviKu3YfrfcR5fxGyDub010bo8IcJMGUK6
Ww4zJNEoSPn5ZJDs32Fyfx0GiWaskodTkXnsayhJZRNiIq6a3NlGnnWWE8z2A/P1QkvLZ6fLS++4
Ti6gHsUb+p62lAI6Gh5bhJ7zJaI+NkGXzz7m/Ep2g2XmAL2/X33XroQR7vYjzZxLr0oDc1SAiE1T
IhzUJYhP/M3mDMfsTEo/xdvjuOTuIJlxx41nz0XtjyU+oydXzhqw3fWanWqVNlmRL6ycXqwU3eWY
dG+HP8uYiCzwr1kCQry1Is5OXvdIanfI9rUsi3yat2CXnySX76fhtS3Z/clRH0aLIq00RkonUumX
lG5bxGMZse52Ziy8Pcq3vTgoV/qOawU6hE/ouafJnh1QfEphnji4pMhmyjrs/cSS0/XlC34UZT8g
mBtiPyXhYExq5GdMZsndM9CjJrogTJTQm/2aRDepC/+CEjuLd5M4EuMJj6GVBSGu2pGcdJT3V7tt
U/4ZNZVsVWdWTNtVQTc6YsX14RiGeMWLA3FtASgKKPbuPakrBVQhegRm0/GUTkYceKY+9nU1Kdhz
o2rEmAMZ9qU7Qd+max2ll5GEbbLxojMBKPhRF7Q+pDede5SKo7z8hlc3d5363cwSxJSyj7+8p2hi
spbp/YP0ib6WiXidwqcCHfjck7XmhrHRWx2UyVDyJ7MGRNB3noNR0kh33ceOL2IhHW332bPsjJOz
kzZGhBuyjrA/Xfp2ZIOqweKnTxMlnkcx+3EsIOE6iOqNZ49A6uzVLf7b29DpzXMEL+cE8mykC+4x
O+1t5W7YeMEuThBxxnWwjw498Z6fGSpuJvx5GSxtcKHyDBW+ctu5IvlpfifyvHMex8OTtfW4Ruf3
KI459JvhmoZ3w8XwGUAJwYThpGIAx2m+LowSH7VpbkRXWEDYEuUYl/yZ1ByxIT50WBjRUHLnS7tB
7vXuNBVp2TfI4CaH8mCGPx6qjK+lWBSh4TZ8NZkqclSKGV5b+1fgEKfRIDcL/jAm/ZWkLcaczEeM
UGwxuVcMUNVfxvaBONgbPFeY40MbeS+wzXzicc+aBZNdlHOPR9IXcu1NTTy/5L1PnBIK5T91RZU0
l85fj2I6UzM461gIbFCDnncgvtJeD6rm9phzWh55nel4vcvPA+7mBplKLi2HzB9wWs1IUVp74JET
HtxkcNJCw2zGJ8yZfiwnuKoVourJ5RT7Q0ucj7kOz7q59xpqM/97yh9InfMi1cRbn/FlCyhZSeq2
JenJ7aCOJGV/j/YAVGCm+NEl30HETSswIz0LEeHmr4PxXo486SO1+SC7xu0oxhi+Op3eugkZBBvj
dUOdiYns7v9l+IP4SN6xDEW9bH6ThWggDzV6TJ6IF6ahNMGTtvwNOnEgOuMmg8FGhKt8ofi63yzq
V4RjomoDQVNIyH/MEuPDswkayDDFnVf1YqKj1U6wOJWCALamve++K9wweU0gDKsJgA/QZlBxLGgQ
OES712CHUm89WOShukLQ/uuTMA1alv6yn8Ri64zO9VMoZ00seqL8IBVV5TBSu8VAEzjuOjIq+fWk
INsGo/J79xttz0tBVAVnl7zHwGpraZV0mXtlRl5FqBFDepnSN3P/WFuMoChH7EBGq37dXoATHaU/
oXju30DWS6JxgPahVsWOqSA/WAuiqhFZBi2gxmLinbIROu0kU5x27UZtj82AqYeQtOHds7HBeTsB
qFFWV4kx0CC6NtcgsQINIyqI/UkdJl0ykMedrAbVMFky6BfFlAB+ufvzOsI8DtedPw0WpHH/OFun
+APni16smJY0NVUeIQZPV+h9sp287kP63A5VFJoPpk5D3J1IUEOJmHL8aJj+jv2VdY9mbBBt3/at
l+xAoYaQDFQFKlLOE5gK1JzLBB85AXTo3yBZvZylhaHQf8soBBEMPfL/O5OODdNUy8VWj48lg4nB
Hhp0MxD7P1jCkC4kIZh51CPmhBlUnZcARRm+siyfyOG0MSOcLmvMrABigaoFQoE7lh6egmLisCqJ
0qhNH/I19l5o5Z60nY/Bu0UvYLzXPmAzy7Qjwg803gzs5jkayu/4bcCltmdL2r8emgUAUZh/OcJ9
Iy7fWdgH6GYYskkA5/wUiTYfthSGzmuvM2BXeSdKZQzOsyTi4E5pRgu56HNHga6qvT0v1UDuiVO6
H4pZm+2k9KaURN1fp71KQXKlPdo2ceZ0FC0cJgRZvlm+c24fAi6noF4gP/Q5otAGY+uZMuOmIa8Q
abPMln5w7bCowqB8arUyp9mEREQ0wvA0E5dLtZ2QoP6yBpNl3CZjTgLr22PgqJWRCjCsXjEe6xGB
EEkCxr85aiYgWL/asxEHF3cMGXTx7ZNHBLoKa5nqiO/L/yxrQlTbAEchTCpwoYNQeZnIaSdLkwoN
2j6eTmqeEV3HzRC2UErdJdkqJ7JvtQ86BKr7AIHqu8S3O5t9CrSsJ9rDzKhctqP/WSqCjO1P8Jb9
UnGWOOXdeOR3a+Nmj7E/vgv2g8/IKrv3zb/iBYIIiFWQc6MNI1IWdn7SNNLQkuH+uRsI9PIMaNva
teCn12iVqwVAOEfiSuALwQljO7tZVhqG/SDyEyKPLaL5odvB05xCM2DNgIPxhxDIQldpIm+G6HDp
uT5sBYp57aUfXnxwMgPxT4iCWD82A8fd6wzyoN5r1XA9lxQ2e0TtHWeKvGvykHibho+GjdeWuTGK
IHIfrurHe54YyKokg6Lj/gwrW3F68wdHnxViUrqHS23HMO0P10QcorWOX1t/CqWmMzB3gGQnUjjt
RgEz9lI8f4kODaICssGj5QqcUMaCdbLvtDKIcL6pZwn1smKD+eyqGdiPc3Se4vh8K3/vzxPMYNkV
mSOSGxdOgMnCipLtde7RJMlGSBO6K13xa0TR/WNoOSVaA4qBETvsNpGXP3uoq8tHN4Uwb5BCSIFZ
m6p25hVq5tllAsI5zA87Cnif/+Yz+TeacAI1c4c3hlUJOwo9r1qVJPWi2pH93HHxl6GLVuwZHJ6V
HejxhoJ3Kk7OaSkonVfdAcy6Kby6AlqisudT2N8KKV3geaVn5qvMZr/ejUZS4hDLOtvXK4WkE4ZL
0Y/RtIC0X/dwgUCQJ6iDiNnyd3EUl+OdcWyrvCms7OTDmOHrFtVTZktXEf29vV1iCFQEd5JCcG+l
Ckz/OtddWa2v9r7fJ5JZzsEqCy1O8k10C6D9ZdNORZCvTszUlVKZEjWO6dycw+eEOOcv+fqBWAKI
/uw1ZiHU0pK85RDH2+yCCTDxDvFo09XEdLVekAOyT4EdAVWiuCZazCnEWPRUltdHbuN/D1l4MOc9
vDQOgRrjf8pXcVe3I9MTjTc46l3/wlfDl8kpHyI6KqKmW0WLwQpEuhwT9SFMPgT2PLDzp/G+aqu1
GgRfThliIkkyX7jif3v1z1DajpQayN/ygqFtzVdI/b7B4Jiarwpc9dIr23L79mhh07VvZ39loda3
XXzHdkChnZEDryCYCTUCKXd1QHoimsAjXDtJvidxokNvfKcGZNQpH/pqKJEDrPkKnz2SlL0usNVI
zpA2Gi6Qml2rZT1YTXsqLwAVjWq4RP2Bz/nlDAImNQLOZi/3jcBOVj+KA1U5XAf81cqsrlKRMAve
B3AXGaNUeatYsqlYpLqveszooVFneEr7ibyFJkCP54/XXDtIW0u4Oj8PeQhDwjqhBl7pPZz9JUGw
+b3cyleRB0XSDzGckkCs0fwFlifJfE87i37GDbBRbtJZsL/yzLMgMaH7BFF+LgBN8WoFBQKHbMBN
f3MjddcCgIBA5VaYZNtuUIW34pIv+IRvNr/ssaD0Qcl0ZjI9CGY2YjVsNivwqydjPCTczL1BLFhm
mT1sRHiIbzprI1YU4OIsL3KD/dqo+hKbawfSVXaq4TudUsMvn9t4ALPgGC3kxuFdg5k88hdcVQVJ
kD04KpNBA7cCZuiecOuPyExaZCyuWNoVtth22V2dwbZGySbzbZ+TOzJ6KYHmzM0jiyD4dVOiKeES
BGXyVCw/iqYKctGLeob3gE6U5MhQOYRYe/U3C8rL8IYszC26+1l414/cX/FNAVplqChxPpXU5f1+
JAvguEqvF0HjkOzKL0ddwTIp7W2DEoTl92IJiu+rB6w4fw0dODc3zwB2L2EvkHHaiPc/1AeFhTQX
bMZRkm7EjynEz0K+9HwtfXzGkWuOtOS0R5l2Eld8lWxSIUS+eLC8qDY9KIlK4oyRLo9x0r64ZLBE
07OeGH2ND7e1Ccp01mGFKQdhbKqtGO2hopu5nj0cnq2ktLvvN5C9tSpoiQbfFmVQfxItfAWrsoEt
DwEtu5Oy4IhrwODeg3tmodito+JdWpQMKB9+OR6gffZ3HLPed2ZoGWog6YOP7VSp+C7ev86RgHmj
wN0lxa9g+yVa+NyLRkdZARmYZ1umy24v5JzxKYIxMtCKvEbCmT7Q0WO3OlS2Ezc0/8pf8YiBgdSQ
TIgAyrWXGU0M2tv7rKFUjhdQXkcUH/1zzRUr7rGUoHJv+wJIVwSDTbVng7W9CujpaGIJeQVzqNtO
S3XOMUdDP80QzuoBwgIn1YeaswO7Gv8pKyarey9l751VTMTOsmxxuGmnKXuVTMLLywALp0llf1OM
22Dv844GIdXX76NvQuAHXDDmTVqnRJ+1WHDQSlpdnjbOUJiu/wcvMf/1+/YjLe+VhqCByXGaofmE
oE5vu9oc5poZ+70fUK7rctN2T0p5DSt5nu2QY62FFzHvTOted98Z4y/MVitYQPpTSy8FSBUbicxv
4H1sCGR+Ag5tmpfLbka7DSCOMb9OnWafyw8rGZOwi8B9hpx4YZvuMwsONsT9hws4U3qAZwkr09mT
sjX1rCxQ52wcH9vFH7TyxR9PI8Y7XD2IfyocTRyIPzhq7b/stqPDKf2tEPl2WPTXKoYALO/OxTPm
t9zihQITOXegN/ciwz8k8wriZa7B+BC9zcE56G8SUoUdbJcqj4lGagYuOyW0+SDyOp/Ead4BK9NV
AZzounsh2ou8+zPg8gUljIZKVOI2zgGwETwIojUCTEZf93itHu3laGgxBsgJVSRNN2fkMck7rEBS
Wg3qPP+Q1FZ/Qi8XNaX6EbsVe6mQmVxN0QHWjBg6LacupW91ugOysDoaim07QpokxhcK20yjVpIn
VZLyDJUP6HP5yU7vYz3Z4urZ+yZOVDicZ/IpL5wl2EYLaMYfqUqCuQep3Jif+I0qHnlKmSzcKETN
SZhWf5WuFRdoTm62tbuTBbKNRAqlT7+3EzAn5Qlb8MVR/5Bk0jn4y4qQVdLGrkwmnS2CQNE3Wh2z
N/qDDqv7Vp2/ArW6phaq+rRpHcab0mXqRB6Bm9fgL5dktQ+wprm22QFguU8uha+07g4c5cgu08XJ
xAnqW3ucdLBEkU7Nwz6Ug69+jHcxO6e9k9Nbr1jCNl+34Suilf4l84ZVLUzSlh1qDt+SFhIy3LW1
1i8eoPaMTiQj6xqioCQLU582wKNhk99IV32RMkg1wnYOozJhzzO/f0RNO2EGfIMP68EgYAtVP0TJ
2pSj8+5f8DIFgvcWiBMJTl4skVJX/rhtQnz6e4iAA33p4a6dZgeNUEJzS/gzxAxWL0ySn7ng5VFU
AaLqESwMcCFu9Nk0RLh44b7yZwwFVVW+fSAIhRjseVkOAykmedvyuXjy6DsBIjKjYHpZbAriifey
QzkH5jl72sSe68xgE+uQO3nYA3fvo7SFtQa/3dk6WJyYoKOcXkf8PbphvoeRFIuQCjgwrh2gXAD5
eYwR0c+AL2RsmqoRCEmKH8rRfBXQCrKjOzJsSacWwzR3365pGYZHpIY9WlOFx32rKThJBQ0xDOD/
+i4pPbGosqp3UpKjRZ/0Lhbg67Mh8AnuusoJ0eUa3IBuR1uAjgAHIBRY1Aw7q7wZZ3acKruwpsJa
n1Genps5Cnq/m86p3cKtaV1zmaVjncAVmwSvKl+ZxbZ0SbB1SfOgB1PGohmldzt9YO2PpJGa0ADb
6k1hsdMdGZ9ofgilylJHNdv5UtvOdqfXTvIpfGxH2YIXyzGvC0kWSnJY5+A9eQ9t6z5NvOF5FsO6
6+UFFaHhyxZI4eydcq1oF4cx8jdd5DtbSRlE4tlt7BzwMMj+P/BF2NL2jvho0S+9dbrXskBVA5rs
3gjOVUfaoU2i8ttnpDB7pRGJGncWvdydnQEe5PHHzsjezHIKONjx2b5+NMhyqzimoaZl5S6RSKOx
MyUTrAyr4Tr7idelsGLxyUj1zR59TQWK7l0+p0m3qyhEd4+FfswPVSeICI9DCv3t2YeYINStM1vH
vXFPqI66mO3H9BHHEowpzfjHLM1aWPRf9/ElyMmwDwZzebMUWsQzTTQEdRnmGoekdc90hBYUa4KE
wlimkiVAwDIbqsPBwTw5QucespatcJIHasibTxAplI/XmItO7yLVk5gc0JyrUICHXutgv8/zz3Xy
u+Dl7VFfF/Qw/M9os22YY2uQ5nNCjW5WAS4QNirgeyEFoddmU2FYAhEjJWXwkAtgsXnVTiy738iG
hROpQW1Riqy/UZ4pEW0ZMtiQEvey/BZ4xsLjDZacM+8NI5SVhOkhHtV+C2i0hKUUW/2x+RvXTZ+e
cWUf+5yWi7i8EWcckRdNMvHS7n82MAgkuwO63YYH2jYVx/OFHjWYsIURUCRkCwwE2lT1LHO6GiRs
pjckhqH7Bu9F4bPgCqkDGHj7GP5aZ8eRMK4OW7QLt1FHOdObvbmY9QogjhtW7N28X/pLyJ2PDaAs
ilfpC57qBSEkNrpms4o4nIa2VO8Nk8QC9ajkIjbhaUL/V8k8y/oKx7p3NaIJmFZoReFYrloF9sfT
GJbMNNqUXunT+JdxKDiGam5h6zvMAh8+SVfP3PmeIPjZOhyxAdRBjyFrwgff0H8tOKYHWP7/uoYu
fLwdEmLdHs/C0w2UMYvQmgY+cxjW4lUZax1vpwAUv+zzEF7fzpYh5HgkTq8HS4ND3Amb1NWhXFx1
234nxIYljcl9m0HAzpXQRsWEzEb8B7EB0eEPa5XLhbL4V0m232fkmLZVqiFYcWRjrRpFLgMKMVdu
MTICxbfZr9uKSpGXyP7rvzplT6v5QTvcmZCGHsQYzwnqWvpEx2xhERhaeJZCb+01+j7owy4TUgjR
i1LJZeA84s3/U8RPT0Evj0Uthm8sMd6lkdjobZY7UgdKRQ8Xct9+XT+wbGzph/3vdiQgqGJC2yiE
hy1TVDpN+3AEEFBZE4SrjUKvpZTnIG33lVHd23C8cA+58Fg2toN8VFPK/4DuAi49FYvqCfqOnfsX
/ITk8HW+faPQAeNtmilagg4m7H81npA08TmF78wHOskQeVhwMaiPqzXtHh6MoDnxP/FhX67dFfua
redXY45gpkp2gVe439aLe+LW5D4ao5KTVO7IudmF9gh1DrEKKXMSzhrLGPcVqLKZ+J1jK4Ux8ULQ
68W1Vmn7VE8s9qHMLJw1o1zaNNGWK5sTFg9ip2eYQQZoFiP4YbTMCzfB3bCP1Enw0yVZw+hEWNS1
KPbWiTwOKwUmrPRLiFbmEpvw9B89hi48v2szLs52+X37neqnWtm4TbyeaxgKrwUE4KpeAKiXpAtw
4LhBouhJJ+HST6VDjQXxwXOzQ/fXh7nJa2uyoiAoTQ5dPjf3bVI58cY9ByT4gv61FSEjr9ScjmuK
fxJPAqVvrIum2Pz9XliCLt7JfyglN87tjt2UPS+RsqXgMjQphdmH5HR0LFMR3S3KOflb7zmmfRFH
SocTaM7NT6AawoF0UNBTpt02Q3+dEUlk1oBkyDe1C/RVEDSF+eqKGqeCjokrYmjMWlgabtxNd4Zw
a0cf/qv3+WxRor5ikx8o7v46iZLMRzlEVx18oVVPKfHuaja3QOIr8TYuegEr+B2q8ihSrVSQuf0e
fAYyDgpTeRT7XYOb5SXZzmfPOhmofkcqCSJZH5bmZFZRl9/LahtagjQst7qd8ITvhRyzy9/dMF5g
LPRjaaZIdfCh0atXRpiA0A2jOISwhBUzLCvhDOs0DFCydtISETX16HZP4oLqesoei0rNqnuoXS2s
6G+xFUea+/xGFzTiPZX0lfAoBGXgzD7H5TMQNRWxZy1Vhxyk8Y6Ww1zYl3BlrSz5F21lMJy/NQ4M
mI0J5xyl7VMcVFqGA4RHJ0kuyFAXp6YIdrhjhE53fvNkT0ICsxOKhnYy9MtEdJDrArIeq9b/d+gz
UQNfZozKqZXOslAZ2FPl7d6IEe7tMw9zDVrqPWjmiJ17w5N/UGUptX58rOwJKbweVCCsomVXKdSu
aLiMvam0++fkH3Z8xz32Kl0E5DJf2MRAbiFVHQ7sLfF+Atp6m4uKFN5MfMoMmN1XE8xJisoR0gBs
XFkL2oJiy0e2tsq4gxrglIxjWPypyzGL5CTC5B9Gli+j9f3tO+TBhTudQhiMRdXt3YHf+mVnHiBB
XElBJeWdMXJviqCk6xACjqcoAACBeIkJyh7vTRiRk6zB4UnUgITc462IUtRYQ9Et4iu04/WY3HlR
3ki3T/0lapLuoNd8hwapBsE/RqT5UyE68AgAJRMEmzj3yJ6Ubc04RLpK4XAdwtJdegzI7E/qHMCM
nTUoHKN4Ev7yHMaXi9qUtlxApDnIPleRJv78a3w1U7LGxeRjkjvTXZaldw+P+jb/+fiHEl5Kp73J
EHBRIlqhb8QGEaXX8zHxbq3J2eNzip8KXLwSiUeNIgJRLoHKauzTXzLAQsm46BDkBjeFQk5R7E1X
uq7GFFrtgv/Ji23OuweYHg7MW8JirhzLem0dUO87IXv1F3exBDhCyX4u2gXWR0LaAqcZFGaXMSEw
/aU1fNpKg3l09AIdlqcFGw7xnG/g28T5rLp3541NGkq25LUhHfzdkx0ECVQQ890muhUmd2P3+Yw/
6P/HGp2CtgDrji40aoUQS/DGvtRXW16JTB5BVLfPemrg7HT4wNt8IYEyPpfa2fNShf6W10ViCD+4
7KMjhFZEFyGU1vYVyKRcUpJSYdCDdqdNtVfVH3d/q8+F+Z1a07RrVgfY16fXzE8yB5FBLqsqSdFb
B2f/+U7sWMwnzQ7OJPpv4tPId2nVSDE25HYaqmcRp4oslXIpUabfr7fkVMEV4ocptPcgLbgAKNq7
3ajt5WY3Ou2YRGIMM3dz4NxgGQdVIjKjKJnIISa3fqC0g9xPx+2XtTanWqIzFyCFM3utBcrtiltE
UvyJMaSnH86NtV56qpuEX+JTu9/puh9DXjB/cFsHZPyz3ynhPO7Q9dReDoIhlvek690pH9fwDVo/
zoyhh7Oc/rFwrzZFC/jGBhVdHuwoTelv1dM4txmvvpSOcWkVZe2jImjUg7UzKE39euYyDxZi05+O
WwO1RqUGaPq3TcK2RU4uH7xqxIogx40+kJPaoXk4I0yUV/jMEOrgxaxSQydw3XOk80Kjchnpq53S
qh7fUJdvz3+JKyxh9G4g2yhaPkfGJcGsOXtf+RUqzJbfqRCxekpMflxfK7q6z73i5FiGHdrIhN+Y
sFjDu39lWx+K8qQnBY50IjGsyJChngWotfSpz5IjnMKdBQ/60AxUoggbiGHRVvjWFRtkJN4EM3gg
+mSjiwyAeTxm59rkkv8UNEzyJh3ozs6CCxslii8BWpQ+N44TRdklybQKZ3hSWiLxau8ANdX6iAFF
qKEygS1kAG1IBHAukp9Z6tXWofRdIm/UdsRwEr99ppewlAFmNzkDMyPWTz0iQF4BgrGY++orsMG5
KdpP2GAFk7P2uuoD0hcwMmXBn87Up+ZXeuLOVRpEOUvViDFuaCOlpdBV2mkUKFhqe9L8ZZNQLk+E
MV5G2gGrAHZ5k7Hvajp0w3JIQGjL5e1sHIxbuVN3ZZ1Jx44syv6tD83xX+s2hadNFhlAPkgvsavW
3EPB+JkwEwOUU5vwAUFDwZAKPiA3rnltn4oKnl2HwZJJn0guFUlZDV0JoF/jeS7AwoJzSYbvpW49
B9Mebo08FUgCRS7ssE9TXpX0S7+uhRIbgI8FUQIMKTB9kKzDnzhG0KDnaAoorooGTGwEYkZ1vKUS
dj7K/ghu63GGnDPlKDETg/iHJdED4fgv6avuJ06bcJO6ygspAzCq2RrZAWPQ2obQLqR3oLk6ayA5
A3SxUDep1ShUotWEGySNVdi7dTc4JT1cS//h5Uddb6DaqFSDk9t3uSCQ0jIhLCqdYID7BqHEouJG
w99mu7zIDZYQ3rQrDwBfj1JQJul7AS7MDz0E2rHOFMl9d+vHaSK7y61+XLWKFI3I98nmUNQDh160
nCSlND/W0nDjgtSP0WOU89cWIRgE/c8wG66xgnuNZjAngzwTh55mSqa9rr0PWZItPLsK7WYWDlat
XLb2uHvccx8c41YXauPtkgTLWtLX1FbuvqSYbdi7R/DJdYDt/B5UgsSgLHX24gDhRHzP04GLDl93
5PQqkQY+ZKdmGHZaqRXr2hjyeaoFRpDpw0IXvOH6c5qd/EauGIMMjlsdQoCa76t62/m0Y9SETaFw
X3gmTfDC9ezcWQRAejnPOfmHVPRH1M7NCOJGbxbHvR/9gDXJiWplcj1SMkv5wwvCSkjd4f4CsqdC
VbVkmmTNlkT0i61XMiDtVxOGKFbsrySDLFpIfs6Z8Ar84WEezCNOwJwaigMaLR4H5OKditpylHC1
pXJpP1Set7ayhJFlIdnh+z6GfP1zX15g/cycmx4unf0x79XlviJnWeiJWs63ALCF7HoX74+J2rS5
noNKUaYngu9vziFC8LQuh8qRPwVt3iyxMvQzTGGLLJbsSNjoWpHk4ioJpsibTtMuxyQD74re/qjZ
U2zLiFlDZOe0mZAJOmi/6RhaZXeAVwd8mApX6bCtih5kPiTj91vzgrkMveT6KZLlG3yEZQGPIA85
DCerErgJvByVD0u9mgiz+ML/VAX+6F6IlORV70Izxv1ejYKSm+dcZsA90w+ah/kE9nnL+xvu4Ep7
EM9DkPz0RPfXascCRkwQuw4af2Q8A0AnOTq/aFYmVDi4V4ufkHHdv+UUdSv9XuGBRMY1ZoCRhL4f
DIl2aIsRBXl4o1uubcpVnHz19CwjsoDmt2n7/aOiYq23SPvW3T9d+E6Vi0Bb9BzFjWbZ0nHRYZTZ
D1Yk3zfCLMt3UEaPGFQ/G8CtJnzIjC8kwYe5W64G35Czra7Wy9KfiyyIeCIqfD0PjZNRnqOghKWx
DaZBrrOs5omXlKIwbP86LAcoZardTVDNHlP3IqRzndk7gnm1ExnV/5jLYmUTlDr8uzUQI0k70/ar
Rl0o3GZ77QLkcDH5Il/5mDl1s9NalNMetRrSl916Y1SipLpM3dv4hzHTlvNi1spBraAFIYdHpMio
RA9ymIC2jDNz2iEQmDt9row0DPLbj8ki9oHBoNUY9R2knWe+LQeZ/dy2HgOmcYnz6xlwik2lSnUA
FmDSpn/E32z8vopADlU12z6p+0+52MKHDARPlLtMW8uCGh8o8xnH4pHH60aeI5T1E5iZIzkSNRwi
uHyW9dVCG/YD6AhFb362cT1dzpZ4Ru5tPKltmggIhx4G5tKBGMGb5yohN/Zc/Xxt5+QGBa+U0Xku
rLoGlQ8ogDaIhbpQrmKYJLSufGvFe6V8P5HBKAZk8wab/eimku1UvwyRPJL95Uny0eiX1c/c9IUm
AcGnz7fonSeGK35UAFUN2gz8P500qMtdaWvZ00vpAunuxDVIOjeS473lVoWuyeS9CK2ZtuBlmc/v
EL4gr0XxQpakpsRdYaFLRnbEKiwWrsAeA/jUoaOtiT5yjnFT8LlYmr1540tsYycP4Zt3S7L7E+mU
nBLtewWwDVfLEj3uYztjqktO9yNmV8wtgFynXqcBdvORz5M9pRLqUIg+BF6/IaUfjfWY35bSYE0o
lXPNF+UP36ul2Hb2tgO7f8e5ftfdU5bYB4SJVubBNXHfPYTSTWdJJId4A9+om/sPTFRScRqxfLCU
kinuPBgrcIrurnGZfx4/iY/cQas52dfoY9nyZ735bNGbFCC7RMc5Aw511YDegPAQFRfMd0a+WroW
KA4JPvIVZe1G/E2avvIlfslWfMsXe4mtaoTJXAxgnhp1Kiu8HqbySYMBkoXcloGY4PerbRrlQ/GP
zua95Q4KqrTqDvQ59NKngBw+MP9Y5+i/WCnvz4gZEDp4bXo5fVKrsqyT1AkSqYVjfF8vC7kxMJvl
VtsO2iamAiYfEam0q/BQg5gvAEMoRukHgq/ulRw1b3fWqoCsUaHY+vShmIYz2vpF7KgJaG50j5/o
ekJ174hoAoXd/B9NfS0aVleeq617WU0CBLyUb15zA05C9f4ud5XGn/FuljVpcLQXI/hy+BSHQPOy
m1qFxwW8PsyjG+/qva8ZIj2/WpVHHHT/1YuxaPIUgNsgYpRo6tDE+D/nLNSCupuP6pmYplzz4ugk
srMFBE4Hs1keBEVnXkWEATnpc99UA5n0fVKGf6WOgEKTx7hlEmpjziPoQI+8Jbo/gFX7JNfgDDm+
Qo1yR7V8gsttgWp9o5NFYgslBArnAV+1zd/+IHI1K5SCWN4rveJp5s5RulfEzf2NU9jfE807yzQX
Dd9RnCI09KKgUVGxr5bicEeq+Q0faG4LJv1bAjO8ASd3LH6Oe/NXkWTDmVGUrdD77Za+AOz++UHP
k0whEpY4HghTMOB2R491LkNs/IIyfFSsMAeDSMYNMHi+zx6apGKZB+NTMyxPIg6/5N1VO2/bzuRd
XcvuSZaYl9pxnoJ1q6cyn4ThwD7jkE34Sub/S3hHlvmH1BO/Gx1cGK4fICTadX5JpPcBQHS5CbSu
NAKIJm1qnkhPTXdMHL/crG/kosUwnkL9XmUIDJm/f1q8K/lECtitir8wsJlj+TjM1lstDAqK25Ho
o8Sf9SZYIMOwQ5LU6/11PFOx40hm5WEvZUNajyN9zfZ/X9RwpRawIoGo2xxU/pbN1SQomGS4OH2D
bW3kIGrkW5RxJE6amQRnT+94QQHjvjuL8jePyn1XkASbnzy3tqyonCDmGh9LFeV2+ouBoUvGYcpz
cd16fXW6Uot0MKoj/GnkSZ2iPqAm7Y1gbpk6q2WdS5YRpmPzzV6Ndv+QOZMlnQ6o0CsM9pga7YFs
yLypcTMrmhqN35vtnN4/OIQ0fTJif2b5a58Zu6I3oY+nxfq6O8PhLBcL5A+3qQwQDBdSY433RJ7M
4vL0T47h1mQaBJNpYlTkEOhrK+eP3loCpJWhqzoqV6WVYgm+AaaAnXZg3l+nUiVbkswe8D6RmBqa
py4IpeQ2o3iLEzoVjFB+IXL9FtSzWaM1EYS59qClGueCiVt4m3ueKnEJWP9/5rj9PodX4l6beHPE
mgoF81+OL2RBuH7Ala5MSxXkyhQeILZ939X/17gqUwmoJjHQkAlzyLjKO5AAte2vB13fPN7i5PDz
kPvbV9udmYz2XW+1vfABsxhuHo/iRE1Hg0hw02h6bD+kMSSFmOnzYYHk/QVcJLi7zAAVfPoNINOT
Jhz2WygPxauJ9tKy1zjY30NtIwbjpcOyB4pMWDBNcQRDM35tvVOO6xx/Vqr1yB4H5i3aqlAV3ZTy
thICmuMrlVL8J/6Z5aoxyWDVZMpF4Rav0sG2vcZLWgo2K5Pq0HYkByvhtISvjWX5SQB/jZ63Hl9O
/9j7PMqszwBxK82rVR3W6M7sDpmjlCMWPK6gV+JgLY+xPncFGvvwyDICi872de9Ex5awZ0FqJFYw
4KLAmqvVpkFO1pWDnTVUH+wp9rXWtWNIMEzmDL3FZBE7NW5tCsIrgr5aYx/1yFUMylSrR9tVnRCF
z+0NvI2V3YFnZp26woZGisZuMDIFv6XoWDjRbl3L5dg9P5xtfXDmXYkRCG2wVfQu/MWemDIqicjB
OAoh+uDGEl07UBaZqOiIZh0kpTzMc+fWIncMmDETmZgOvuEXkD0tmuVx9elBn279lc8FS05JWMRF
jpUrLjRcbQx+9OqpAcL40/lP1hy3eAnUhr4uYXx0LuVTP0jIS8prSLWTGs/fYPiR0WlJ3s8vNQ69
7/Hch7/0529CnLQzgHD2QWjnk7xs7SuFk0ymwOJnYSwOukIHJn6Azo/0nIdJT9ixlzOo5aQofhQV
5t6+UTsGT0s4M2YkQKLzSFxRbx9DZsjRwcP1a5macMn2M2jjoiRGP2AMAdeknKksM+15cqDzaZS7
YVmC+bru4UFkhwfeaueyQOXD2rS0SbxqVutxWH+h2gJfCpFyi8MyT1yzVInTFjw1WqTNptG/81Sj
d68RIhlKmfFSPk5m1so/hDNLISXRVcd1WXAxsFGCAvp52gr9Fi12maNCCfGpYnK4yVTOtVIy2JKx
ny2AaxcKpoSbhJHmJeyQGlV+Rxjvm3QNVkKWXuBKKMNhZNUFgTxitRiUgxwQ9S5Rgii6qhrTN9nn
D/9cfkeTnS6/WSihxAsXxdKjBnmucejCDJF4Us+jAW0FE/knAjBungy5OsM9CISQfbF6auO44OnY
V0iGObivt9OCWPVXwk9XFET597SQZCsElqOODGQBUP3l51BzyMmAiXtT/yhrKlQWqParpIT0usDl
GhTrsHIGOcuF3okOIDK/c0nAsSCJp11uNT5b4u4OFIYGvKYQ96EKsjArH73z7U3fERekXcl94vPJ
aWwp/izTarROsZvgQcooWd/CANRbHImEPWGt8579WVXlXF0ws8SFHiIZ6Ut2/giItYEjTVuJzTbc
cEnNS/lPup3wO/LWQ+lnOM8okbrXMgdopG+YB7UcpyLTjxZDXmU/4OSw1xzOLJrHyu60aRjd8K2s
562SCeMRSdG+sLad/biXIbk8oRqWT//APnbe99zUn8j7vCSiA/gAHVMaPdm23EfVAVryJ6xgQk+6
m254/G7Hv3+Bh5wT10D0BtgLfoRcSFGRC2xuXUa1cuu065WOi3LkQkStry4wVGfnuh0UmGYXwDJW
Yi/JJkLHbsD2iE3VXu2Q9DMCIOznN7UWmrC+zQtoDB2sWA/wtaZzsaqo0x/yu9UBQTTBYeKpC/7x
ECalRrApLF9Uz86jdC8a5KBn93ZUPOQ5TCUQiLswhyZqbyqCb36Abe2/+PJfH7UZCc38SLvoL9BV
lneaiCgc6KXbVQrN8J27Hmw2jy7+AJf26gT9zdWcRXJtcS+sAiNLFZ955zvECx20PdifGiWtm0S+
ipERRLk7s+tk6VRmLvn3sJ95xJN+qOe6wWg38qZn137JiNJN3a8MK5XrenSM9ufSve9I+XsKuh2h
iuvTQNet1E4xmk1jPaZ+1GjUOcOWUEH9A7h8T/mXFffTz4YsOAhldZBEcD8ZHvjD2UyNtK4k8mIc
WvLErejM7WUhQ9l6rFDcWvbmxud0rL7WB4o5HbcJHUjOWiV6yubHFrB41u+FpanlBtnRho0Hghus
nDk7RIoq29hwrQRxVD1CfNObF0g/eX9gPMUE1/0NAY+lBKgcKQwiZLEwD7bqjGabNV6FjHDuMX46
jk8Z6rcrzgvpp0y4UwFV3RCExujxyWri7n8vj8KeQaIagB7zCYRLYet9PCPslc/fGZJg8JOBA1Li
SV39iMYv8IVAD4uOL65V0NL6qY6F8tQmiKyDYTvBWed22B4xjpPXa2Mj2w02da8BuiqjOHOZSZX9
AB9xKEPYOXb1c2DaDwyN2e7AmAg/SUMN4O1I9cNbBYXwhHXfepx7/DzaD6A9+8UukwJvFSNK3MkL
SFqkW0PDi7owgw8gtAbW6RwglkAF+yjd4oR6PggSRqzRZ/MbGh/8yVIkE+GzYaagAckCWXoA0h16
Tv5/K1vZ/boM104krnvGNVwlpApwzzQ96/KJb6O92wsxDghCmJV/YL6AGBZ50mPzpYJl/c5FQtPA
GC9TygPOup/Vojs5nyQE0tgLsSL179PGSWtQ5G/uSlAV/vyraAL+EtMK+qtsebolFHCSwUyvhY54
bdmF9F403+2csNfRxkPgrjKUYbT+NqopbDU142HIxenis0bv1/FewPOFm9k5BhUKk17c6rP+Nnsc
zyT0CYHCBlRZaiAh4PADeGZ/swBBw9wZ9sTb2tz0Lwj0ksmBtR9f8JDtpTgYCY4iceDOqjANA3VN
dzrr300aUmkD/16yTzv/E2pk3+Qr7cqUvT+113Hfs7Z6/TYtDzCk5x216VeSAOGxoXwK94mzqTUn
fnMQ+B8SmhbtTk3mwiIeIrgbsHyO8mj5dpjZXBmOWD9fPQac649ifX8eilXsFjY+xegfz8bdh4iB
Kqvx67dGn9P38K8pohUqKifmRVksnIt3dbzW585ApZ0zz4ukZXpXpRH6vRaJBybP6ypS+/tAa5AG
lwXfaz5d+BWKl/Eva4Ec5FSPLUvBiYZHQEi0/CYsjkysNNJdEEZ8QkgNCjWx9P20y4cJ8VO5KtaA
aJFz7bN4Zdaa1l7bzrRzIHpOqRcWI4sYGEPsQzH06gmNgnbJkcljWD3tey1DZmtqG2lDAX88I6mJ
7JKH8WQnGSQtQqLsZL0nk+iqGlXC3GrzWZEgjDXiTXz3oRXBak64LqwPCDo3p1fS2JEXEKSpRShH
fth/49kBhphmcxcr2ETVfVtE5ZZx9UMcu5+KHJ6AKg0iIMRshVrWlOsGigbmxOsha3FOVOHskDHY
w8PD6q4vtw0MJ2J638k+/RWvZzHLF9BOu4Rcomgy5jIuz7T/WnfsutpILqAIVRcnIof/MLXeLoJV
p377vRc7BkXOXfcxr+HkOeZVcKNzWOqhhZlrmfWIsyF4AZ2aefTV9QT909MSk0GvlZUpTNnM4EbY
q7NGgJyWttmaQ/FKbC9ZVmKy5VOwRVdABEhPSo6sSp86k8bfdytU4Mqy4mEwRHmOpUdXQFNIgMXn
Lpov/OC3XZwufYpxAI1ABNq1KKxCFTp+peyl6m7EXU7mOQBSQcaRS2zGMAx7seCwCXPhpEUS6Oud
RbhTxt1X/1TUsvom6HUB7czEPWdfA3nZCqkJdiL0WNK+q/4iSMmSIKGoWlCwVB8ziD0fc6c0pyoZ
UTf5LMky9w3bh4kP8ThCL9YjFjdwKcHyqvKInIWImcqYWmPV9HBxh/D5QMxRuOkXb14gCTXFxOxs
AEEyzBRoBjnLb8xKaVntLGx8FTFiel7Sme3hmNWMIGkjzj9j2EAp7AE4/RTjG4cx7GIz+3tMQlvm
x1U3YHceofnEhzDlbWHzkVs3XGeUWdx1jhVsxWbt6FG3Vo8pSZRucj+JJ9jLYhDU3jxtkA5ELLfL
gWQgUfrPtkOsQVX0dMvke3/QG9jLkPGAGSP7BX7HiMzER0Z6dCG0QRcfc/qnlP+c+2jDNba54CE/
jWYtCwi0d/+IriqN075w5JRC0ZoObit+dznXRcdPvgmhrBtDc4o3E88fyp5lAegAJKXfI7X6oNgt
3/qABhVwvSO27iJIcljxXhhwOuzcnOssrKl5rL/Lt81lKyAXSM7r66omN0QSaGky1zgsJ8a/DUi0
4TzPfDcmutMytTfJ1Jn9yTiwy/2QkrtnI3Tdw8Q41Zls0ue/AfoVkB7hAIpl1/Yv1QraATGsl6hS
UbDV89scxv0AHauunhivorrS3oOS2H62WgZX1W9Nu8q2J5NaJkzo2VGzTJ5prb6ee1G5EFp7GoQZ
3MqGcs7E6ArT02NnVDuXAl69CDOrwloi3LRVPVPpKXsgypAB2oIir5YxY+JfQ6fJz59LwCPbxhVb
uKmCvVBZUB9lTTEFFJ7izxPeiKdfBusIuPiJHoAfH0YLKzAYHqKOcGV033oSixuC2gxD07/6mDON
Cr8zEC+bpJy4Ca/RHkBD+WqURrO3qfqe4eiJq2hAtojxbOdCrH0KjnX6hPLTzUhjFhGpSM9wnyBz
5AQ/xJjDofmdJRMKjDbWUPmJs/Xc3Ba5hMxhLAMkR68caL5HD8mLyTUNmolHXB+TAvjwA3YJcPhb
rq7tgl+DYL0KKTNBa0+0HQ4frBTn2Ak4L1wxLDMR3BRvdk2dip9pgWJznHqsUzQVgV88szIfVVI+
trO+J/KOpqCEAcFfzRtprSs/oAE97uQZtUoJPDaC+7bzSeWTeqq5IsElIx6VRSqxBffXs7GK/pQR
3FttbEwklVRbw23Os8OIzBage6WXMsnsT/SDD3Z8YbYiDxsS1zb+uiyRIvMfdQeaiEl2C4IljItL
wvyAKAxfjCG8nn7egycIDiozVMA4dK5O3FZybHcm7FbY/ATKn+sfvZ8ZEROZMTxW2KP6Fao93uGH
RB+Uus4zLoMZCeqVXTNt8Vl80i9sdIBTWBWdrR4wBXzQCmkeCC0j60qAdYOMVUKxJUnVUmjll4Wm
hORikh5Fg2UYqWEU83bOzrCA/PHtsLDha/LWDsCWHLG3ONSkzLtHC3Lradc8oqU1JhMojygIUa5L
wbffgmN3aiPbve4Z1pwAEpU1XJS/frDHb2WmRqZjGsjDE/nbTFbZsEEPyTrHrz0v7rrP6i2Eix8e
B3ovvQIcxqdmoNDGCfFT9l7cK3njM3VUS3tVNmvqaEHLXWU533cO1QENLU2pIVVyvOVIfr5Mdx4U
UmTHga5exZtq77wqJOuHEVhnx138s4EoBW3aFuL6CW/LO6c621ccafciyc1Z7xe96IoIokXRcM1H
bH5acUcYbjOfoamI+R65vuyBt6iuElHP7YoSuCvLpDPnxwwDAtPr7DLfLnWr64awLPmDkRmOLTLq
2RE9BLzXm3BwNotgPRtH3v6vu0jJWe2WcGMuYaijNZG/kyb/IOOCWVZC7KLrZOn9/CbMVk3rIW8N
6y+UAEbrA2MjYkCqjnZ80VWrhdacSo01LKFTGK6YAlkr506TtqDSZRHVgRvQu/rtFPozqZ3jMquf
bELt5Eb10ZAfvQD4qmdU4hMB9ec43WSyAJtIrcv1qwCLjJXUEL85IWFVVEFDkbvIemd69N0n4MbZ
4wI4fjREURjROiir5wvKCZHSr7WDwncNge39ox2fGuhtNwJkls1zRdS7fNnuGk9ZKJCh94d2REHc
aWNZD9a0IQwgloAeNy3WiSmlPdEu1ewCn2XN6ih8w2jM/gNFOoukUCQr7MGg9FRCuG+fwu/zk/jm
f/13XRHgFaePzIZ2G5dliRUUKRkh8tUdmij5CAKgrOb69K3syj+VGS4luvzofwdp63AlTNvUEL9F
C9fsWo3ZrL926I1CIqavvt0M2w29+aAFEuqJTuoogFXszHmfgCacC9R62m41f88aUGXCe3n7QZD0
gmduj5Qdsc8KeYD3bUlFgKHnR8m6qz08gZeOJbGZlaFkeKKVWS2pGOBmFz4rw7D5H2iK96oXex2c
PTFNaPhMKfBlHETjGLaz0iEdHx00vaZyni/p7wXvuCbnsa9QlkEGQvo1XYTvZLSvP7W9t/DJbHs+
xJOkecnSmWa0k8SwulbCpaMdCY+kV1lwJFPgvQHbkA2kJXcI82UHBN55BxVfFrV6dgU9UAhDzkcO
k6Xog4uQZh7kinMw/vE3BP45mcJ7UaNP8+a2099xEPu+bzMo0+rsEg+xspTujfsMfRbOyV7Sen7F
Fgu5K2JUTtmWuGJ/GdE3yr/MCh/SpthukssnGVxw11Oj66YlX658aeNGQevxrnMaXEYx7h3pexEB
k87bjjwd/ZXke2Nv6fyfCjt/YIcSXL63xkrzYrfRVeLfsReJ4zEIPjs2hy4zDxi+YIgDBoCUMx8+
I0EVA6ASxgaGksU/3RkEQXxtKfFA8wLulyyUEeW+ZEsleiIinwumFvD+SIJZA/WwwIHWtzPl0LYO
TDJUKPjG/WndA2k2Yp1uoYaTXRhOdIZzNL+P6zXIRJuVtEYFulo3/juAPbyb8gmk2kPmA7vp6XCa
06KwsGBB9E/5jviHag8fePruVT7j5deS3+pF2SiKJNLRSS0qgXASOmrgSfWvHFzhEeufVJtfk4TD
92K7E0Glxl9Ra8/a/CNW++ZEgsseudQFywgbljO+anSYXRfi4OmGx+0mMqGXS4okOd6YYvEEDqK2
SV1oe6AQ9IAIsRyz8xjFZojNCGlEnDUoUh9FRNt5PSmxNa1l5vfbmNS4gmQXvPanU00WNrQJMKr3
vpkf04E5ENc2mLWg3nhOHxTDTbNtyZb91W0yP+I3LOwbbsPzUKQiGSVLQ1eLOBOwf0uzDmnPMqIP
FmpjGHi137FF9hseeCVbChaXc5VX06KJmJ9CQlA2EoHDuz87KvyIoMC3CY8M8TVz6CDGeQzoiZ5L
howkSmZGAGZFBqZLXXawGcqQ0y6XriMF+21zLOJEmdoray8gH5HY0PEtyjU/CH7XzjAUrAZWEjib
ZSaHevvlAO5gn/dTQSoiVw4wW6lDybHcS2hgHyJpG6lTCNEJkDT096F9t+oRI4kUFQp2ZksegfZb
gRidrDmgCuNgsbR3XnQRupu5jgUpO2/RjfFuVJdZq+tUem/YXaGROo0ig7Es8xwNcFGS1QrciI8V
IMfDnyQxTcG4iuejT9miT/d3tLsLx9jQtjBLrLsF/sP8oKzwLTfns7v5ettrXV/L2kholB3VgcLW
kjdJAhm/rSsF2wvWKcomcN8FgQH0h61AwvPxK0uB1KJO1nRMM+FN1XxjRQBd12YZyzs2asqa0kNO
2JbgTzTJ4mMg6yid7g6BftSXtOwpAPAIxLUWcLGODJncYOuxpaHyxa/14O13lgeGnPO0OWqKlXaC
FSb60KZhDVaWb4+guACUJVd9LkYonqlXN1DBLEoyFuYIVguqcnWv0Jax3+X+YwCoCRxBBtooptYI
UIgDB+mMHEp9+4RqJlVtDyl6VNCBU5cx/dcbzrt1VxkH9JJQgppbkUJzxUUxuQCJu1+R8B3K/h8I
/+/HRKf+ngOJYww3+KwdpuNxqziVmi5/VDhVh8j/83I074coZswy9Bvi0Po7PCdagsa3ec30lPoD
Z30Ha1YLvlOUjzzPTFuDjE1ba9gn5ntSpP6RinFM5QGKv+5ZaqrT/bbVPJdtV6G/qiBz5vFZC/CI
sMkL2MjCMifRgXT2uiJpjrIxooUKJ08VyZPOVo51NCtt2g2timLCMAluXDUNG+fwmo3Ug+0rf59f
H4MXcVJ4+LC8ilUgreYWhuHyt3znFZcdE886K2U9TSlmbZvCDRcMSlbX5S8yNpa5qwNhkh+sl2PV
gvNk+Y9BkvMi3rU7lwmrSXbTG07EPDQiWmk0+GHMU+NVlqQBuTD/eqhk67C2Kq1JT/aHVfyN0E8K
c4swLc38R683w7SDlBLeaajmU+CfDHFMJniCMbl21SFcKUcQiWlvP9yIA/VWcp6CVuKPiwy+OdMY
3kHtJ6ZfC7ORcioWqGB+iCC4uCfXhk1Y0nSl4CIUpUZBq+dT0O5XTDw/ccJtHQto+5K3x9cWorRn
/CSkUgZYHgXlg7Ta/u/lclZHG2fKbHHopMA58vNg6rRxXIOuBg7Q99Q34zhTJ5cVeNpYTUmtx1u/
d8jowYnjzx4/dEsZ/CKyAtWCG4qYxfbEI4ysAVjBpDgjSYKLV6GNxNPyQ3khHBnqgcE9p9gVLgV4
DjpJWbelBTYLzgblT9SaNOue8oJLTZfqZLy48he74Wnl+aGNdjDGd5yYZLsstgDuyxFOj9j56BaB
cxhxQcMkVv1tu5O/+TaRW1QRCMqoWN687pYrRobkXjis58skAYyWXsYoWfZgRGZwzQKiAWtUzKOr
8W+YehXNBbAvgmw1AEhhTx9087q8Kcs/IUme+df0wtTVVMmFmqmIObgULLyQ7koN65DeoyL0B/xE
GQmMOPxT8ztQ53Prlt2yo6YUK/N9CN64i9qVZSQfWr4R7Is1gq5MvHNKi4dE0JSgGm0FRo5JOpLN
wNGdjW3XlTCLEXcrCRnAYa6Emax6RgNz47b2kjhhlMV2IfdWm61JMpZVkd0UKsYKuff76+nU9YO9
VTpNTr3KyNKrzLRBC06jAODv1ltMYqUyXIfR9nGdiGAc7/FEI18G5628r+vqkj0cUyG0MBucqOji
FrcAxHPJZJ9NyvcMjaOK8DWiRYZ4QYzFrRSNFRfQf5l96mdvYhbdfdBt2U56X15hBgWJtD0HIY8B
K6mED9sNtpA6nwlXC4tvfxoUz32PdLIaGqcghdliATMWG3cFj6AJqwZmiIRO5yeFm9DUT6M+KSVk
H7UxYqjAI6KBdG5cT93aAVCmUrF7EEpUyYc6LwjysW6xKKI1yR+PB38UF8CJJ134hIXWk/C0+GdX
qdmMzoYVTFhJndV+dG2Mp/bQvrIJmtXLyp9v1zbXLQ2WI01NhS8Ue2ddG6zhjeEAwlEwF3S3wHQI
MeftDP1phaOozT96dV5uF7edi1SdjBirwFWyFF5Ss7twqxcen9yUJhk+gZpUQ4/FkB48nMh4TUlc
fd+OTbJVmU+1oHhjEoAM7JSVojmHjSZFdcY2IisUApG/0SJ0vsmdo4lwlbyGEkhBTo5ssZsvCUGS
+Ew43fCfJYLajMOrrzmHiH0aTIRxlhQNTLhmk3VMKJ9JJSmZ4OtnHtJ9+Gm1b1VZP1Er5vRkuezP
PsG7wNuCZJzCZlHktIlffXdYatTxri/adX1hegUzoyxfF51xKf3GuqQK41ttvujKxH7/ijBj0HDx
l5Ryp2hxZSm0Pj89bT+zbh0y2hl9naDXeI6lCG4rgtO2mo2P3e3gdXThJ0O+DphcTi57MJChMYqr
Orl66jo4GsdZv9lnGUskCXm4OrekV1E1XrzI7/ZlcbU+m1knvsqXIX+ylfNUPahGJKk4DyWXYWqJ
B1FTqFCL2qP7vcw3x4XYhrK/QjXqgtNQ/IddLKOduUTJZGZISNaMMGbCiuxrcDQ7z/lz7sy+vBqQ
aY0HChCMLAGnydyy0YHcF9PtX0nYlmtNrIaIyfDiLzfvUwUQj3QPF+WcoTfTWq80f6lCOZlX1pvt
FeQobDhYXakgpApMHqykW9kjFM7Nwf0zWBDBzyd+e2XgVj0Tz+XxuAqWaXN7ZPkvgnS6BUjD79Eb
g3trcLsOmk4NyVTPE5HXws97wPt12WMVLKQXwuv8HvITFYlLtrnnuipJk4FB7j4aaXwD8BeDf5iC
PfjGwjBoRAQ4b9zUpiUgz+z3DtG1jW4iiV22+VQTzPO9JpexwnfSwTEjhMunr3DhvaITZKS1ivPh
+Vaf331sp5sXpE65gT4kLzkDOCCcK0C7ner0aXReWNf8NpM6AdNC4jr1TyRooW+alh1RDY/+hDbz
jd+d84TFY7rCjHn9OGzVkvbUloXB3o3H9dj7QUG89cFaXezUGD1V+3qAf7p6gejvC7+1C/+2lnY4
60i1qKUoc4P6Vxx3pDbKNWZATplkChhnrxugvWZU6Si59s59WTUpVX5KSO8Vq+MYWZkSjg/ZTQj4
wtocfaIc0xQKHo17391V3l/BEfvvR+P3eHhtE/3A+EMVy8rRJLChnCfLQ3rj1vO1mSkLDThfY6aD
2Nr1oJERu/J94nY6YbRC++iAvGHSLRLgwGskRUdM8Ad8SQJYGAoq6Yk91MAFOkLgAcZ7ma6iNmG9
Ie4+tvHEBFKXVOSPwbHrz/6bPfy2Y8dbDB0xf6jKyZ16ri6LMovSgUtEkH97dD4laMML1wR8g6Ga
KClhae094rdGtMRI0ulI3yXB7d8wIGKZSKdJh+FvFMYrQGjV5gbe2kbZPoREeZfBuqshgjJoCoj3
K7wjYGivT4q38lEAN4SotJl/Yh2Jta6uFOqP0i2KsYWM3xyDEqTzpuTcuLd/KAbd2O8vpYDZ1Nhn
SvPYrmMCdJ8ikFff6kdWXS4FM4lOjDPSny20cP/AUVSFc/IVk9ECksHhAKHHaIAhmFfOGcZL5e+b
HAVEkkOpuFwkkri4NG38zULiXgZtMPG94NHGvec9xFCfrGQCvNxfR5F1e7bKQOk4hLUslUVDPRfT
tb5wOih25S0cP86YAigydT+h7tnDzoMBBi1AOH3X+DSIBE6D6FjdGtACc8ZrVm0PV/wfqMf7bWo5
s0+bz94DfLsNtA2OJm7gICMBRhbgshyScQIiaG0EQn7HV/hiIr5K3zQnGwLer9Sq8shEsm2Klknp
l0+0UHWg5OF8jCLo0dS8dxoTMSY9AaHzdQJBl1+iiYBvaV+NTU5PF8DaOViU3LHbaKIe1NMpgjuM
nphgQfHTcxAmAO3SElkmcISeOZHSfEiEJr4xoEplfSzxEDxfdvKXO1nowfbZ/hIZQ1mJ9PYo9eZn
dw1YzrMch17qOQEDQw1EzPTb2V1uQi2UGiqNUU/QPKhKPY+tJewaCAmOGQP/u/dU2oej0d2pf3PV
qNFs0eULlCfUxbpn91oxzjgVhOsjDBJXIk0xIBplxf8zYYANJYH14KHokx2GCg/sUkr93IoN750H
uDnJoFh1cwHjFQI9/6w3Pfqt+3OToORvS1yL403q3WCBV03tAmA3MWIjooVPAASUBV/9FAJg/g3v
IvnLU+EEYOpmys0TPDAkh/UH6vSdnUciWG0tHXXzuza3wXM3I0VGnAkIH+CU1wjRaIPMJzpUGJ65
gos4WsmUfJp9oaaiw+UpG2yoibgTh6fliFKdzWD4CSJaM4pFDRmICtIF2gQ5AjL7r3eitJF5pTpv
na1X0ps4NkcHleM/OlKJMI71nc/JRQCwLzGyBPAwv7Z3eu9L8HpgxWZFOBOd0sDgUX24RqKvkqEI
TvpL+SInoCs74jL8qLXKuftCHS6pKBoMwnSCknQHWRBFbNhBynqFiOGpZMW/Fw/gdbCA7swbAAxI
lCVgCiqlt9S1iJTXuuWF5B/TMjjhMhobapmiCJT+qoOCMJVO0uScKVBAzkdgLxKZqH0JOg9cxord
PiN57RVtpXAcblZZShOUvWlbhIqW8K9iow8fdP3TbPnI8wfJQNXDdr1012PqxZTb2YdrSQ/h/x77
B+74p5+tm+SyHYA3sSURh4eyckBJO761owYVbWMNmOowFxG2thfE2OnClF7oYw1Uoh5KGS5no7RP
eaTSkdYHgsMBx+3SUKhfQbXHVnu4o4HMXEZ1tH5B+zUoyleFY36zlqjDxv5UwXhHOrNrZp6aT+Zc
S+qr8/Kz51Og+GDg3ISJKiZXrcWPlfRZrt2KgJiZQ5kMnM5fH1dd5c2MgzIv+CkqlXFCaV1+5GSq
Y1b7GXM6l3jljcTbY3s1oStBYTZprOYF+PqE8UcwNFyVAW6GwvbBK1Nv9OQE2c81b+V4jHtcA4pV
wIWi6w7NUHj0QeBPvgm2sU12BeikVFoXZNDrZ+aYWT+UP34PGW9LW6SXWJvJZiUiROw2Y/pWadPW
/Ye2GeOR+RT3vZlZxIipHKCkNr2pj1TwkEKdTcn8GvUX5jQ7LTiXyWoCZGMeXjPFGF5afKJtUYqI
97xolVfXFJyHK5Cvp+exil7l6Q+atC6atQiIx47E8F3wwBNX6pBxokaOwDVXvWBBj2680C58f/64
v+h/3/KVHOnIVyaCowZhipJRFbcgI/jbW/vTfa8hoEV3hh+rtBggCuFIBH9uEh23cTVjBdj4GgRc
PWxUqEMqTGwLNFGJMEnAGeOVMMih6A2IC+8NahT0CIUJNatUsfRleHPmoTO5pYkrDm8VDZI5aPSQ
wVUqM0yO1AT34+Q/2436D1yNUE6Xmnp5kcmpjKIUsx2vrBCUEEZK6UteNdEMgkevDd6PVxxHkNxq
3t0OmtflEjoJBIbfEmjeRX/JY8j9DIf+GeZ8FjLVwABP8/8B/2jVup2bKpiolZhSqvQA02D82vfv
fhtuJL/X8yaOjOEGMfRIvNyzl2m9vStZ5ZnYt9UU8Q4FqUqpno+hnwv1hnzviQmE9LaXoSvQVay6
o/ONKqw++BXKUpBEdT6Ieg6GVB0BPKN8Wqz/kM7KMSRAK0bYIYhXJhukY/nYo9Vh8PCvzXHG7Xci
dO8B+tyBChbI91i4mrHEhXEH8yS1kntgX0jGnmy+hRfJUXWSDxEC5FUC7iPXLi4Kcz0cFIQpK6qk
l4uBG+1yjXSQFAq/sp4x9FOVlkefxKD/3BCHlCkbHrnoYa7g1T7JcPm1DrSNZwcF5WFHKWD+2J6R
l+/trOITjfoeQXBK2Pzs3KvfVij4lHckWVcNcb6pS8C8s0MKBtM/jiqjWTM2WeQnPf1Vphcz0ZJ5
cMVvwRzwgl48n40J85/kJIpZN4MSPpV6ZpU/w3l6GP0sxzeFJzA3TmjciEXifeUU1oQVRnpY2WsA
Ti3RppzT17EXGBB4biv1LandP8Pz4VnaM4gEfza12ZyoXb5ykSGYZQ2wTOzjX4HTdud7W2fOwejd
owE3ww9DPT7hBTNCd1L6iOKtpIJYlm+k0EfsiptkalBexmGU3blERbp3mJXeMKHEpByD5Jgoqhzg
2/pgN3ipo3JB1nuUOO8AkG6SCEdRT7PnzFtqpo8El6OdjbfU+EVzG4DHxrxjyQIkrgu369ZBdy+S
U8uajqjpd9d/V1b7vJOwHe94YRJ8WiuCN9pQRCBiMh+dCvyVVhh052EDGgiNbWRa8o5BR+kPmHju
TXKV593OEA4dW4L0xe70KuW77qs8pCUywjLNP8NmLbpUGGLqdxFJ7HiZBKIhUSRSlRXZIT3K+MZ1
2GmhcCcEmNHgmNRhiZgB1ZN+0UL5dS+uSQpaWEl1KJ3ficJwAI6R01I8G/W2dLQSld9d1La4yDNX
Eu8G7J5oH1Ks3dMx+xjo+lDAsnHaKWezVxf/XYbCJFX5NzRgTE8eHIdTyR+QkyCYHVjfyz3NyCKy
0+Heex94g2g3wOyLDNemO0JqnCk3FSlOcrZwOZ8PB7vQJZNyA2iAu8+2Zhc5DDLo1UwwI0GcHfvh
8xEn+Vg24Dgd2CGL+xp75fRW/gDVuuDVAyujjPWbvFzfVTJ7LwKCVOPAPvHv0Yf28I+q8yFPrAM2
GDg32QyAIeLOIeC8Y1HBHXuTu2+p4PsdzMpR+34j86PSd5KudLcru6gSwNCjoLCxwnU4JByS/kMs
zav7WkbGRluL03lRyx8GT6KpxDyNaJZ0hRrXbtuS2GtN9Js9zPK5sXF5lNjdtu/G9++/DZoHVPw/
AIaoit71t8gJ6PScW02fOzLm/hUNAnPzoUq/CQwJd0wscJibYgUyV3PBDNqh8eUXIZyZrob0p0m5
3lRCMqQeaaJd9b3knudYLz/v8XRW7XtvGKzWf1LjnWnW9cvNKRyJ/ME72S845sj9sUYKk8H9zMu4
BM99pr4lRfzMbEGIuStLV91exBv7n6IeXfshsPZ6xAvhb+JVtcbmPKxVjOkJtY87HJCHfkQDjqZ6
TKi3EIjIo1+bn0eBoXlctjKePsgFZRGmIVuGbsjr88WY9tOOwpfYGsHAs4EJKxa3SBEifeVVaBaj
AJtLt3wU9C8ZnkxhQqLxY2yxAy3qiXEbZswmGr9oJxlSQP8GQy2R53DKqeW6s+yoeN+rfuyAewT2
HIetuYds7jPE6DP/ZGjm38/3VDiY9gGRCQZnbwcX8hOYOHodkU6uKq7o9aCLEvkdRklMDps4iiIk
4/PDR70Tbv2y4/ATrh3jH44gsNm6HuqTJ4buCLmibf11IU2GudHUgLIIldzAAfnmTOvK/byki8zw
IbYqyHThJekb78GejvgpO3GUtUJxhYsW8neyNQOUEDD0E0pdSI4u9WAOaG3FqZHt/5Oh7VBKf5TM
3/96z4SBfFFfji21cvK/mheCm/Q+ZPC673OvIYA+2u9ygnsB45PmkFFYqQChFFvjBMZUPVhTXOXM
6Xviupx2BYJ1JWQLbcZbv37KkLWdmElsnVjjGKH7UUPdGmFYsLcMaHWmbsbY16S/ED1tNGPygZs/
yNFV8+ikbxP/UgIghMRarrZ/aCtuZYd7blzOY7+OpjUKw0zPOSZA336csRAcX6Je/s+Gmya/uFr1
eOg0bU+59uMV4NQ7S97jX0qqCgLpp4rZisFY4iq+INXFspx0oekqb5l91muVpU0DhVDDzFfdnLYo
tjeLBgbQGJQFFiGlJTAqYXncA9tih7I2/X6wpZ1BrBAUwmPkKq8PkFbNlN59tMgRlB/dZS2BmNo3
C3WpFqDh5HmsNIwxQNZ2V9narPEIBJV6pMYJ6HhyVVysVhEUA3FH77muzut8FN3nrGxs62ZCry7p
2801Vi0oONM+R93/izX4I80ITq37/XMLhiRZoKnIzsFQ8BoCM26xqlk/BVweDNDqHgTr1+M5QzY2
bxBwOhcpW1Dte+dVQ5SCTwTwnZhDGlYjroavnD1INQx97/mU58MryeUFZ+RhXeqtfe9/0HFrKRSG
9zB2vd172CQlolDm5rCXRjh7DLD7szw3a0/EBmtc2tWoroTiPokY2dXWHA6WdY6H3ClISYwn71K3
yvD9ZAu8t+IYWhF21smWq7AmzY/obmdTaeyclCJ52OUqJ64A5qOe0fnXQvyUmryKcW8YwGREtMgo
59xHoALgE3S20sn/s6bX2mYlTr/k+tq6leU5VbslWZPkn0ttUcJlG2Ak94gWouKDSVUvSaR1PYeM
HgPOknHSGuz+Dk12BSMK9oyZw3l04VhRsBtYOtV0BbHE6QzrPdEz8Fsu/NI1jhfKJeTz7P7CYJ0C
NPDxJXv6HpBOtioHfgbZ/6TgL4zoHLpG1HBBDQg9xNVQELbSB4GdV9kt68zq6FMwgx1+fh5bdt/R
jV8og/uJgl7g8szVv6CQ9Qco9AyOFvE0kJIKiac9GOfOG5+jHrw/yuq/B4fiTVpn6zKfMeXJOEzF
BF0NZh+FbkSr1OSiD/llmaKNi6L/HiYVdDWij1zXH5TWeQwUAMtB0+BeU8Ob6YPe2CMOBt78PqaH
NQzBhLzOScjUgTfRhTJgWHdePThT8Bo2ghFNzuU9wPsizloe9K7CRCZ3ga68H4+gnriMcAjHdi0g
UPoUBYlpuSFgi2wbwJsDgWr+Wy9wemrnCKNPlwW7ak4UlEuOd9Grl9+BFKm/Sc2k+vEEhY/59Ulq
KjUL8/8h21yJqPRjTVGSRLZcKW47LqGkW7ZXYMD+4hjag5sEAZqu7Ea+2CMydsUvo3vNtc/hsYTz
Qm5u75pOFQTqvEUYehKip+tsYK/mQfEbgCOdDvw2BevIh5yMnmCIDmY6scWWa7PDjxNJB95iNbhl
rVip2XpR2LQngZGOlxybVkHw/eXICyohQ7Dgb9xiwNqWZHFvzrcP2X5ZZ5GyVzCwgDWLp1UiZDJq
4yMqQ4rKKS6T0L15bR5+5rBWqqhIT29cbSrRoTP0UAzcA7bDtbZBTxcMcjgXwUGcrOwDkxWH11NV
tf20l1ccXOdtSvpMgSTLqVWzBgwq5JVRAFAcXFY2GlNvYLgvhyMpyJQYRo/5iQtYwYbOQ2D7kBgU
0Jaqk7EFiyaNuNHFL4iAT7ImIBnCInx2y2Gfup9c9czZBB6jPS8qbC9mxcvTHO9nOuyooyrHsZNl
qYJuAJJ/Zdxuqg00AdNjevivFUc3NQUyCLcJdpcbZdb4+06WSekX0pxc3yEz0hzUWLWOTJk9flWU
02J0XpPZk+eZDA/FAoVjsEwxkR5PMxTUdYGdM9xXu2BlXftgBKrH0cou2n6/Xp/zJK72eCIOwLzh
Gt2RgQnw7Vme3eg6o15K5MLk6MfjG8wAynMN8XKS9KWwgCLHXSH1jD//MiwznHSNFT0SHBA96SAL
smI2TkAF/B2AoBlyw7pJGdzH1sP/oWycUdZ/MCwhhV5dp0eiNivmA6xVRQ5GhXpdC82u+Cb5VigN
yuZ9f1R/0w0g3xrQlwpJrKTFwXJDdjBEP2ldW0QA222GeIXBgp9uyb9Qb2H6eqPZR+p1YdQCpDU2
YjHLUJmT2hwhb34vedzitONSulNVstFKtdXEadDSFzvy713ab3+NbJZMskPiS8EUYiNlqACs9J5D
Az1MxllEk3qnJKfENMInK+UE1XNxiZPxKMnHfGGPO2uDpTJd8Of8dJLnF26Cle9oIw74rI5TJnAh
h9RMdSMCnEpn5VH5TgG4eLAzM5lPzz2B9DaP+hF8V6UJXZWSnnt6dHF1KPAJanT467qJJLVPsUos
bdezKr/PIyqDHjsyuWBL5cwkq/e0Mei9+/Hmfo8vi9QSou9PT4cGGInfCHwEEICFsV8Oo67BjRpE
TtfmKWEji0epX2At5hRutclfzrgMLM5Bqnd4jw+1oMWLTsak4gDNQMHEYrFWHTuxD1ctyGl3cVtE
GqYNKP+CubksJZfi5XwUr63D2zgeWJxuwLlusUm7mMQE9qHCgFY9MeJYCiMVqiVRGQDXJfcFxX7C
N/rA15xBRFlc5i0rsBNADoaBkNrhcWnf9WG5DoGyelHELISh9sGLQLaSQlg40ZJiv4yGolcGCcP/
ZcywaerLx5d17zGaX4/w8FZRj1meyGvO3F/vLKKJAZzQIYQDRAPSrayft+SgBRx8BV/WtANyfv+C
hIUUhJU1C/je9wcH0l2djg1QU1mauSqVbMR8JnbijVFzJWc7b/J5R6NyKwHrQM8GtDyutetR4mwM
BoJrrpDLj4NZcPZ0d/M74qFVmT/pfqKgLqR4SoXrAgLbN/yRhLhKq+mGAMskUUk7EjjXTLGrMQC4
GFhbBtHVVIvcP3356dSwZ4vBIVaNk1dVBzXK5POIAnIyxpWZlamA1f5FUNUw98VxxLhF1jgbcMA7
NjDOescdEy9SHEda+5Js9arHVZ+6Q0YUjCSVpMOjx4ZL4ilHdkse83YinNenfOJK3SWRVdUDImGc
/clwbNOJV7GqELIGDoZjnGNSzvZgyPUJy07vlk8esh6/Fi/gJX2UTppOOl7CJZX8Jz7O8onVDXd7
05n563/ixzc8Osd0vo31Ph4qVMbNwqiK6eKjp76POgdN6k4E+TSIdfhe13/kX/I3dO2Iryh58wyx
BSTRv3ZjXy4Q3J4XYk0S1ApO5ZyNFC2O5nm03n8QppdwNpMqg+BuCDm/PSGM9qv0n5NHgF5r0Oat
5Sd3Ha15ZrBWfUJiGKCTtFn97E0h8gxVFIdWb4xZk7xlwGF5vSbUgjfTy5sbAvbDNhUf9BJwTpJD
yYimCLJKZ2pNr+DLS+y1JNcOqksD1e7+sT7+wr/XCj8tvT+hBZ0GJu7JQgUWL3yAZtpZ1UkAxDGR
Q3HWuF7Z7KDABuUYcRxVnjY+x5+Ymuk4KkI07jMBlXxks6vUwunAA1FTelOmYBNVj6v3yMl+tSJm
wFWk53SVxWhpgOGIs3iFxYuYjoxmplltt6HJsI1w+mjevx0pAYUAAYHmLChXiP2b/417KsLHgqbX
BXc/O1l45ZRypsjfG1nBHRAQJZRKS9pVmN8KM9Fsdzsw3SHZb6918+R/VJa7W/PBJ46Nqlj+Kvx4
2Xvh+ysRYGZqkEKDw2Qg8EZb+WkbZcWZEG5HycBZ9QgUQ9RA0gVFdga9cv/zrpMKxqqcV6Ne8har
wd/bDbnaGALL+T+84Lq9ZQd9I6szjnURct02sdQcqacedcETPVsQY4diIueyXkBXrdYuxr9CxKN7
cDNqtvGrcn7zI8+jU+Erfwvdvpko0JLP1rArOMnNnxFSsVwwjxI6LYJ9I8RxtZscgZDSCw0J1xz/
Z2zrCJVDZmtfEumBW3r3/AcFWf+qWnu/c2JN8efQA5MGACYtQNd1cJQDTmMMZD9u+f3/KTCKwu1+
CPEArOmIgPPsZU3TVAnxNlUHSfDxF5tjeGRhlMblJKfQx+GyVoJl6O0RYhA0JY0r7ObY4QU2130j
JOsHN7n5+5qgEoO+8Tx4OoyJl3r6xBxG440NZU9Bgf0F9ZS1bFWngh7dup1dP1V9o7Hm1FnlEzpp
B2ruvLHDd+2xbSjuA7qkl/oC9xy3Lp3gnnjiS+tsvkZg4vcGhujZU8Hbi+YwOwP1HQzNS3NrJlhE
l9IsaYfltDKpU2kj4hMV58W83c9b+h90gDN8DeH70t0X8wAsBgX454Y3rfa6S7oUmTB3JbdBIKZq
uTDTzB1aUNEuqPHSabNUJ4LFdmFgTXkLj9f5Nwl4QL5E8jHnqlHlBkrLxqXRBMSvphvuWNGZxy8t
lcoKJ+cc2xGetW5wYPr3NZQNfxGUKBmFCU7Up+30rCqgoFdZ2xiCldmCWeJekp3KtzUMhKxO9LMy
Dae10mIbdAO3WBdYPxRT+r0qDIV/ASZ6W0whe5x3gqgrZEMJ59qLsgjCDKazRugy9LqK+h7V+u2N
4wuJjx8kX56J81JjRx3ApHxY8q4OWY6g+XEJgozSWyu3Rh5j3v6mLNx8F7m3MHHVvepncuu+cI3Z
aEX8Tz5ENhiZ8xZCp0Dr5+9gZUPOVG7pwq+K1Q9X1Xiu1LjcfhGWiI0rk67xXnPHGbanv4NctilS
rv8Ka/9ROLxHtciNbVAFXPDQRfBZ4FkCa/MB5RUTxGPZIFe+A2pLVWFJG8ZMS6dz1LLyqe86JqXs
R13v06cj8KSlsXo1RbX95PItllNEscQLb4BvcbcLM7LBbRxjxlkbYPEafOdCdLXJyGyvtc6Bg11/
zG7OgutYNX6wE+QTRc/8pnoOv5HiCQBnPDQQURILzjzSif3MqUzGY4ji7sqiJy4B6zGGqlngxvM6
Ti0OO6K1nYpeOdX6XrfbF+JARiqRt7Xw853nwey2Nh0olPR0siiVulQB1YxZWzbr76Zh3Xv7sWPG
TYGEi5dcV3cq5fPO0vBQXeTg3pzcst9LtRxi+4pR7069cCRe7FWBrS5sWOFX6W0t5eKFzijR3J7B
nPquZ+3wtW6dR7y7oHgOFlMdHl0eAXk8cgtaVUJRpkxUX64nrZwxieqCSgTwRJulhCYctwweIu58
GSYMC+zKoeh9B19UgVDxP3C2B4hc5B+geyg3RX8S9c1oahpswkBsGyJgQ8WUowuFRSgNqtsyE4WU
n1WClrU0J80q/Kc5VL84WCMymTW4eEttDFvCBo0B/hvOPhO6V+uwdIXupEaoBscKG5JonxrB5XA7
F/Z8tVL8wjo8VP1hixv6m6L+PHC/3bISTvY9S60OwWs1x18VCLx2EBLraP/lWiNaz773l5Mn5nMS
QDk/9d0j1UwpWZly5zyCY2HhiYRRwIl5AtxkvsXagQqYLbuCwpUGRkanCZ8P7mof3jr733DMg4ev
U01/AStcYqvhbYv6Zx60rXCuAZWGo9wUZARuNVdDck+1ukcWhzC36rTpI8wff+efBClddCf0jjVV
V7igykGwABAMqM5eq4Xq6b6GHBwUlPBwmQAoJejPCv47Av5TFBo0ae+ZTPOnDl4EShQn+4jb250z
Xq9rwIUq8mzDIYxXGprzB7qU+Vi1Rdra2ebCwxub9R6tJ3UbjmMQpHTjXNsy6+WU24jGC+udTeig
homBVpa7MqRpR7LdcFRs9z0gjwfYXpSt9cKp/6JWmKnkAqDOcWkZ7vwbTr6rm1LSYKCRfNTkFvso
/f38HVVyPURrLeD5vzASVR9q+7QOAqui/OHoBTcY2O5iuO8mvKFOHs0IwP99kYJqPlu9dFiXgsTP
HdcsZYSxB8eAZxY/VUx0Ut2iKVUMQ2gbHimqL/5HGmGAHhStX0/SQb4T4lbryvdqCWMEkQLidN0N
JdYe7s0yi82h3Qq+6J/U/PhfB8CwmAGCkbKjziSB6HWxJjwsxw8zcy2a9VAykWcfGH/YqhaeKZyi
iH8ckSLWjmVSc1Cmi5ToyqQDC+3U3ocr0OftZmYoyvsp/6N1xY6v9Tm/rV1GJYxzur1Ief2MSbgc
B2ZsFX+y8sRig3xji/Pwd42xI8qFfUN9dmu/hxlfmLtIpYRE5zapPfI5Ulpo0M4dDGnXaJEcYl74
mEuurIKmiHZnMv+hDQAHd3X9jH9YiHUUlHkzE+F6f126DNfaf91S7NYVHSXqbh73iLgvbZFqKlkf
2kZY/tmHWO349s0ZlmcbOEnexdlvnwD2tkmyLo1YpFGF0pVIPaDb0h6/oEUApDdqc/NrkWykhr8U
yh999YkMcwqe6nKRWO1NrKQvyQKr+ZC3ab9dDkOdaIgPZZq9iidB0SoHD7nPK32un8ej6e5vppS5
9F7u0KkWg5pQMEUdKGhFxTvGia4nQR2IAFV5RqbjxWqM975IJNOVj/59Am9w6VC4YXFeH0+vzgJ+
VmPz/ezxz27Ft30EUXCh6MSQpOLr/P1cXIOSKJL83KlqZHV3JpamiShwvBPm9GoZ3WN4awEbahHi
JHWsJhNUk+inY8ExmMo42xLpDzGl2Ntp9RKk9oagaQdQieZpx8iywKtC6GS4WUSAtLD3FDJpmOXD
RVe9kDM14bHqHBXvCLnmNboyt4l+kdN0pBJ5zWDeK7KwoaVY/FSv3q8vgOia+II2keeKZwgAd1kX
FE9LV3hcf6vwAiKEWdwb/3wxE23i3RAgKo5l8elFli8GpSeCvMC/GEGXUbwLmzzjbxniER/VY1T/
Om/lZDwGNbNUeP5cZn1YfSJAz6F/FWED8qX6qqWt3ORot94O9VWzjSTJPoTkb5ejB0sXhB9M9crG
BgaSuiIzOg93xszsL7PhIv7CEMoWnt2H/md/TA5Lky15Qb1msrQHCUuqscmqCH4A6prwKxhGWcQ+
S7JLNPrYLlRgSYEvT2wwqgYvWmUfakWzu1lUZQdGNooVb2E5zmlSdO2Kg8gzAITYiJwsswp/Qieo
aQKm59Q6VBYMJxnHFJq5MYLir+ZPi1XDwi9+nLRRfs+gz51SXvxXDiQfStLCf2GPjJPPiokzFYef
oC7rrJLmWD6/Z4/z/F6ouLmCbUDQwfoK8+m2XenvBqn9zWAUQ4Ng8Mrc5JgAiDyFXjHvot6w3hME
1gXjI5SuIjFylFHx0ItalgDk7o8DJLkiLtmKTkTnx5lhJFUyhURdceF0L+TdVYpIlWS6UdciCaD4
Q7Tuc5OrTrt01vr1HD1KCUO9Rmb0RalNbTPxF5/4gIRPUDWidn004tn81NjtkFLob+5KjIp0aEbj
BnNBEVO2C/hpKP2iaWbabHj7rWcHxjI6W11A2z3Kclfr+z9jRFgefrRF3J97Wdeh/VSSP+fhGgu5
chnYm4oCg2S6e61Rsr9FHWfgMpuPylR3BFYgr3Ijgm1wXEh9fvyXSEIdOINJbCYB/m+lEW7ygewc
yefz57/Z6+R8N6HUoZK+ihFrofTu2VDDS0zx2a/8nE1hjjzyEOPbvQH9d0drkzXWQta/JxbiS8q5
/BP6cw8Hp2OpUYOdnEa3M+1bAVcI0f4E3kM0qiNEYMuPl4GnS2GE2XLM0BoeqPear4VRy6e7AwO+
rgTXdFEKFXlEgD8Sz7U4tocbhpIVjd63M3vB+gGpCiIZ65TGI+Pybob4c9Pb5xgzq7CQBLDcgjwN
tgftU3Wig7d8Nw/zi15KSFGdsoFfD1G+Il8hXp+sYP+Afr1s70OJyhBZt8IEeQKu5PmwjV7F8JAT
9MWydVh4fUQ963MFtAZOwqBfQYXxQvTfFAxa6/Pdadq0rip4fgSB/+e61vmXQ7CbiJhxDvB1Sc5u
fKorktaktQa9eDFFDHSVWvQBzIuuZ2A57BQN94ZxpBFBpJmRs93B9i3Qsm9+Je6mJfA0rcJi0MdZ
QOnE3d5m7VJVHl3jVg4Dy76zhQaC51qjOEOzHOgO4N79gGog0SmHP+mUU6AYSIDGlLMHemo2lAK6
4TpS8EFVFL7Qf8/swtL+4bbiLzsn7rttixiCWAinvS7bfUBdDOMonqN/CzWtACHNC1F0u6lRSQly
ZhcUxgO0YWqXV2MNZu2bPpwoD4TrS/XcHAZ365JCfaF5JyZefGd/wBwx40CMXPzP9r/YweTmKbwV
G7XO7zvBx0dwc5mPtH9w6RHx0O9yCBQlBK+eZ2oftI2E/s3kHf0OlaXwUyn/VCYKFcfkzuDodSGx
z5qFYruALLFgJXxbJ4CGsR02TD7qIVeG+7V2LUPaaUOxQmzYYSECkhr0fjoK4xXmYJ/y3GLpHMCH
ZRyeSkcCnSOwVVffxEdffD06l/w3yF/bKxb/jxhG9c4CLPlUkBBxmfk2PrVsbb8ELlZMHI0UKKV8
lD0sWsbDxCfAn4XHDq0KYbRAiEqIfREBzpJeh6eH6G04h/a1Cyi+vRv0chDDnB4T23hLvBpPDJ6L
kqGkg3nIxQNh0iqN2Lxu01rnXJuxa0OSP6T+vFB9NAhjsDJQfemBiRJ10oRNlQu28nDz8N7Ekyqx
2UlqLNysHPbNO1ut/sjjopVU96yi+t3DR6zznxm4T1y60dYVXDaY2V402a8OzgXMiOeBj4Fcb4yU
Za6tQxSKz9Oe7bhybGDekuQqoG2Ql+hYANxeAZatdiDI2ZdHFRJ6TOEeaM7mKOuritftmZqAtP9r
perOyxdQHtP+D65QQFIFnAu3yrdajouqSmPgixrY2Bq7/fIGAjj2CoCa1Zi2hyxLWsUmAyfQvXdC
RC6Qfgf7J8ekJACNktEckGIiLXlZwWCWzmeKGV+bcuGh+87QrlPIuE0PwYmR7NH/akqGd1n645/D
9Y/rbrkIlSK8OzCPnwzvKWpvhxsxdf1bMsYnsMGwshP8Q3zHwl0wHo83XsbILvyU6q4X6PzC2SfS
liV2CB7B1LltoPtpW4wWvGmTl7gei1aINJzuf9Ut7/d7rm8SjRGU6ACcK3DGQaf/jaOCCmqJuxGC
+t9qzvZ4fORoINXZksmD8IWRoykQJvYza+wQZkAQapyC3GqjoQTRIW8kmI4CwSN2Znt0XDEfI/Yc
E4KLg+kG1F/dGEatajnqHHiNQIMu6C5ymibF7F/R0v5zIgpSw6TUMKN82x3GRrgduIXFnpVZI16n
uXNKV3GXVLalv/GbphO3i+7z0h/P2HpGHfR/L6OYhbziKh8vVr291FQblKIt5MWkvOnFew+aXSEm
jTMZTN4vL8miFg/0N2QmCKMXJnmK66o/0Xg5lxh4oi15HKVaHjgEm5cdI3szzQmTfF4KV9ygXH/4
GPueq3vyyN7E/1s9ulKc+GjrqjVeGBgbTuSuSTEQkaiccP/iKc7wwFqoJ11ZRLqGl+1fbnsb7Alm
LYDxuLqhx+DOxCUilc0XKvxuWhQTbVbRHvjMnYICBrK6cgTgBX7YUiE+8teuegF54Lrbt/6xFfQy
k5KyhKhvIfFHTRFAclL543qKfE8S5CmmO+VrVbmzivD6bVXvB/qRoCby25MWJepR4PnliDqJkxni
x0j511Rg/wT0crTIylA8Kh8vJbOpknkX8566wg9+Xd2A6J1Nd0BhWmV0URggQvNuRT/3Of4ImGxj
oMKbmolCYNnmcHzAG3WSeaO8Yqjy+tcgmYckTwY5+6dp0gpe6+pbTyoSE5KQ0xGsYkY7owMlbGQ+
95WPn1hQY/JAc9iS7yM4H1/LGUQTs2U2KSQgiXYtnjnGCTTa4yaD98sjvnNjm8TrtcCwTrdi2zkQ
L8bTZG4XUsWS44IgLL3qSCEB0ygYOv5Se0xfHr6gXydRdypwd8HZP3/jB6kFhWBZ+Dn/m+4EqI9Z
PUf/I4TlI0MbN935s1RQpd8Sd80gnMru/LzD50QVDpgegzkqU9mxOFMsX2oSDLhUxaTYxgO+xn0C
MOPvwvXgqMK2ideEeTYkOIySRsiSfltAhw9MwU2QiYbzoT7tq2IVU4FINViiny6IHGGAZxntPJFm
q2l+Wnx7QOTqaTtWO3UmoM7vLWJf04dWNBmePHbj2q2DCYKOPJuGKKVothzv6/PIxbf+I9phXLS5
8Ii169ubgZz2AOaINxvnMy8xwKI5vROzbrwrMIrrCKsxyPl6O1MKylz9CDFH0MF/nXklUXIINS/a
XV5/tUmLPpFOi19aMEeh9zGH2w0+ghQ8D2iNM6SY8fkc0DFxw5ImxMzWMV+gOeJBLx4BWtK6Tsd+
VaDWu/NxJO57r4fvfbIfA89wcoFyVl4W7u2M5qYTVQ+eA5qM6dT9jrOfLXUyngnKraJQ7nEP+UBC
nNeMC/uohqXQFpCRrolx9vWO56Dq83KhojR1BM5sv6/DbgFDQ/ZWiNTqfsqPmAD0syh2ThrAtJOE
hPf1/4DuBpAxlgNJ05UyYyM/17pmYy4MEs0cyOwQNgKd7safF9L8YJ/RE/JE1j5qNUl4BeunDsRw
I8FllqZGSc5jQVW/TGTQm5+08f2Sj87h5hVw9d3W5gnmAT/tQSegoka1vgS49GEAxF9Rosc/fcda
QCEPDp9abapx9ySfUIC+u68ILcT4oUAcc6rFx0sGoTdHV20OYyiYvCwy9fc10m33UyPdVeB1W3Ee
Fr59YLXGMZpgLqLsNDfq6q1bgHjc983V095jfOTQinZGLQTPkgE+2sNck8JKKoB5XS0RukcnFk7d
EDP67VsYyor2N/Vg6E5n21wPLuFPsgopgorIELZJ87nvZSmZMRqrPyaDFGEKoO4dRGeUHATQB+Lc
SjcpSR0ABzsX6zemWH2m4JK/oL30j9RwxVD83GjrbslI2ML34xpVv1fA9M8sEN5p3d0muksZS1IX
qVVgzku5u+SBgpvMthk4FF83OrO1zlrs5V6//IeXGzzNQj56gcWEhrHLRXEfszjAwLXcL22NrFAc
rJoPeuLev2HQHwezhkNclRECWkjadu+PEQF9f9UDUUuV9CXK+WEX9hhkKB9gVxwfaPlz3HmNflz9
EXU8Kl07+3xcVhUJOpzOPlclsEqP7SoPY6eFqgf0O/uUnXva39BingVlCVNGN9ObLLgRBRf7yKUV
keI0Yzqd6B03KBTclm2kMgE1feQcfU6y27MKbGMnkxG51kkSFTTyebW4setIEiFh/TgYOsp+QdfZ
g0GooUmY3FyoUEMhLrswC1whsArRYU280uRNURpo3hD4elbxMc97KOAnnn1caT3IR+FaRGoqtRlM
cXVFOxMTO9cfWEOJrLi264ifh5/D4gU8qHvP3v3jusW4o09M231fqrTjrCom81D3Em4Oe9rz+0Dj
C2bD9l9cztCSfQM8ZtVSaBK4mvMpiucvFfOZBTGH7z3xzfbC2yrBiApgebXaJ5Ok2X72cqYDXNrg
PsFDlJsEyFFp9xYyEeBxeQPT//cFYR+ZVxTyvEwZr14srUpz855YRjLUbzB6cviGE+w/J4dR9VZz
uLHBnUJpJ9iF7lqCWEvXddDOGzGz0oz0iHT2K2Y7JeIecuDJgpN8LIMSQnRQmt/5K8mfOmq/7TZq
n65u4XiBePZe9jJKS5lEnjU2lo7RI9jb/ZV2BCufEm00jrPxTu9XGJjnW5ey64jP14annf3LGxUu
4toCk7qKa4n2LsXj27QJlLIJzLaF3O+ijVdnEAmgNI8u2n22QaYGsIJI9LrmaCdAJaXX5VT5lXCV
vJE7fMJhd0LdUTT9JOMkYp1+/BnKnRRIKcEn8xL21Jy9q9h88YjFxdHpVylQYqVtEjA2reVgRT8D
4EH1sC1wVw2GFkD52KzbHL7MgIV79TC+5d/Ws27TW1FY5WNb1xIOhxjq8MUTokVFA5heG4n/2Xjb
YNhAm8YypVNE5NtwUNNiUrK0rsOPIFX2BFsUIamRTh29PEdYwqfPq9a2FvsevUCZbqdubXy7Z0PW
/nUhpx65V6IZ1eVCWR7SXe3JzUWmy8Rh7bKLcIsjVlPCr451SrPOjpq3N9wJfBB8DGSNcF/Hlgot
pSBqYhAb7FhUSaf0HxGlhgxxra3Li4Sf+DSxeuunmLX1dzTVCDtCmuZkgpeGsYPaEbjOf/eBK900
A2Mn3K5kSInXypE7JpJNGCZ9ekDP+7Wo6E5m3ONdQ75QXdCDDLVmfXOtqK1qJAd9IHpZnGWEcR0K
5xCoFeSwGI4sdVS+iRKCClSl+gjv1kIQ4SpXBaQXDaf/KEjpzuo8m6UnZ2C6ivWQrmwSpqd5Rvnh
8bNf53i0NzHxVwXyGAWU8b8/LwuKUA7NHQJn1O9YX+iSvOSA9cUC5MTL7KrrhOPYk3pgFNxIfki6
86t2tMtbnVKR0vHAJBn4rLszAMJlY/igDILjmdFZKhtTqdJBgCV8IU6g3F79hCYzq5pyeAxOawwt
udtZKBRFjZXasxP/KCf3/xRpsSD+kvxDcFfWfV/RqjTb8ZRUNWxyTclhwOvEYo52BFNlu3x5j564
xqDpmMjwtxrR1b83qakS8PhECKt5flNzWzhuyJI0O2MEvkK6qBTE0w8phjGwmpRj92sAhR3CkEW+
lCxlnnhnCsBaCTC6aDAbz8R0HmYRes/PLSQ0EtWIhOwbScMjmy2zsECPl1rYQZ3vtWCb0r66NgRg
r9v8o5JiugdMdQLccS6qVFY33whyAZ3QNJwd73luM4NZ9jeODC5AUpugAbHxqa+mpZ6CbyYuUhzz
hQREUr8eU08Twkd0QgoXeQhb/DYgENwxYJgm6caMRkgu8d7BlZJPmCdNnxSv4274QNc2rTXy1kTw
2cvbYn7Vx+XLeMYjK5i5zXRJbzQqrTqpHKZIoj0kvaJJT2lZmUAWiXJGmW4hfFBH7kN9tNp6r56e
X4YQ73SEGigcuKlDE3R95U4WFRJgQhN0ufwSgY5nHkMKWDL9tBTbo7pA+OcVLw+xCyjxCBqNnlzy
1SW5slwb0lBt4iyg4dAc2JQBnxIBcn+Vxy+BFZNLsaEGJpu/GalG6LKtElZai8v0JYEfDTgl97MF
3mabT716cSri6aJkANjPyTZC0fqziZU6t5/PisqqSaNjVM0KBT1iaPr/N1BdDy8OJI0LNbJH/KnF
tqM0EP9DEyP/KxD6158MSLSTm+pO9ILC8jatnhOF+rCWvHZ2Afz4/8gCPklibB53yvwzNVhy8ECQ
wagTlL0/WzJNnu2aAMd2C5aAvGKQ/fiPBhzFWVWBSg7xVLSsq1jedcak5H4eEju19fojHuZPBQDT
rbqeRTOnfBIP70Zaca8ZuOUghpEEWUuPApABaeb4vewdu5nbA20BG9+ZUAIlSkljK1OETeymDcqf
A1GjWalB1CyAXlLAxJBxXipaYQQGMrhzB6R6PUx8IYTsJUrwrn6Z2xjzoVNuACIA4S+IrpX+0k4z
sFH+N3ahz39YH4vF6KaiR8jotFEIIxaukKFIz+tRPvnVjKIytFVNlr+LOAa/vS/T6sEELuHDl3Jz
vTJrYOXeY2/WNx5ZU+snIl844tAvZi+6aXk9sao0cyzCf9ocpQL+vzWvJnLmQUrkGpf9Vfl4SvFW
hcVdhiKAUlEwMhVSIv33LhzKn8tiXdMjdKZWMxABajY6DAbyYxSlojb44Te5YeXamL9VTbkOTJ/Z
qJPKhyeK6Ok7QKBUwxehY5PTatcgloiwjrQHcx3HpXR1y+mnb8bl7Cie22ZR9rL3RqHT7usDVIZb
x/Fk1JdIgIwg2o0MtGVWetkJpTsQRXkdTiKeIUOy8DpQm2S5T40X5g6ToNaMN2cqC0Ny8m7XD/Ii
xBL3Y5tuHA8M/GsCfKBz+jXFk5DRPDXF4QVkSoi4F9gZUprFdBzt0FrLSU8orDfm+UWjoKIjKLA1
KAR2hAXMOnhvTI/FXa7x/OaQ6f98yKIVjhM/6Qx/kwePnQcCPB5Iu9XAaavs7T1Xro41MeGQbcyY
WWNazQMXRi5BByC9Z8RJm2ybISm3tWwwdR+g9X/5PT0bijOkZQTiRlGJEkNiFlEKhg1yVfzmgpw3
Tbd3g9MAXeVwykxS+aAasI4oH2/CPBIbYYHZWG1DX6YpNqo6wBMhbuEtWG86MnjqPGzyg8O+Zs2Y
ePjwzuBWXPTI3p5jQRkarhpqMeyorkppIaBKEIADPk3D1UH8spUliqqDf4IKYunp2Ejk8PF2iMCl
FrTGa2jGo6r61VHHtW3jXR84Kb3miGLqdszqmgFAeevZ3Za67QEzxk/lLg7QZJmaqRP8JBHI+w+a
VN6jqxNQXpvFUIXCl6vNE7loaojOgSNfN9eIIpsB29FNBF14Vhw+Z1FlHCl1joCngRVcLJcyY2w/
ABjcq29Qe0dHFxa4uZM65PamYXnUBTIC5yNBE3CYHzCRhUI/LBKQLCatNZiAt2bXZQJLC8DEM4UQ
QQKbuPgMVWWc0xeFP90TOqsQ2xPZGLOY8ICImhoSRwJZgvENNK12aoUsQ66MnaLI2Jt2Ws9zpzJq
fMvqYJKPrv/u0M/h1MBSF446t4TChMuSNxLbd/N7uvpXuy2QsdYXCNi52SdYxerV2wSY1EhChPt3
O8JgqTZEE9z4xI87kRtN0OhAnTvuGaU9fgHxKhe4i0MFrnhVdyxqGsDIRIGo4Maw3GuBAcihIk9z
cIrKxYhzy0n2pxogx78++zfFReAJ2nTBb9swT+nQBgX5KKHzWvzQNwuBOwnU+8fJLP30UV4n8LO5
HOUngHrXYPbRbu+VQ77iSF5gmQOVDFERvMCuxm9u4cY8cn4uYeJyfJhsb7sJXl0eCDGfgNK42C7K
wpJrdzPR+4RGB/nom+m2aIo/2O3MfQFFYOUhuvC0gwwCBbTi/vMitPatp073YrQk6HPf4Nv+Vz3s
QhJFSfHlEPfvWXFWCQj0yaA4JJYeDaF0hkwvE6XdkBooUYXxE8aQJUTYKUUX+8k/+ymJwriD9qf/
mu3/j/vn1VNE7mSdArTDKCoiIJkDy/3xD8yxlGJ5KJ4fSE3SgPP1Tc16VXUQHg4G0MudoYPwOcGO
V11ARmA6AjLbpF9jxZqzzCcx6SW6sXjoNQPMMWKJv6QxYRoz2+CZtUAatJWR02l0pj01/odkF1Tw
+Tw7PBg/iwSMxdXpxPBlOQjcxKAs9HWBMO+uFkq3u2sqXSPVHk+mBtJ0w7c0WMVK61QSl8/yghvs
HklcObOYI1RKEZQ1rV52Jkykryvr+39oDVcHTbWqTJu9nITKE8KAD65NVzQ5j0o2juHZ+328ioLf
zAk8Yur2otZqKu5Y4OWbyOJnW6ok0aHLdCyNqvs61a8WVli2Yc6DZgPLZZl+NWFlYjlRrujuFgyO
+u4FbLATsrLtUZn3tKyrH0TNcl20ZPBVAfM5DOEp/jf7qGjT93LikwzoLUVLWfHbyzGLXZCdeLtJ
Vl33s7nUeTDujAok5ou3HvlNw+V4wXXGAaWiMMbOz70B3UXP1Buyz/Dj1IwcLS2dMesBXR6vjmrr
goDa6Jcn4NOCzcjPw/+tQPRlhx2ecntOVikMaRL031HyiR10uyEla2VHqgBcX2WChvFHBxOta1uT
GMAgYEtoELJZLNRfJC0SGkmGVpJGBGv+CsXSnbbsCDJn4Jj8MC1opkE/HXu7bvMBLmbmb+RAhKWa
mUc41+wz3TV2w9d8EUA4xvNu4ojDn1ERiMRpJdf1QfDsvEPzVcjol+g6Jc1Gp8/ihw/ys/DjF5f0
seIOPE0SHWaZ8We+kIx6QhNy6AmjGe45okUTjANs7N1M+BIAIP8Mo/JsizeRQ2fV8HGsNtFLJZ2Y
mpf0O5S1Mt+8GubKaLalMd42IEoZbtOnkd49fVJqGEnb1E3lzDGKOlrOKukKpjDIAP87XrpmfPi+
i3a7W3hrUNbpj8ymcxdrTGMig1Py4V2cWAT+9bhkFp2sSOWPqJCVzuzbrtsalNjpEsQXw8NL+dAu
TI2dEyxbV4IMku4R2UmBKBhsA8O1YP8zL4hJEG+KFzFV8L34L3SRc9hB3u34tcNdNZzTd+LQ0wts
NhtfHjR7wbhlMfxv6c0+WWYSpe1t5ng+jksdxr6YzbTqLVLPym8CMdngtJhIJoiynF+Rh8+aZTpN
6vP/D75BSZ41VxiFJ/fXKKEWVjsWlhCSaDxsMB8+7Bi8eOY7LME2HQIgxUGblvA48DR4Y/07FILs
TSzPWoTlc/jZIWH3PDaijwtGCpBn67mpU+uwovPYlki1gcvEIQe72VusSsPBejdOkT4guE85lhDI
jlsA2MVI+bnZWC60UhBfcuj6nFI1oVrlHL7bQoqZgvKs6RzvVXzjaFo3GUyqOfErfQQKQlkebvYm
g+E/BlPkzch5sGub4Kq3UNiGxHmCTdB0EXgcwLYNqEvJR0ZdxH8H70fSqJJnLRHDnsqwpvw/unY2
oBYWFDFHp4gjxlXbB331bAgwrpNfefEpvXYRgrtdWKM/VNsM8bdnq8Bb6Y1LJ02x+NVKYDxt3gM5
WZeey4dkVf0fg4TQ7g47Ek+YNQx3sYsKXEEswkWxsRIZnVVECDg0KV8navMzepUzlrKZcxZL/ZmG
W4JD5fAN5aYo/ac4VRUGbnagWvqKSDY9oXYspVg5hlATDhujGAH0UCYDHkV5XOQs7MefkyEXk1bt
YYOh4EKRAEkaCPMnqDwvxeOhmH0vdCDiCA7m9+reMvogHSBBaM3VR7j0pGic+D0pjePAi3k3/Okx
iB3MYsjy2yFeKSh+e9q2Xiu40GNEwFtfSZtekeFH7b0ioA7ihnrsNCWLn8cx3vzkyXsNauPVk/os
rBQNwQtA8ZiQKnLe0+I0BGsKRN2etBRQkyD+ziqU5iHI0bu7BDuoarIJuJbA6X2MNK9CgWuGE+4E
zfPiLUpJJfRHjCLygr7m4Q0vla/ZFLkRkAh1hXPM/apaqDJ77vHUaQoe+Fy61rR9u1PeLtBdmBe4
YdY/rmB/eKTU3p3v/6zRx2OhgSWuV17vDeSSMErH5Ibchkb1kkQXmz5yiOiIDFnNDNVTT50+WuPO
MKqZw7nu1OrHynuP9y7jQHddiFU37UQgbsw9FJbG8PGBQbB/5YFCPEOa/BhCLvlF8HPKNnf50MXx
GwPfyPULfXI6CvPNewU3PU97valKfkIJaJm5Hfn4WSMXHNxc79kolmfsZxZqDuQ+uVBTNjRCV7ow
za3xbdDHKTPxulyM3IODKULf5vRSgmnreVT03MZZ5K41EC3X9OosVWQYdq7SnzayyTiGW0Q+1z8f
881qBIMqiei/AXPWwG6NbUTPgZ+1e59o5Mz8YwEGkiwULNsScV4oLCPXO9DKGUsrpPoA/6WAxKRY
mLAUl000sn5rbO0ibZIZSLyqOWxU0m9sn6sROTqAofHwHIC+nh6eGVbr1ES1+2ZDdr65vjK0D262
zNts4tSHEdMUSQnFkvKeZhX/v406Lj4hQO7pi87HZc3br1vXcfGsOqsnPN9LnJFB4h+p4bQxOY/p
+rtZUpxm4aDigWgpguiEeVFLF9QNVElh2pQkvS9vu2C5QXa7EFn3+xO7hwOuqteXFGE8SCm+K/15
XrwRCiWNcGOrjQhR79zu5mt6KbgRpJ6mHUTf6xp93R1msrFiqbaV0CWhirG2Fybc+8dsLtE/A0jw
NJbcIT5l0ub2gdRABPjWUcH/9hSddROBQzQAdgJgfH4t3v80fe1XxhKkauT78dEoEBCdE4HcnpqT
jy0pzru7Z1goLty6M0vtkr5Nwly/Ck9bNfPnPpj4npI2JtyBBFEMLY+k4lJxFSHhNSpHdoKrr3+f
dqsexQPTlWZsF6L1JUhQTKeKoVTkRzbM9pvgfLvOTbDpOmGGK+u0wYr+STxJvbkZu/pAt79A4WUR
dXsagk+Va4PSgKlRk2g8TdPqMCJY174qrNVHqNz4jiNoki3EepAUC0CSfce/wmG5tZ6USC+487Bl
BLQ8ymXm8SNFQBtEWxy0GElnLF6GglBfb9IBSkYvWt8uAP8L1QluwcyLA7q2FZzj8qapSUnHuy2b
X/FU4DXBPpjivi+BkEdwJyyycfsrZAke5SkiuXrDz7rUErcW6SPdsEYIDgsNlVyigYYpXovHpK1u
Xj5/P/J0MRENIuBvoLeWlXEXvDv0snTe7M1R1iJBXVhvwVWxNsLZCJs9grQ4V5EdvSbYuf898U2Y
UlAj/fPpu/ETDp5ckx1UdlRJvh5/dRf1rsBQd7Wy/UALlSbmKZJ10q/CDRi/ule1Y2QrbwrQPmTT
bBEU84GEd0wwROC2q2yAcrqlrY0dDXX2dNY8BWjEJKxlWJnEkx4AgqAYY8yhxGsWp31V/u4mD96u
GwoOZR52Bu/gt3K+aqZodfTH+KtfSperHENbUizs2f6OLzbnxlJ6CuxyjvR7aOME4yqcKpjEAKFs
OqGtCuFCga2rCeV4+xc33iiUdZql0euPW+yWkZRnzyvs3BX+PR/yR93Y01GlOS84JFh5q3LWeKrq
X3/rOZP3vFEOT1/+TM/x8e3I3efBLSGDw63KKsW15l6b5J61OGXsMekIulCxG6T28P4ud7WbqFPz
vlbsuLIW4+oHmKUvu9xFbmT5nGz4oIcBkRoTJzQ8LQO3jrd19zVxpZt73QQ7MtXySFO6Lbd9qcM1
NwdwgWeYXtS3WMqasqKSieXkxrfscrjcG5fxWPqth77hvcmOSxOXu3+TJT8BXK350YSaFVs54mrR
q4qcBd1AMl582yoN8VwvgUdano69r+p5TTQ4mHG7cU+Cw8KDBj2tDyd2nTMORuBoyQX9eubbvOuB
34Z5o2Lk3ouL0KTEBp8WVA8V3XvJURJZt1KKL+CFfpTWLYFG2njLZn8UJtnAzH4eGjnXmO2gfcew
/U2+BaD51OIjC1bIcLpNZR2OUy1yTqWsSMxk8KIdcEjFvi9nIeniYCzlhjBm5mGR28zWGsO8kUYo
AjoWW9JYJg3O0BtSs1li4S96y8NesUiruuqyT648E/4vY3kG5C2pL6eri7PoE6LiqdSrdi1HRxB6
ugXlmcWl0/H1vL95LDlujQdhdrI3N8Tbm5k+SfBXvGflAgkYKzzlwZQzbC82i/tYgnn4WmymtmTB
e24bSE/06grr9U2BtMcib0lTTk77tTR72pHxXJ1aIOATsYgj3StAWR7NnAQzANLJ9paVufaKpD3t
9v9CjrxszclKsK8rQHVtiEB7bbqOPW3R2HuVeh5BW3TAP4+6Pt7EGqb11j5KuTXPceiGi+tmsNxS
BC2q4lLa4w/1I693ESX89Rf+fVUtgdhhxYANB1g1bHVpV4NPUG5j4rhmyYYuVxnY3nYUlsF21C36
w3emTlErzz0jamQKTcIZ3kV49BUPXMIhXHzpuHiK6TEYRhxNuQtMNE4+g2vpmnQxWHS1/t8elAO7
t9pUFJWNHU7DmJc7TQTI/DXtHYtkavS4QVMYg+ESJH3KnCE85VsallDVUNQufst/pMnFsmaw/uF8
uiovTqJ4MjbvAg09bqmnVKinAl8iCQUqjLpwALwtSG5UYj+As1DwhQXZJOzQlPMCzXr0KfCq7Qt5
r87OyjjKgWqXGvkm6uh3q7b2MOzuosM/3KYudXdpZhGtRF+6z0gdAr0L/hHfmG2gxWDHsFuxX6c8
ZtcfnHs6zYv0kC60vt1FxyDlg+//lYlmcieye3JNi9Kv7N+3NzRZ66tznDiT5PVvH0svSZe10m/T
GwTf05PVy6KfG9tPOnDpQtw2ASCF8Q7D3J0XnGLQ0UczCeqaSzt8eJ0uUq0OscstfRMRC+ubg6bZ
1gMYT0W9BZdLY4qubCevE1ZUwjXmTeX5auS0l17z6UIugy/A/10eeJlLSyT4pb6MMApSlyy7OaPm
P8mIV585AmMhg0HbxFy/K208dSnusID+LbS8qVw/OrVBwP36YWWd5d2jVPPP5dI+MLJfgtcFWR+7
BBMQwWDXSER2abW5AYDeNCDf5I8jZCQuxq89OC5a689t8yMonJQFAhANTfeNZJ9hRQKvfH9BLLVf
Mah5H9RwWFcDtZ2Mb9wEJ09CXls/YR3zzfoMxse8OdUJQGsblEZEDXGZTd3slRVJ2t1Tis7oZ5Qn
/+l+vw/QP0PiqWPQGP4/X/P5Qlsn/6d7K7ArFpmqLsHd3ULc22QMyhUhxnSUKyx2LlCy4CsjNP7s
i1A2KWxEUayBeeiyXOgnIGTZ3NqkeB2Ebzp0ktKUBIW+ckrr5S0uoVdy317+FnFU+pLq0BieUVjl
mGAz4BVWqXlMyivAQJ/+taZSDfeVyN9tkQ6BP8uqMm1c9Jxm8wgArjA3EJeLshrvEfy0pmvi43Qy
d0Kd8FKh2KeeSU1g8pxCfnN6Kn2hZGQ0Ch3cTs582kVh//mwKavclry0M8MbLuWSWieI0QqrM4fj
T53gF6tsminljPfxOFIXXg0byU6on22Nx7ARr8EiStcS6Ru+B8+SEwA4oB99+f669iaVw7Az9UAU
2n1/Cv2BuNHUr5WUHhZAQowDCGqAa+nHqgW2oIFItwQLJeCy/IP8L5Ial7bze1TJ4ZXIT1F79PGo
wh0lviMIPW/iPb035gRoaBcGjakoNNfAkfdF16adEPrNcxmQ0M+tlzRhB6nDpq1hBB+vWmpcqJYX
iF/PnpPX2RI8LdcuaWs/sNdEETVUx9r6Ps9xEQs2qN5d3GlC7RmOltSYcqAwVAWl9oKT4lzNWSBX
DOceN4l8qRipmECAUpfKO+XPksjjW2JG4Roa5Ui8m89PiXDCYMl7jvvVQ+JtwmsnLOeiwYpDHAJP
EHQWvjihCC8mzl4GLyR+sQ/J+zgkqhFdMKtfbwp8sdubdJ4NEwteMyoaPgIR2AwAKn5INZfxMYxQ
PlVYWfDECixC+nIoeFH5I3dEDfrJhfpaJhzSAyNk5/SRbh3RwDK1Jbe8GLKSKMvEm4XYzbWzfu94
vin7Z0/sj1NIodTJfrTBfqY3vb/KACwR8PkrYvDy8+ZsvmMOgddarGv2Ac4cN+FRFi9MUMv3v6In
LgWJKpFLYoIySVScsHOPJFF8ic20rNZlKxidK1pMGcwx0+dflo5gmTZ9o3TR4fj9DvWusogxnJF+
ptpaZKHO/mLYGdVQpTpwX4UHQnul3dyzPjFpfxM5btEXOJhBkm70FK9GEWu4uBuSPRCHe7i7Y2hn
GOZRJJsS1Ml3foOwpIALwI6fIqxNfunXxsxRJ14X4fvyBWxUbMiZCrc53aJkH++dIoJZ9NAVuY4/
KOjFeKHCurH/d7+jB8/YvrKeSoz/kHe9hIL52QrD+p/Ik1+8Y2pQWCc9XqM+ViLedOL+E+cSKDfe
cLudKq9tC3Khijbtb9miJtkEitAZVjA2vyT+Rc91/hffekS1sbE9iUNu6YglwIgrJsDNd4nS7Xuv
PnlXMN37M6FJi1nUPtC/ITGQCWx+W2UNrswg3Sb7+RVBVkoDT6A9DX3dGofTg2dqa8XLa1ycdcQy
FMA+lX+YSF4Pwyx5oqoenjg5uIp2oxmdK6O3pqq8XwsXZzHHTtQSx0BGsvMe5zKx5umedMyGiRk8
YvC3OxWYejyDmVpqtr92lwMoPAZkV25Fe0Nlkv2hTus3w96slGaTzTbrW6Fuh80coSMW8gKEry3E
ftclH91HDahxBddSKEdz68nUKk918ZTLXnD7sHTYlkPM/8sVA29TiK09Hf/+z9cbRTfmpKZg6L5t
tilArlAkbo06/HKN+w47fyAH3uA1/SdSVY9pq3n8T0OoBTkDuFDzrjLPkUD8xxQTkeB5WyRi+ylK
X54PRueMh3GChXYORze4MOy55MQe6nUakqb/GdcL6ujf4MYazRmivPLGjbAuoaoaMPT3dv7pjzf9
TV57s4jgmpPYtnAHMPjOxqANTrtYQP3waZ1sqpspGOObUP/cqMz44MmIdN/tFWnLADY1E0VAHOVJ
g58JkIvlPrjFrzbo7oGeL9Q/4x/o9ffdcSJ7NhZnT3S6zuD7tgoxPItn3FI7Hs44et7LGA2zHhuV
NHMOSTVPp9L16HbeFyi/Oc40Sk07WnR2kGSPuetdlu1J1eUtQYlgT057OavasYJGgQNdWMJSppAE
baSaBeih+95pldhWJNnZSs1VoOqUwaNa7tlzxTmFIh422Rhc/Y9iT8mWjDsIS52TprDkiZf0h9cR
XwqgEgzhJSBVmflDVpMhPNA5GpRM9sk4l77obL+g2MSTNOnQO9hh9gisfMh0y1pS8S4IO2i38bx4
pG3/VCWyqkWBrtSFxpHhlCPFeOt5WverG5puSegWlReTT/IClw4PHGxU9hiWqgZFNsbjBNb/Jqxf
bXxZoy1xgmljiIOdI7M9DnK0lVFOzxf+eyc/Ct0K3WvpDNEpcJbK+bX1VUYrSmeBipd7NOCs81mc
bZbqd1CXuQt0gzwQ2svHJAK8cs1VxRQ/caXR1pvO5gXwom0DE+LzKEDMQsZeZl9HulqvDLWRB1q2
lpUA/p3RZ+QdXqke5HN5hsuPBLy6qHQOdHCIDh+foa0oVuP3bdDS1l9LmfXBdcCmO18QGSPtN1Ue
vqrIuwqHkWiMvRx+0nN7oJ1f0pn8C7j3XrEYsNo9vi4oaTSo5JuD0mJ5OY/IT5+h9a0iQHATpTmO
odCJvK4LpPyByC6i9V6e7e3T3d/5Te+diBlxbjYaj9/EUmyn/vx3zWKkHQEVOSXBHhC/huVo9nS+
+RU+mK7rGSA8CyT+6Wk4qWqP8xTxv1pnblV4hv7ok2qzmR0+4OT+Kw6BGoxsirVf2044ibqgkl7b
NyZYeWs5veorxXoUfe2nllTh+FxcPxZTBK/6v8IKIRAcEQUhB28OPcKAWZdjptn6pM4inanEKbQb
HVQ4uviRh5NGFh91VlE6p5bQ5opHfCAuIxJ6XCD8/2gGfW6GV6aG+pNAQ6zZBbNLwlw0looELj02
2ajcrqW+LySFYX2IJT8CWOl1ZEcXnKi9gWYgR+EFaRSDoXBitcuuVwoRVvo2RZ/vIcO/AxgW9O4z
xnhj14PBobfzWLME3jaYLsJK+RzZwlZlQsupQC6ehz579g82pjcypIbFtbRTqmZkbhM7jiL+aNhz
HPMs5SU16lMvMJNcDmYo78Y3mYfy+U02lgDrDMNQn6TE13gQ3tiWgtZDgpvyK0InJAd94O8LSztZ
3a992ti83ZJ4DT1dJgbgiGzQHoXerACQ9GmaqZMTvdVlEVA+g8Uq875i3nia0ojdLaEae9bLgRaC
AksdCEv/bsUEyL2v9txr7WyI6L0LANaWkC969g8USbohy67t63XADMV1RRFmuoHIQb/6aTU893b5
pOVYLqANuOgGEcrSJSNk6SJjSdVGXJ8/mUPRs/QukW5/ostzVklz8Un2ZzEADG/9h7R73ZLwFMq/
IiUwzOMOK2kGVkLJwQDJsAmgMrxh+exHKM5dzkwhnm/M2Xi7sEbrEYPxnDMRvHDhxSLNAB4pxVIc
iL41EHNONnMcMv9+AZq5mLSGdMeRjxtUNvYIx8bpMrT3a5PehV0mjog/FEINUocQHE4t33Xp5zBr
q2Ws2rubKn+6se6V1VFdaSQ15FcAiln4tuQSO4IZ0uhzo+Drc5OibNDAa+lztQSdyOmanhT/iHja
DdKQHXvNvV6OJ30Yhy7m8BjfkChF7A9ohQCn9sabdUyyHBzz2fG9aNSLg1va5R5V5qYoZM8inmK4
d9zven/5pgizpUBUpVIBrmpF7HE9ssazdYNXgcNLZCa6RgzM0LyH+pUV61jYOKiDujLYJja/BVe0
dYaRYOIi42EPG6AK693rPkzeb2A1lgJtaMpKMsp+dNQaEJsUy/jJCxTSiX6uLMKMT+7yZzd9YipO
QKkQCr2wXJRAkTxUXA+BMqVIVlZJU1gSLgIavIYyG/L31SuX9OsfRDGG4VJCX7ib4VnnTdKJg/kL
o7yKLNrUBgKyW7DN/R8wfI5QosIeudrYbzZwsP9GEpYbTo6iDwijt3qGY0+iWjWnQ6P57EnASerY
sQ0f/0STK9Fp1E2tuYwRTvM0LhmmjZ2R6m53La1LH8E0wdJayKHGcEvq4Ebr0voBlypOk+G0RCHN
Ci5VCOfn2nleoKGTZ/VRYixElgu5Cw/iv2RWj79GoPP/kIKcZaDrUK25kf96RUoYszxkFx92HjnP
Mlv3sJFUdRHdifdW/dO0fTg/FQLsRSIFezx/upvrJtQxYSmLrVtJEegncVkanKFVTCwaeiLcXmCT
/guM/HR17To5fHh3tbcRdkz+MJPnGNHveo0TOXUxn5/eZrGxUpTb5rK4qLFJjV3hEkmX6Swj5HVH
00nwUgOKVsiDvxOgz1UzPRw/4gtnX8tAKbit2vCSuN29uRB7Fr4hpIfHfJrwYNoLIpgCddyx+ow+
Q9BxMje8MbbEorXrKtidtvsyALyTbtnvncXoWrFAXzmVoycsiu1tr5pdBsp0wqgJ2mDmt9XeRrTo
XTBFUY7g0k6/iWgV05DKHeCMkqPNG4ZgyPdVxYEEW3ZHSP7FhTFI2tKw+vCxgdHu7L8XGHqPuyxc
z0Df0F58/sYRcWRew+icX2uRW7FSZLWSwniP4ffpH6vV4cVcPgAWRtFAlodvirpziCpC5YzvdM3I
kCYUEp0OEZQrEqBW6FZTLqG3cL53CFOOQibXbapqJyZV9FH2mRXZKmMvh5NYAO9D83CPP0kxFE2n
81UpU6oetgk2qVbnWYQpPBadrxdM0jfFe4hAc42sEZxemdwxNO9yTjqoq9o6UXjA36y2REu53WJR
9sv/V1KvWVE9cKRE8fIHXs5+C/ztvFzrsqf500hVa/h1F+iTRb6RjsgbsuRC9Xspa45jlKIMh427
ie/jwZJBRYS0+iivKWYp763N5x2NMJeg2RueWnbqYnSjeqVR1xrs15kyHq4pDd84hNqatj+fx9xP
TMaSljEqBX//sbwpvitkFpjtI+FDitowAUOUUTHe5ZJ9RE7JGC69SwJ4FSfOzZvXOB+qXtCs3eYR
WUW89Ad2JlUwRG1vsDGm5jEEokgmHQup7RNIENsw+dDGZpgL3fuM/uxto5U4w3xZ0pL/ojl4vhxp
XX9BhztkJPUuAtgsFnhEExRxSzX9wKI3tZ9WAsIWXbWWfAnYQNM9Mi7QEMcQONTZWq/RySuqAwkC
PUw0pMUaf4sW69ZJzj/EL7J/suSphMkoYrC4jGnA8OcOXGahWDuGRVRUPlfwTilaLT+PnswuaQHk
beEJwyogX/ju/ngyWGzEFRoQvyfEeVEPYRjtOWjUxBQ8evO8XygDV1m1IAd7CWoNk3UTegUhv8vH
D5jJ9jG2jkg85PgyGur9iMrkJ0vaFthSyPw4fKzIXvDdJJELZhwXsKrzLUmOp3IEpCv98FC2C+P6
9o3PPFs7+qJBtiH9u4RTobVWbj2L/5xhR8hMwXe3YlJcazn6C61z72wpTiMSOxvLNR6rDt2be8JY
o6rAkfgOMgDe6d5UBPtQaQOTzuTJCwdizPwsMvivJGJ/hBE5ykPGvhvGKtYqRnKZLVBYAr7dnZyY
z+3YkZZ0AKBLq3wLJMsfdPdq+DRLzLo4WD57z+8hNraB750w9b2WjRdPxczyOpa82KY0Woie6kte
7zz9McL1IoGCfxnVVTbcSoYFWfb2Ix+z8P8tfmoCyKob+vIKscjPJNKhWnSUQ8oi2hYO2wS9xr5H
R62UmlBpPdMhRgZQsJiMsmq1Brl06KJDAturPXK8brEm/bBfFOp4cV2QGDVqjmITEP1t1XAcDths
aJAn/vqF8hyVQNMgEqEarsImQnvgrPYPDWBAF5CbIvuew2Cl5HyxojNcMSXIlNuTb4QWncslhado
9j2V2U9iiBOPyHl9Cixl7VccxqHEEzCFD16tcdoW8brVErjdfv/CuATjyQIa1wJodkuoFwJfHPxs
cKNmUDgdPfPIE5eC7rJjhj7WCyn9gwKcNFYIU7YH9lcc67DoH9i88D8+MJfSZ9pJjYs5g3cLeHl2
g8HKwh2tU8wcaTbaknqX/gbsyazPikamnnSzsm26Ib2o5w05VP6RTD/iAiteri1kj/DumO+Tha5H
0Qg7KzPfYjAHejbnyW7SWqiq/A4If1k6Kmcx4iMfIGuKvxA8FjjKyD9PEPDq1welz4/lG4ECG1sZ
fhkdWn0BDV/Q6dnC2PCBQcZrAh8z3//h9R6jHHWKOF4dm4lJcFkaWO2EEK8kcTZLfAGkzGXUGAHc
KW+S6FiIU6NJdKxFZQCk9/XH9+CFwlbWmdTKi8wg67tpmJh6XV5KP/JuflM5ckc7gph5MqR9FdLN
Ro2ZI22ka+d/3w3fxqtnPCTOGVO3zbXMz+XgHp213vvd04ndmK8MqSTYWA6EHmEF1+Gr2+3QE9TL
WMmG2D/8ht+8tnuEt3GLQ/GwjQLuptM/uigEkMwPcjar4CvTkr4Gcg/MJDqYuxo5Klz0o6nVVgpp
q8OzUCMRtUYJs7uqVr04uzWFwmLvuGMpg5wb0+icoWdMw2oTEpHLmSFBpKP5wt+MA4d/Gew1GDSq
LzVYbA0IITZfUJ+rVldXJnpSn3SdrccSJOULt9gsPUAVUHlUYgSE1R8URI8/b/jx7wxLM7wjYwEi
b3CNslUxcNgQBZSFwahYtaQEKZVWt3iW/l1hHnTb86rH20bNRXgSE/ROpd+6+kepr88mwbh+bdz3
2g0pwvrJXk9ZWSjkBKoyZ7W0LvcWujXFm7xBBrCW57VqZFivAQDwLDrniNT7KS0mQoMOxoIcTLk3
X1Di+9SP0MesR36coEcjtqXhqjwy9dTzBQkrfkNKiMAL3LXqff0qnr0rkdnN6eImpKC4g0MOWBzn
koxZe3Ib6h8thiPk7SFa91+MK5pyYqZCCHKgkrca2mpN5y9VLbNElRTidcqwh8SpXjd1gDDmt19Z
YPaqNmtZaFh4IZFF5P2jR+Urh8nCLbPLhyoOoiEeky9TtlGnQJHOEbw+EU65sTxVks8cHygvQ3Y6
b8BPXaT0lzfe+4towZNfdzDF6I7v78/pFlyKebatvZ/ahI+mUU22CLJAX6I47141sURQd1TEpt1r
Zucz99Hly6sWKcH1yaNqmePX4rkrr7w0IIoINqVIBKhdz8aCTBJ4jbtgzcI9b/U/YqtEABRfqRvX
Tds2rtazULk/7jYDYfS5QhtXLvZyssW/z6P3203kNU6yoIMWsOwSBagfonCMcvYjTcB4ftRKbahm
U0TTXNYSLczjpv5y4XQDOi0FkKa6EW/05DOPazo45yZ9mRw+0/QYLzozNnAp+xr1oM6eUe/LGHuk
CqzNhnXA9RasQjDqf6NvwRdBMCe+Be8gdhLlb/NTC5rTnU/ojIczFqO24MVtPTq4W9twv99HThmK
nSzrfRXWa4G6lU+KlUSUd9qgzBEj3yavrip05iPTJvuX30VdL6JnXnNna4YNmVlZjTOvoRQaEFN9
YtVv2oWR6GIAMqL3OgILQlLouelAk3C55eONentoL3ixXZpo0Tv5Dj2XkY5aYdM09i8oWXL6Oi4o
rjR3ZK//fg8TSFIKF+drRbqMkpLHgbtgthzSPTo8Ft1GUphkXiZ77SFeXqQRS/riyw9xuXR+FGNa
JckFZSOWN4Age/xgLoGF5tJ63yLenjvQ4E9gl4uZOmE+geUprkEhzxdQ0tAVI3YgZqReGrse1fdu
/aMgBO6VivJHhCO8UNwN9LFOa65TZ/a9bkdoC9eO/fYFUhysN6qXVzOda17bZNkT+//+WIj1AfLG
UJTqMH4qEko9nmLZmk4GTKdnElZVvwpSlqC2uvyu70EHHgvIRBe4/PvUQNPWOyQtzY/XbrGAJfGc
iQygd1FVedcfd+YpEkA2uP5n8JXqDqw0zdhFAbEd8d+W1fIAA+6+5UXLQR0h3mbGqthJmmVh+uSM
FY0i8SV/G+YVRQZCoXv6XlZaG1l98DTmZK8HXBe9JK+pSL+kZOJycsFU1Sj2szeXhVhy78Br0gBB
n2C5l1/UNoXuQvMhN6+Iu7GdRsq38Jt3Gqykdg70f8VZeEFGzFzXP31CYK3MYn2C9HHXMOBdq7xb
fKlW8qlZQqxvfUHyveBwVT8yZmZkhCamoU3RreMtwU8ENA9Zl3gUjA6GUb7GC21SJWQYLyXRzV1t
1ERmpII0irQoLciyA2eCM9706mytzQ9njTAhvLcMt8LNg64pNi0JbODQmPO9i98b7qIhslj4b3M8
qgXEYpRcDaEgkkQX7y3HrYEMeuPiC5UbZWBnm7TZuQCRUACH+BXw78q97wmJmWWHTL35fJaseynD
15mFfjlqcGw7CTzaMbiqgB2UJXppYYyiULAiFwgJWy1r7hOfHpTYEMd5Dc+a5ndr7Hswjhm7HRtH
obLK0dbdndseAOlMMbWudlR59pgx1koTFyK4HzYTppiBv0ArCl9kRb+lT47QRnMXaEV390CpmN5w
rK/e603DsRoJz4fUf9Z1Oq44X64JXEsDrRMir2Rn4hoxatUtPxQu5e/iSorzn5N0ikAsJYp9Wrul
vsad5aj7CLVPa8TVRbegGywzghLsTPChY9xGFD4+CGfIFOPV5iiUa47Hz82A/ARHf5r6lzvYR2fE
iKaHxDdWYR9pTaujQfhlt2EIz4gPet6m+Pf7SsMFYxF21zOtlHvwGuIYlgyfWNZRMph9TV5tcM0P
HJkOZm1ZOGWl+stvJJdKzxo6EoxfgJJ/+lvEeT2uTy5IAibIi4DpU+pBYdJy8oyNHsMn4Fei3auh
0i3863ghNPqbv4JceqYptrbOxyBnWvafF2ZvTwEt46HarCwrrCYUQkEdviu+zEjaJyv8QS+8FRvP
nVcXEXerWWhr1MWwIzTEHbfqCw84/lCXk6XrRI98e1FarvBnLdCtTfGy6k5UmrXVEpUnu9xdqW/T
wZiHT5C6DH7zCxzkavaTkCKf6f76RfJT2EVKdeyzFMRQZTO4LbHg8BRmBIrPKTwdQFNnjsjiYway
9JBhjP0y6G8NYwegZm3kXTwDe81PPBndz5Qf/xMVSGSMqjeiqK31WT7ohFlR7lM2pfIJCvdlMbxu
QLTRaVBeuzeCROjdiB5jMbadeQgHELyY4rSAUF7H72Z+Rn2+2MEJNCvn9U7EVEeO4eP/4rF4tued
vqsL91UI6e0E/pcyN8HX5Ghp32ZbRsNObh4lvOBadW5dbz56UmHJL8tNHnoGc5BUw399Jt06EEKE
A9L2bxm4Jc66RuRY9pmd0yANYtzy61Z7yVSh6UCuRmjNgRV79/xI21rXba2gocgn6P6EhOSS7FgA
K0TM+/J7VFmSDYfj5yCll7rh25UWPi48cqLJaOLF0Z8EHu9WVpKFmUKuxS6xwg99ve3iDkfJP3Jz
yk08+qF/SX98UE3Gfr0m+bGpTFb9nd688W7fm596N02DwHXz4UU7flAa/Y7pzJtzk1iRR7a8oMxT
WLzJ99m/uIGmUJ/FAFTQhc8YuvJnbpYPrgyx3arXq1edfINoD5iF1NqLThjzFPWOVh7jFtq5CfjQ
7DuQQI+gvc16xM2PDODkZVfuM5hMNwYRUrs8572N6e/tjMDS9yTCLionGQHt0Umsx7F4ohQYCXsJ
Ccohonm+h8jD4H+BEHz9yI4RLhVnidb7n9BtuWM2sGmScWTVQJI10BnxNdSSoJwVbk1R5oc1/c+Y
a/W+ck7p9ORo+a9eM0sViE7F2YAHZjmsynqhlwEM1RcjT/x4nCRQ7MfjmjSgZOaPPVMBKWhH8FlO
8EHIF3/25Mm0QESjxZkMhMXiT8P9+ZGFfPMVRqVnMLuICoNzUEtd4zLczPOSL7663P1X5XlGYoKg
EH5Wn2BFohFYPp7X4s9J7DLfRai7z042na9b3NE/Np3dG8gafnXGvcl2x1dfdwGQprbHDl4CFLDg
cpsRIJAksXzvxPG/oPm8b3FyKRIw46hXuiG2MBDGxR7XFmcO1Qwazk2Nd00OPbxtkBzY1tVNeKck
jnZRC7icA8vjS6Ve+M3HRGyb9GEVhRwEsNQlcNpUQya/M9vap9y+uoXL0Mem7LCQuXHAEX7x3sQC
O0FhBRHPdlBGUXi0pgw3fOjrPbAjujGDYI9ASOY/9HKFC/eXVKGf9O9cbQcOS8NbqzyPAaAKElEf
V6iZ5SSHcNPwMyrb+kaj5JD0FLG0qAC7nreaCEXnR3cIjJMFgjNrzOLQMzmObBbwyBwu+2/Mf7mQ
Yz3EWkcv1D2BIDnmyNZpDvMtCJE3V0HDkqGs8evKtGlTK8zfzbClxKxWQ17fOelLlw+E0lZTVLyg
uoJP7S6Mx+/fkWypPTGq5iuc5xjRpmx2F3rEE3E+/lwckJpAZ+xZTSoG7Q6UaMhUhr0CLZsNWc0N
/kQ5vikMN5gmorV2qrZ4zOJX0WHN0+K1V5CopuhAtiPDCryg6nWx3fV1yn1wQC3wagwPhzyQkiV8
T3SixwLzb8FjopyavyJGYHs3a7r0Rh7lnZYcO+EeSpTkcOm5iZPZAHDRt44RDIuHSf9QkgfYg3tj
zZReC5uk8UMax2QGq5n7V/kfs6dCA3pufSUGGsO1surUYKNVn7zUiDtVBACcVb2tTTIcZioWxz27
5RqdLL/9ng0I4CjCsyv2R7/U2EUsrbZztVbGy/z655DvQCwlB9bawC2v86jGQfrBLwX7VJVFMZJX
qq3aVoq3zWSraR1JHTvFx+6OjFPXzVExpfkWgCrQuZXt99Eq/6c5hKDknFNPsSjk9cT9CfzqEkjO
momHzaOch8PzWIlG7b5+PIsZpLBzRu+99BHfVNwAdm3LwtFmpc7zwLTW3t9Kud/9ckSsOJjHqxhn
NBdi7jinTC4EG8uo/ZBiFiAfNsRz3BdO5GVCKhjZOubOufzSc66zZZndZ6Ho7Ja2GsNY4gy8wJ+8
IBuM1C5h6tkfKOgnwI+J9vuRVXwSqm3fTZ79u0jxG1LENLFAG0WEkYp3JSD1vPQ958WG+UcdDa0F
3roTBgBrevZ6qIBLeai6OcoqteXoCi+Q4LeYpxDdqlxvRbztgi4sCVfH7YE449C7S0S8V7I/dUCO
Cf43dY1UhyeguDofiKR8aASKCvTx2LavfSyqBSP/L9hlaorXMm+AwWOoXZWr8/dS+6u7/BWz7kTm
+KJ7yQ6QMJudxFS87Qlcv28btFbHe+f5ZFOvWF4Gd7LgUPr2samCPcZ49uuqyeLQGMgxQRBkxhqm
xtsB/fVRCxZ8rpe0eqwGpn2z4l/OVHElbk9+pqHm8vI5nvbmElGYb04F3kbLyyjus0JZdPft/56m
R4LJGgwI9WF0MbJjS/AZ40gW/e+VRHwto0Gd6ly3Okhq9ekQjq7NQlLrjYBqVxdFW99iggPtrna+
IYlEmffGCEEZzz8kT6QjWQQ6/USqTDbfFRDgQqLnIXJTQNS0cSNZuO7hpxMRtHVO8uFoKibkJq6+
DXjKPcO5SIK1Gxo6FbyzOoOsDOjHWP8bWhjrg8M7HhA0cdredOX9Xy7x8PurLnS2ZDF8QqXNO5H8
d0wZ1FyyveQF9a5ZeGd+WalaIj9Yd18p31d9bgv2AmYv+BOBB+NhgGDe5AOlDYmiEvKZmeRAmO8R
m7IoAiQFBAmRJfoe609+yIlyRuexUkSk4G+yp3ZrR2bFNk2yxJ7yOofs4L0WY5ESeCtXOHUCxBYg
YT2kkpb2ibLszhQRhj7bkq3NtLS1AsMsK9tTsTye/IqTTBcIZJZCikT81MOm5mz5ilJr93QPXHu7
miRMk9fAEZ8T0Nffb76BLIorU88ykU+JoNmtJI4DQVN7bUjGIDzxVikyVoompJccl7owFVFBw6Tu
P977TxHBxeysUj0430XqZY7ELF0ZPz2SDg2TMgG5hqIARp4cP75O7rwLJId5hf2WW49JCqB5AytH
EH7Q7hZypzzQ2OD6zQ7BUTJqobyTX/QYzWFUYpZUjwGf9a0gnQFEjk5xGLWj/InGNfFetGHh1GnG
1EJABSfp+DX5X7UvJp0retJYwGCUDb0Tt/vKUNNchG6je0w68BjQvnIP2jKG7XBqBXfjQsnl25Ox
fSAKncJOI54YJjbI5r45Uhzrz5DJpNvyE/dmegyiDFVPEJqb6FuRgw7kd3LhuaNqrDJH5efjdfXQ
x8LEs9samXD1ZoN1hDHLkFGbTc4hOCKaxvCgYPS3hTkjft36qaHKJ90WxkLCfNGg8pnhOmSsjNxb
OWzeQmVlksqydHxfix47kdzF1ETirYndV6+v2Jiy+z1sWehZ5IPWxBslTZ95wP2AFFx3/rH90L8y
1//cCbY/yho5Y66SOdcIvjEyJHssqgwvlEwVeb+YUAEFVewgQHLHjhu3X0oGLPeFTBift5y8DUe/
7uVgdhxs3y6mujFAp3eOT7uD6RGXd63trLoZMMSD/YAEKwzH54cLaPL/5C6JziPPT4JmfHMI/3Cs
0PqaeCA+0PD+VP1w/7Miprog4m3IrB61hkMVZf6F5AeKbAlmqdxmAt9YeZCvD9B4ta7PR8LmqlLa
C6pZ4rwhUKSo+oGPIDwCMVIEf67MQNVNUl/LhGSYLCjyZUzgnTZjlrTKJ6MhWtj+2BNwiSKi7ye0
W8sEIFtyZH7JH0mG43pOrZLez8kFDS2MGoy3YKXFfZR1iEBYaXntrn/HK3xBQCgZFiw958RhUFC/
BsjLlDHdEx1QMY9K8bH0ljktU0RJ+UjzKE7Q0NwBN5nsIuMc8GMeT9yzWBVII5axmoR0BL5ZjrQJ
jlLXdd/W+RbX78MUHwMyIjLbYjUTHKfbDBjBb8Is58a4Lm6IsZ9n1v9/0vo95yWEYzVM0vzOSXMn
49KmMNeg8Ua3OfP8j/LcIkVO6Fx8HQt2vheGNLEw2w3qvow56UWDItzRWtS/STofWi1betWEQnNi
WRXXmTs0VOJFbBd9YJZsk1Qky87NLLZklqikWRmBdmBp/sWfEin1Dl3NH6hbYxejOai9DUbRYZDc
dgSPTQQbYkWekN2zCnvCjeF/tlZ4R+wKS1kUOFkWeI+fYWvC/WwqdxttjZxyDl5CnGPqRZOvixdE
3pv06oycTi+UIrBuyhorwmi3jDbrIZCPhmbVW9igV4EWBKTwESDr/yKzdLAVlcaYtzKKZ/PtfDJm
Ff4vP95BT7qKXl7TXMtGTteRPWqS1mIGiAkvKhkMhxVuol9lQiyeE/hOUj/7BBXpZW9W0LF9rKKD
sDNeuSuJx+sLSKlWH/0ziReEyDNral97xcuhOdq8xJGjuyhQdywNDsM1cTeD4KtziaFNA4Kyf3XM
kY/Fmal6N8d2ZKIB/ffdfn1u5SKRvXxCsOYDxJARdlGRAX+7ADOScLErfHBspTLgclHNBQbeGeY6
gNWxFJjb2p3ACpnQBGPhq2cqkF9NMBBkCIvSwAn7tLZYhFKwXSlVxchoMNP7NEOUqN92SVS1HjbG
C4JfT479AOtU2f9Gm2uxee7ASWKAAfkqsvP0QkfvJZ90kTIZTwTEFZeQSkZ0sTOGtknVJpwff8Ur
cYr9Mgqogvn3D5C1y353iJmnto+1/rxBC4WAqZeLTXqH2C/OWQMxfFhJ+6FeHCmIimvPY+n3M7Gr
7s4J00AW4h5BSWJYDBDXPqEnh5QRZWK+hngS2OeU29QX8YOWG2w/CEG/okFA1TQh35fPIjMOtUE9
KzrOxJTBl2M/+tR1QZ+dJBT4GchYvz41ZjrXYCsPpM1hgtsRrMP5cgvcns1527XM/oZ2RIbWwaCz
JMDu6jVqnQ+rqYXFLpX9orFQVc/Xsd3PVNyeHMLL4ICp3tFN1HantkEEgIR4KcRQoQ5IohUg/j0c
bIsjOl/rTqVKvv8r9S04485RNCA/amC2XGp/LuyN/4gLIKuL1+eXEBzaSLNT5b4wx4xhdh9Jd9oJ
sxbkXmy/ffA+VJs/6saGsGPy4OtGIvPcE/RN2rmh0Q6jn5eGptTDGdvJOBaCqQevlCb1HsUgAEUn
DcX8vDgTvRohgRPdT2Q7CGnEgaQ4ng+KY+Amj4sxvUpNux8f5OFYBi6nkNVAGPL1b2N/dcN2wGXo
B8VhqkD7HFFGHNm8ddl1wmCwT9/cTz8LZU+GODNpwWz5IehN8XiH/6r+HDM9z/niYAkbBx+TPKft
tWURKXb2VT7mGPaxDoymYMBucEjl9DT5Ds1q6sLWPRqcLOh+qGNl23bEw+gbIWqyfpSQoO7QlEf6
O13UuU1cV4UxQAAt5QtaNU6Afs5nbY2q7hr345D5UpEMT13FfVlrka/W5T3QcBUugbl+A5GlYNzi
V5C87C+GBNpNtavtxbBJkjKAHj9Bbgntxx0nMrT0XiOy5EuPJcxZ69gdIT/D4zjYDRINZszeabn3
fNmO8TNljoaWtBVaWiIHnoBA+OnBYzbDR0YOA5fIHk7aFu8rKkhrq6gaKBC8vxvfq4nT0WblaE4n
8m1r2/8nloJaql0bCYADWWcEHd9QOUmpL42sCiy8DVOoRlR7+yZHKiYkeOrTsTKKL9ao2MZLtZE7
wP2ObGRXimJ1uhT9iN4hxu4TJIk0/n5WXMLr5+GlSoOAA66HsjtozIVkS2DC0cuHMPvJOGxZUjd+
EVSpFoH6Cn1kj027fxFnPipBDd9aPlCNhtgOzM5llr2n9dLxn2KJyR/DKsI7SzlAUARMKWWzXT6f
hRRh1XbViSMWJCl2TYg7wMh7aOHSY3afsHJ9x+Xa7UeQHGC2dNpRuo65QijiEY/0DB6d0hKmoSGW
J2ahfiU0db3vmplrIhy3oKA7TBXHd/cVmrPVNJQwJL2EQOV/KhMOvBiNzHIVtsjoITYPLAbvDTMn
5OZhlK2QJszRREyWnfM5yzWN6cGeYcrbqoXj+qzeG/sonPJKGBx3bD4TwmBqZMFt2tpreXZnJCmw
6PFC1PxsNlkRAu8FVRy3jNjxCLOJgC1MZwFd4qKKGYyEC53BoITZpBTWsKRg6UN7nzakAjrvtJ2w
8EaADFgUhyN2budBVju21JoVkp/mBzpQF+LXk5RiPcywU/QJ+DjZ8Esu05eklpaLD/47eE4o9Bam
SRYQ0CXiV1h7sFMGDV0gmVmd6Nwy2AEL52Dn7m+6Y2mQ8fnfd3dba8ubGHULQAK2o1iLD+Ah6JW+
gjWR2LMVmQDfoWFOqk/Uu7L29pmll1FV1uC25xxIrLI9QIc/8CfV6ksTT8eTpM4alEvlIvvlO1dy
DzedMRbYJ6Iucm9yvsp6MlOIac5O9d1x6VFANJTCJFWPPzEfs+b2TAxW82COYJ8rRFlxmPko21ij
9zX0tLdP8HI5KVUe8QQH8MvAVu6maXpbTPhwxyqocN1laSiLuzliEvMyRmdr2XxMl9v7ITRvyHdC
JtKgUGXA+W7Dh8uZ1XlVdiv+75QKzPLMGCQjOnm8pjQNJQWai0JK1a1LF+sgA4tjRt5i+3CxVSeC
poP55zJCJW40fx1y0BOBW/Uk6jfKM977SCzMVtkjbWCWv/1q6JFwTXbHFvIuIG/c0JqWVSnxfF55
TGtmv9BIAjkI3oOq4gOd1ChTfeX4M4iByz9mEFxdow8P5nBRzhtonu4tw2JQwqPVsOdx6oBa9xOV
m2Vo14U/ofF6LQnRcJY68Zr24ff+w+Nnijj3+Z9hsHALxcbDPvPPRisXIFHro7U/xsrDWx2ZxhMp
NiyUC3/A0CAMkBVcUxVDJTL3i4fXcLAlO62NkDwq0hB3fsNzunRWygxcqG9bcNZwEBdAcJuW8vI7
uX5Mp3gMj8WzPA9xBTIPK81OeNrwcPtujAeQtBOcOrqJkXGYaMMDG0fmaz9hGsRbQUMw35e1x6K+
8bI7IPAHxAA6/x5XjOJwgpFq+YSrCvsa03VRVEWp4l14x1DxwQbnfvFJ6QXGP+1RjcXT6umsBzQq
LPlCUYuw3nprVdH50RTXtuEbIVEI0a4x6N5cfm+qYfRWu9lXrkzjOBABCSn4E4rA8y4LYVpBNOLR
eB8HLD2oAHWf90kYX3QhOH491Ymzs5GLNlz+l3/ZelcCIV87hWZVwUWE3vuNnbNsBKmuea8KkAVi
mQ1G+DN+/rrrN3bq/tBRHZfJlxfP92bU5XWaElGTBFsif9oyWovfG2kb/oP9WLuo71MmP4vnv1DE
CMV63IYjHr4Pap/BTxBgwWUn4MpK9CI7axmexMDjLEIRKctpHwWWLiczRkw5j4o0J1ns94MzXuxS
KhQHU6k1EbvFhgPDK69zqGuAIZVxtRElZoDCWjCdcof0q2ZU8R5pCnYhqr3b9RhGYaj+Lc3AE1Fi
JfZ8GyPDjnEIZ3eEpH/37zEdzb+YAHCC8gHoDBRWCiXny3t8o+37oSq2bdumMGmXgr16MWuLtSwl
94xMDRN4mUQQMs7YMsNpqRvYi6CaKbX9XTbZmeyfqeURU1JnAvAa8fJWtkSnzA1vATkF9gNrRIqp
cJaCnijnSeLe4zWx+s3kFaGcFFllWhzH5/hgd+dnfYKG4xzQWWuRCGuWmJYpqNjnD3k9BOcrWrim
7xYIE7Fn36VtSgkAnZTY9bs+PuhvvjBv1q6x8pt1lez7PsG/apPVmqBCRx0HI9TltwGNYuPvp97g
zT2uEhByov+RZDlLDGwOcnro+xLRq2TSOpQ31SGY7VrzK7+z+VUJqLOQrz6YayfstrkvQRprQQN1
/9m8iV0M4F41TPtrwlam0MYyjTtXEw3V4uaovjniFBk2Io2u1lHPFIcwtSRQm+MrYiOUVCMQw5NY
ziQIdR7JXjKBA8u1w21OTa/7A0ta/ogHugDhujc10XnqklacMe/UTPIZM1qaR8ctlk7+cu+TSj+n
mSR3E+JVF4AlmJiQapylRiCTgDZmfgPIs72bclkMSGveDj01nh1hkp4Rc4sBN859JlraoH+9eqtm
kA8RpUTifkEQM71fwVdrPeZtzLHWTwibaTlT1jf37eCz/FNvGqcF3BySq1zfMIYB7kpG0vq0Nwj4
IWafisy0FCT1zybsTX5hUkjykTJcG6wC6wyRd8QYe6pkQu8xatB8mQu6DvU0t30ey0/rWtolOxgf
aYRl0Eq5iMf45IRYThPmsT7tdyYDaOfkesaOT7qrTp4PwPJem04sKzM1OvI2WCgSUlNXbftiYzo8
Yik80kAI7T3jICVMfJpoCR/fbu1dJaekM01Eh3nr0TmAliI5ZEqYKekXpm1oYntjuQrVuFbI5son
sw7PfqGDHI8UF3jOMOkmsyGTqtZodb2yrcPkU7Euu3gWPRbUhk6y/LBPUGSOxGKWas0fXaz4ZYND
c2zNezCUkppqJGsBm23yyqBJpfLRx6KbE4V9uMGe3t+tXDmYrherrYDjBCYI3elVG+AR8Sf9LMa+
oGhY0EamfABy4qSvpZSWCY2RVuVE6RghKOjrvF3Ui8bo5lRF+nj/7K+00AY9Hu6lt76HhrVduCDk
Y5wOWH9gGzhbURYEp3Pa+hQgqgMn55YW/w9boytkakiDnSzCLbJGcijWLQzKwSHqT8qICG67SA6k
x2BJGfnVguu4BbScHdYLznUmqUuYue81miblmfKXqmV/B6W/tMLvtny0MlDvJGHl9sW9iEp4Gp77
GYeKiRmnAipXmE7AdRkFEFhxmHsWrOQcDKoc1LWIpQq3UdIEMn8ZBV8t0yQy8xs3esncfu+q3Y7l
xr71sqnoJ0ytIk8Q6RVI9UL/uyMtIOclIn97K3FTqvbb8VWhOslTpXAGZK+Qcn/ldyDFsfJt3U1X
u21AK+OL+8Pu8hrWXDBvkotTDyhhEmYONTxdjY2b8qmlp2GggD7DOJOw6HXkCanyLMm4L/4FkH9v
moBczwrdMGAzULDtM83deIT+8aUKk4ICDHS2aOtfSdkBwS9hRKMYq4gQy6Krb+W0otodHBx0g4DO
MyubM8FvvAA9ezL3p5EgLuX6513nmCKqc6/X4yEBIvr9VQcE3jENaJicMqiGMVG5QmYc3mE/nhtq
6yPx3nMXvjF8c7mtn07ENscAVHl8inXcn8ne4c4CA6mqzykeMl2Gf2rUy8u0bxFBG2uVbECqkQb7
2tCq/bfGWs6eKFYqxtS70Q50gtGGUajIIt5K2orgFrBR7BPkYsR+LCNm8ClgTuSbt5MQyZHhc85G
D0gcO9kE859MtgASuDYOjHaf6cpeIUvCOo1am/PbqwDyoTWLWlMgiujTCdskr1/M/praYvFCx6gA
Rm1qIyv6xk3Ab9nM+gXE9Fj397kO4owhMcobSUHayF6uhUWWJW+/Rmk3FKSSNQoLOlDNuz70sFxP
rJc0b9uOfXIlQdSsGgPMhtKGii+DpLXo0bzbQpHAeayxhvmXfjQzJEjRc0PJDwvgRR4x+QT0f1dE
e7/ao2FMGK4xXtBx4nu25vYFyVJtr4uVQeJ2lNa+Lb/Eklk4PsmZEObbr4ZFvdhDhE6l41jHV8Ii
tJX4cP91LwPw7t1PgN5FMxamow6PtHwV/bMdlYsNKoxDzIFcXgV9xf/Ra2tEHWai5SFCr0BiLDBs
jPUofkJusHL1oe5yEsVEqBE/EG8OmOFIegHGuQszSLhgWpphd8nm9/bZ8tx+DBcNDLXf+Ti7J4IX
P7C2pEiulhNT1LsDdAd/VwsAHg1xPad1U/mlqHobHYEm866w6pkKvs8B4aFv9YZX9KpQk6yCJ6Xy
v12mGHXWLSKnUCCssFnacr8zr0Qrk6Mik0TSYeDOq27o8lA1DuZ3BNAjmky2rF1sQjqyODuPjMfl
0YS/vxqEwfimUNw1SXiM8iUmcGnaqyLP6xowZkmI8WXb+pA/w6N78DGNAxbQBH8Px4PLW0Hqvitb
aucyAUmRN+AowAz3KIbrlcupDW3kYinzuVyE618m24taqWvp+YmD+cfNl6gCJmbfdN1hrDEClB0L
0KhGRM16Vt2jKmTy2bAnVSGoCgV91RKcT4gzdjwHTXdQqB0f6cK2THPrXrdPQksUCprAObIEAbg+
1qZeRxNc26Oj2Yy85al3OG3DOvXDntK51MK8DwcJ/v1tql+UkTpbN5LhXmIA5wleydFBoc/QaDjW
Vtp3epTTWQ12gM9a41FXFX2MbF7EqXqxxdMQSJETVZaTGVfJUG5xA9SArUzoKNJXGjgvsUwRdQjs
wsr65kZy4fnqKpCy7KgpKxGVXH9KJWRSZqfm2WWBqJ2FqXPLHI98HLkXtfK0LDQQ5CYZtcMGqB6P
o3LHM3xV9hBbAhsCYETWWShT9L4u9FmKhPvHVCFQbwzy+KBaEC4g6DuxfpgsEhd/NR1iKiW/efm5
JHgbHD4YPu3fNYjwC2GdXHwYN5SdnUfSj2Yil9Lzy3qATkcLCc/OImWWfEbOJTOBM52iyRC7hi0R
iwTGQPUDaBeYSz7YxQVz+Cumfsyj2/0sLpHpDjfnHiAPCdJAd7rSyxwqCQlcCcbnYkeZGElJ2tDm
OLj5F3jPnbIyp/VrSPIoapzAaSrJbAiaLKaThqX9LSqkGPnwqGAffWCItBd4KjIJx317T5gnabm3
Jr2rJUs/j0n4QSFumlDoEx4xccgbpxx0hLYGyplS3O1qsjRy8NFcP6KYhuK2N0x32YDXC6zOPpMN
GgXrR3xOWt8z4ZK82+vYB+45jvdKn95804OYEbnuUz+75kaj9C2q5svg6Jm6Cgr98gU7WMl7MbXy
wEomhM/V94pe197KRJ5PXcQo7Bu4OPp/IY2zANevxs3BDDw2f0/TNyOR36LoPm/Ases+qarJwcPo
8ojdszMHZ5529Om4XHaJLcNFw7PfOMCL1ZOXoPCI/6A0AzeWko//v7ebuE2VtB4ssTwYH7+tqoSb
gcdZE2IgkHvzNe3uPPhh1t3tmmUL6WHzC2L0O1Y5LVTEseBYJFT+ARMjVFVrNz3RrNWZE49hASWz
thSXh8wOUUk8H3dgccgb2BLiVyLZ//wW63L0C96z1BhN3zjURPhruQSkftTXuzv/bOpINitkocO8
Tq+6o3LJLMiMpjU5mFzynHv7f5iUM+jvxu0L4DydVfHfgkOjafhz/L/MWViks+d8Kiiw1zcd+ClH
dQnvdhsLj3kY4B4sqvGjU3YlCbvzHUpV/VSLwWv999kZvtl5bOU2Cef+DIoCCNdkxkiPGh1KLVfa
Ati40GAAbMeqJeHH3CjcKaiUBTbYdNHFEQBsIjr81kT/RIZJaA0R6eooBAObOuu7iiLbkzq9Pk3i
8sofn9U/YhtFE5O4Syy1gnU3Uv8ehl3+EQ3i5GyGtm0sBmUTlkvK1ZxyqYFaQKgQf6CuDPKizhBX
AbgqykKb+zTaWcYSx4Sc2McSLDOHATJuF4/4vzTz5sgEsMH8h3zGa4PuutKyyrBYTwwq3VbziVji
iV8qbi5E/ISZfUYUhV7p1EobVYuyffJ5bDkCXRoikO2vJnsQG8vZzOl978+549KYG0ZIl2F9ur6u
TIYOci+zj/5/NRYi2NnTGWbi793ny0ghK2v4I4ZR5mqcm6lal/hQvzwo4O8ICwpjJj3QKqcTiB1h
Y0zTRgGTiZup4rG2B+wmnjjkntOF0qkGAkK10QZDuK41iQwmRT9ciRw3RU+153ATM9R8jWZlSaZ6
EDwH2tm8VPeOQEW/NNse2yCGum5kkpAd5Xv7GFpRO2v4Tq3vazkRAMSiGdBG0cWBYNpMiLcjKz5w
t1jpU7irELgtqQtY7haE9kTNj+i71fTuWibBLSXLNUTePE07+KTO44pVbi+96EGWyL4BtlPOhFCX
qB+eEG15+pUn+SgzqH67Gvcwl8H3yt78FZwhxmNkuRwpQgFpiEkf/NYJCFLZEcTtK4MLoCFBhzw1
tNbTgrgl0YD/7rNuWPQWNZzEDbQhyU3Cc8ZWRpnMnLTG0s/KiniHn5Tu9vgWZF3PTqGaoTVjPbD4
V1OAHuzbPVDnWx8dbJnWIefsDE65asG3a8425PAVwR217/zwi4I0vRxJTgmUZ1MXqPK0OsYCC7vB
PxY5wE9NJv4teu2QEzw6WiyqpT7nMjw9Sp+oTWt9Qg0vg4OCrH5Us0F6UMXZ1Nkq7It64kLidwfN
KXMBTSRt/ougeuNNhz41iH8FnWVkY/vGdNfzjsyJlNjMDsO2A+sHLaWyrztqswitOj+nKxYFDe6l
fQzklG/hdPkOcvApFFfGbppH4HOsiouu4TtMUvsXpzhxmC47l/5JNe11Bul3BAC70czu9oKlcqYu
sRpaG0tOz2N6SbGgETcp0HoDkAFJkmec7OjIuwCJA49Gsep06YUmDaoQEvqgk9e4LwuRlAD29wNt
pz1MA8cu4v3z6RMZDixO9I8d0s+2VcOL9iBNCygYpy9hTsTFwcCm3trJTRL3IJdhqX9ldJ5xlW3X
6y2W4dVmYTWnxMDUSY/ZxwDuy8yya5q8J+V5Aw/Nac9A79RNi+3LXhdtUGVkxnVd+fgq/oppXFmI
eyueXxmQFXaTpfxsyueoIK7nr4VVKLw6pkJeAaF9O3+syLF2ke4kPVOSX40KQ5V4snmTbDHi+6Ks
3LuAqNVz3RY6VzTp8bu7BRZ5Q3FS6CHcVtcWF/5imQSaGzaSIn+vAyqyQCJAFLtHbYvP2vDeBsU1
s9DjAezD2JxEkJEK3L+l1RCPB6HAz9HzSYNOWZDPsKrWQdao/WRfh5PBcSlxZH6hPPscjkG+HzLM
YcdRQUCwwUmkjMUsdCnRx8MrJ7Df8SkIAU3eq+P6RAMnXqLlVEtu/gredrFj4EMcUgui5DV9dSzQ
VYj+pretbAsBrM9O++rBneMDsdx3vsBK4MsSoqF61LUEOv4f1BspKfgg2xSZIzLKAvL17LUPPo7Q
bHYAN3GqkWRCyjy7IDU2UZ/ROTh3OkmyX8e6dwh+Oek147SWD/AI4Smyxobg+1Jy3N6+D1YD93Ay
QAar3QCsl35DQ9EsWkn03NnfcGm3BzD8vGX82HESJlcNSL/oVmjLZN3sWXZZMzhSmnGkRD6KvrJy
qD6nLPik3WPo5Cy1CGnzddIdYC+FtGAIih74nFLQRG4eTPlSIbiH6PIvY51K76Ps4bQW64nPeRWD
LvD5LIOm+pPeUoA1vPrRN2BzkDJXaWh/Tny7Ipe5i4aboSBcEeYLnVF7vZsKCQcimXoL0KgAC2X0
kuabWBnc8u9Yqrss1r9sCfqcqUWLYaqILckiv8PgFrJQb+PFF9UELC/Cp9fJs7ZOU4YqZODcg4Uf
whW1MafLekxmiEvH0yLwdfzZBMYsxgTeEk5zdKO2XuCriG+JTVZgaRtsvttmG1Cyw5A6Mde/Q+Vk
3gYsEriAMgupW8XpKE1TNQ7dZuDxihFzNcdzkMat5huvGyUQiTRTb7blSo8FjtLHpgGAOa3HkBsM
+DWehC+/7efMyVfx+bM9xR03bdWx7Dr/LGZjpukBhsnIhzVnowoulslr3PUKwF5+olM432vijtXm
vpEh4J+1X4y7fJuqoCBB+M030IvNeHNlQgmz1NB6qfaUQA1XxOKFlGpi1FepfmnWXBuOvzJxobb4
TXDK8QwPo7fbR2QjOQEG4fcpSr6bQynZNRls3F204iGA21geyKgfP2nIj/8BNm5Q6dqVYcs4I+uq
VrTc8Fs2WFxMe2Zwetl3yJOui4HNQy4JgZDU2mVO362SKMTNigO1lziivp9gfTFGa4qHgaS/XJbo
OVtLQipJf95b5eeeu//l+ZvVn4EAaHoID0tYesLd6sXEv7gwKbiMT1L61JacjLUgltA2JP6z1e+m
Wa7dWiIvIB29OlcT/gyejySAaLZ0ULTljU+WulsE+FOIsRidmU3EE2mcY7HnALR2j3hCgm8V2VFq
4PluGgxWdnEl9CCYgypaeJH7zykgMl1KGwrg5jQzSgsgwVyfQgjeTID8FrfozynohjJMVoc0GT3G
mNg5331zmJG/uarcCskkZLPqj5tLVbhm/DJVSvCw5WQmX7PBDuqQo+acHrmKk9KsOZsp51OPaFUX
AfW+R4VE/tb1xqTgM+ua9zeNMxI8+rkfJ7a9QTBEGKFYLZHpYIek/V7yZ/c3dAHnZJeEHgCTaBD3
VMjCaPa/5QddUVWclzCri2yNBvlplU/3p430AZoFxyBTgl6g/Y6GDtqrsqfoX+K6/fc45+PbAzAr
yu9Q0V7HJSoSGGTyGXCkh6k/fXytNMDcz5MXOO5hIE1x9+HjJ1XL5+3Q4Og776oFhmMbNcfRjJN3
5P0MaE3ii77hXlYm9GV9OFIDWhb8FscXaSpfUgWm3Pb2eBqeqiKJqGyq916aepyLYZt9B55Hau4L
V78LlIKKkBfM88XwESMkrktGyPkof25q1hzhqfxAPlsdxx4Ize6ZmXc/LsgqzsMVIZDJURVeRJ/6
YRn36igKj92o9fOYYT8047o07JOyZ0yg4kqaZ0p1abE2p3qOpdrjLM0YisUeInZAmYk4X69CQC94
5DDOLJt4noRkYzzuseNIb0Xq72QfuMTDE4hH7w6GdekBfyKqCRMVVfKeB1EC4f0Cd7eeIMsjsv81
uTro4MQ//0NvRV20dQeVMeRby9QzWfiFcgjfJb9Pq7DA2TcgT6ISKbsDXWDVRZV2WqsqHpeTT4By
YHgvMeVGY6xsQOJL2slF6Sowsqx6vwKlVJK3xqxW8IbnGI+MyNH4/4ktSaNGwm2Yn1Vj7KcjDGGO
uAInmfgn14BCPKC1I+5xMcJjt/mJwmNaiv1H2xvWVre1p9rd9hm4pYZOxjkuMjI7VhZSHaFaLjdV
Vg7BSQHOVEoLi2Wvb1ETWbx84cWxNKxBJzhYbLljYnIapM/QRHeXwowyXT46EfxoASYAqasDdqRP
JIquio3fL6k7XiXVxZNAWpSGH1JPwNxVYvCrvkYekf7PkIVcm6paHDphdugiR5UihJwRMOetYdxe
kWHkIo8y5CobgzicO2PUu9MourssAj4fH2/Bd0dizHoJrjnMnsXdxm53EwzyKkkZQUFy1m0TKFf7
cEiZcq7K5kX7pJt6molEh0zacpmhYffDqq28C+pQ+n4x5va6xkefdg7SiDs5UidRcZqVcyM0kY1M
zVl1ahm8zUU0rMIecITNu0ZMTiylef4HbEeov+ngy9FJkYFNj8hPRMNt0NkBy9tqf4WiScU72gAC
Mij7eO/JyTF3vrgwDiQKgoRegKnv0EKNDkGdgjTx6nCxCEkv0wGLo1pyZhaDV0S2juR8GfAZLfYk
NMHNtZPt2eCedn2V5u6AJOF5LjzADIHznZwGHfWH2kAOKYfz0R5xwNEjbdEvqVDhPGJgieKDunb6
mnIZJzxNzL5hkJWxN1L+psN9LYMkyap7C31XigCkqyUDvEkobbkcuQDsxV/3XIEd76TaTUPvtm1L
dzUwagforHTh+FC/JwAnbmvG3NMOLy7szdxBUVTXYDWe6ZcpM8l8g3H/LED2FOc7ad+97I6z6s2y
rsTnA6iwwSQcewcYAcXPVsWrFV8XUj9h28HokJlV97VJM8qceZQ8I80lSKtNjJbswLllPAACwBX2
y80IhrIB7GeJpsi6/Xm9wnpBVghoezdTu7fJglc63JI+bkF5h+qXVMzU8+QKhJKgij28slp0R4WU
jYFTpY9ww8YWN1lZZF67BRocL9hMPVKdPDv78nyPLkUHOg0vfS+sYb8c5U+M2BKI7cQV3+Kx04eI
Wu+J9Ap/cuHz3ExvebbV/WgeX9zgDw88DSHes2WAJK+lapr41Ps75xTvdAtMC1jlqyWXBh8/VZlH
NsLxTTG6oS+m6iAEwQWzPzGDnaG46pbzcpojXv3VCzOcCOQ0QPNohvEXfMo/TU3LuxXQ3bWp8joH
r56UaIwolsZFWf6QyfYrDtHIQro//KgoMqUkanUBVcXjPB7x830aj7k9n6q2yrXF59cReD7kVISS
+4+txn6ZXX9KRzfahHZlt2Gr0QeG5g5W7XFZVHsP504BzPOYnbjyKYJYvJg2XBpqusPa9mROKVgt
T9Cu/GLXGPL93N7ULQdqa0xM+KouXEDe4nMZ6QkP4r7o+WtA3XK1CZdANXN/Q/iGv7WVDt3k+kfT
72EkwCcrV7AgbH6NRnwDWkp7/JBwJl4DMPJIYEYQF1h74M/8NmtoliqYXPyqKwl/HIz2zzN0Yh9z
rs1elTtVoUV8VcZTfMiMoqdh1onKdDV3pG/PCUTgcv7enqL1sBgAawgb4WBiy3/CGr4ZGu5im72x
wY6XktS3LHYl7WpjjGTOv5wqe5nT9W3lMyZ7hkwQiz4xA7SdhPqAc4kXn/wIf4N5ec5LtnglW2Om
FsDmWRUSUevEDEeNi99aPsJJlye5oDB/x78IWLN3sOsKSF4skkTHsLP3vSk+Q6pFQBJnsrXJsY8d
C1KwJVsqSOjR+cIK4+I4dTMLtckTSwYdPXFCEdwXVZFP/MrByPhKIbezDqfznpyZaujhspEjK5cM
fuZfnbBHk4DxF6NnDrKZIWDUyEMkrufsntwpebXLLh2rqTHK2/LtMgf/++VIiFbdrk5GeHf6O7D1
cJcPAPfV/u9e0378Uu29b0OahmeHiV+mQ1bNQHmkMjYOhJrmmzHXbpj0Sz6KaRFJqMsbT3Lh34L8
FQ7Y6kB6z2kr924l25LZZnwFB8sFPa04GayeF1U2SuKsbNy3J+PQvUU6YNEiT785MSG3wPefRJw5
5sdgGV2oeK5oXmjVBwS38mUH6Gamdw4oTVCpDzuCZbY9CHRLvQHREtOH5Zr+iF8L/dcFjJTjsQey
kR4Qr8uIHCPv4lqfxAmKfUYIT35wggDCAGvbEmm9wM0rV79xJq+6SMC8ZbmFWZ69NOZbxH5xbhzu
s3jn9/MSiQdmMtoNH2IKrJ6HEJFwFrao4+CRSwMaO1LTETlwIyiZzUohKUEXUCYpdZijfL1L4qmk
JCxQ1JK6lW2C5TvfLUGpojOybRhME9n8sPow1pT85VZoBXCwbem+SAMFUPP0EvLvCPf406CB8Rrk
GdU76efV7S2f0F9Yp6FvsHKfT3DPQ3+pPyZRD4rG1asGAtyZMcHSLBaA9dtgNyhgn2iGRnzs1vxx
3/eBPz2OESuM8mYbDAioZ6mL2DPDDJA2gKKuGLGRg1YTXO6eh+Dy9mwRcrPz4cAa/ovn1lBGodqK
yay8tBDFpVG1RmTcq1O/Bbgo0oZYRUA4NF1tEVdJ/t3Jm+q2h1bE7Aqsl4KplJlfveu44O61Wkg9
GJDogaHu9xxVdG4gUHQXlmypuKFjY28e0FUbzv+c8RnlfEegD81YxNcyvfrM/m9TsAywyO4RedR1
esnFMWG7P55NyV8sCa2IF+ol/jYKUSRtZ0sXGF2ybkCtdtld2I/jj6u5iTduzowAUGujI4ZdMpJf
QSz1N6ObCbP4+2nRKITXoREuIr0GtjAUFFhJRtf2t9CJsyIWo7VDoVxqe05EYEefSXkc/A9eIiPO
ngZDVt7a8AokR7rSVTLIDcoz/mTCI0r7pJNGi6ZDc7IbFIY1Zg/6hPk1jGSufQMY3F5LziCk8Wva
8JaZQKrfTUly+VMqEmAZUuJHfrIZwDQYP53SZ4enIdD+Vi+u+yrm/RaI1wRG90lUdY9LXg0P2Bt9
lVMwuq2V3BBbFF/2BkPTVOzwteEa6ve2O1Xc5zEtUgfYDrFKN5nRBIeWuv3jXZPwlEtzKg4eptW3
xFPNOv50iPNm7U8dSqManyKT/OVcMcDl2XlH/NatBhVs5hDJ7dkiRTPvj2k19mz7/ZoI3CvgUMgr
/uL71nnVUK4McfherGVVbeqYyCy26xVb05P+4lpv1SjoMiyNfBDv7DXMwa/plVCGQuoRgcr86Tc+
trjsEGgT6yWK/bAf7PXdX8XUuNt2l4SYvvft38ZZuuPdcy7ATwF8X1gRRYM+773BsxlsBWqJDG5A
Z6nL3WE7aixVyL6nw5DPzN06tm0XQKbXPApfkTcWDXS2xS288Vkg1iZe79wTQugSAoNFeOHsgVku
B+6sm2Yb6AlOLkBO4wyMidi4ZLhfXoKZMp8Ca6uUEk1P1BvL2fWOElMg2BhcU3UYztCl7r4xBhDJ
bwaZi5Xz+9ST3vgTWUBWja+mZKZ46z8hrG2AKJFkSudp1LOIc9keON9P2Hm7e89uCRcB/+Ol0E7A
n5uSEhoA0F7eB4tvXnTMRCWMeAHoj3z8RgfPiczSYmT8Vm7U4Zgloa7EfMrJ1XA0ctsFMlsm1/cg
kV/sAv/4HKx42Ayz7iG1c9N1uErN/teFgy1hvsKx8EYDMeL+35jnS+MZgR+qEIzfyWTFKgXiHU8z
+py/lrHCA8PkPQhds7NrRWEP1Cp4kGkzWvEa2F/M9LN1nRvNIslH//1wtmO4vTuiXlXHDUrFZLkL
5JzzmR4GT8R59vb6JRuD9y6kdacQlfQwT7MqfenlwkLvn5EHKmxuvQiBOdCJUQtxphun8h19AMJG
x6gyAr7/ToXn4jS4JtxA9+XJzFACKLRyKlI2yyV6JAlK5+LXGX+ujIx6lJhm5dV8Q8S8oJ+IBmUV
Usjy2aZPPjUMwOs/DqiJ4hnLHXSs0zvhK+5NlIaGsFLQUugamgG5dMrbk25HH8bgz8Wp09eHwvcy
r+ZwuVDY7UHuzabUWip6q0irMoFTSMWzxVXcu+wy8HhYKJ4KRO9ovtd61hS1CmiOGWQcUUVMpI+H
rqDlmXrYlaXrV+Nc7pqb9+mV0SLf/NNKUCIBWRt1h58ybnJYzgUqI6NvBRxIzqEjT9zc13n41KsG
3hctd7cn6kHjtQSUyUGWLWurtOQD+JmJ6Q0gNVQqP1tTecyYcUA6O8iNGtq2MxiZwm7cKxmZCz7p
qpwFJ5dgDO4+gCeCHB8q8nf6tZl1TQvrxu5WrNTUU6AoScChYeVSyNi7zdCOyt6oFnO9v/F0oknJ
KvKpHTzRNrkpxyZ1naGpsAzYYLs3bwkdLoEXZ5RA8a+QNLDP5FhqvGj74O98gD7IDYYICCLS1bpA
oMOBqO+gypidng8IKV6umBb8IhmOQlzKPhZpQyN4Q5KMYDxJ/FB81Z6Xyw9zfG5K9t+Hkj6rre5k
yV9IEbkomBiGSR9277vCCuHIUfK5xEYlQIzZeaqP+OdUGFteX5UebReqNbudNgxDHnsS6KrQxonv
lD3y8EzlYr2L91+Bp+TMXr2dP94S2dD/SymoIjQXjSFvzi1pi36awx7npvklioggc19sKyvhWp6E
AH2NCNueLFcLvik1USX2dnhktU3YxYjZ7AS1264uGBwgdhweAnWrWfAFUYbrsVAPlZnFEG9218N1
Ph/94vHOGvNzFJjOkFYUsozN1G+YLS/PS8rAJwQmtNy2zudAhkXJ1NjWf2Nfa4H3aoIc0k9llnXl
OrGtAEGv1H1MoGFQWlCVk3dxRF/PmyF6vBnWg+wLU73kx3d4xEEgSezqtL+HojeV0VnLi2/t5XYO
7IgGXN6MLzJg2ZD76gnvxXygJz4ZpbKcqVVa6WiP5pjOBTfAxsIk/afXm9Yr5IMlckuhPCJPwcOW
vyPLLCOfcV7JTrTNjpkLzwBm3uneSFOHaO6DNhzlKZfRuUsqh5LMTMdmicyts22+7uCiVmNp6Uw+
oK+ERZEOFSZxXlaEG1HfOyyUg2QVgOFcGKzJA3PMsyAz3jnn5aGCbEF/GFpcV5nLojU+aEY2G+Lb
gjpi/S0TtaSCiKCAJhTYRMrjjhtHI6CuDYQIWbogbh9mhfDKzAjWjMFs207LJO5Lw2HTSxHXWahy
24QZC+OS3rx8dFFTbS8X8wWzeQb8+6x3ElEH55YQSysO8eH7wTuib9exoXej2QitNYKTAB73yl1h
+OvHMxdZe4WtnMiJmSQ5x8NBLwZ6RyFRLuaZDn7wLcS9eYjPDjQ7nWZoHTI//WfGMBW4E0eqFZyd
mYLcQpvR+ORI32ym1dt+Fk6vchIjgO+8iGBYv2W+nhdZ2M9jajdBILXj2qvBIIhI6ju9c6pc1Bwv
c5kMbjZ3r+OCcnx3gihGa8xyFZld8906qXgYKjolPOjlvmE4sLZpx7kDgzTyzIjr2E1Pq8cZxK8n
UZK8Xu2DJRZNH2ZS2drC0QVNw6c33cYujTreVMWXd1IPZCqgBqYtEdJE3VCHtPe1d1/8IDeD4WQC
rZt/29NxCeh32lze3hFHrOF+4domAL8aoNL+hOe9FRChdq5txwDVVjVdTUhZSvFoXJ//J2JSrgCy
5AOlA/NVnbdIf4br0y8QIXTVSR2n29HEzqEatrr2V0xWwRFRKmQsQXE1BXeVbjybboYDhDjwcp1B
vAmtX1I/CKZ1RqgdXz/onkpgephzVZbCXxM27+PODN40jzjEQEERg7jSWAX4whL0cX6JYmLpnWhP
8+nuvniu7H30HFdpFYnc04OgcH6gQoObCJ2ltVrF6EFlvrzrVrI4G4o5CbeLKBsGGgZOTpnJj4Fm
Z8ylL3aC4is1fYqHQfVD+DP4prIv/DA59J3FB8t5tIokee8Dx3Y2P6Ts635RpBAnhVK0nqJZhJgR
iELIaxWiBFb15Uh8EAeT2VqCVrCZBgPWLft9V4M2jbDxhAJBEMFctaoQqs5w+YGLFBZStTO8sP98
tc9/Idvr/Nw4L+o8iwZ7jB+N32qKvq7h/QJMypJbSmQkS2HkM0o59UqMwtXng+4HkxHqYoOpX4gm
HlJGm5OgsXDS3jymfX2mfl/IFUBR4wxVdeldBORlBpTAhksBuahhP7XYVtE17LMlMnvIGlpyTO8Y
ufChlQDc3vYf2ZVeYyQgfdo3GdiXuOR/tn76wn6vrmcOyhG78CH/hsyMVx/rLkHpYd2RWmATIYe+
+wnjeW01Wg8gmh8U7FncrHnwDUJZ8DSC5F1E4IHhRnl6zoUC+DK8RUR39glCLGP7/ZkMskbdGVF6
zs4ZGlDTCDvNExfbeu7kp+kR8a2XEvK1VISxkypCwkPdxqgKJvAVkc0DyWBtJy62pffFShkeZZWr
xdMLv2yb3QA1IFp17ONZiZoimyeOJxgYyRza8hQwWxh1xG6B+tAL949gQUMoQUZvy1GbChb158jK
38ulowxBAwsdFmbXbpPn2rbhQ7IsdFWNEGBvCBE13WZRIvJIbkUbPipRmXZTTrr+axcPjfoZ12vv
AAz0y63SkWK+LzZJU4VEILAnV0W0/v/cQxLeD2tE1fmP6IjKVX+Ssryyv/BzeDfVVSNuFtKyTXDc
LdDJOBl2uP7xX9oeS0MIU/41aQk8gmt4eupK+cHgWgcGIWFdDaU6yyccT1ec/EIClg1UFNGwKBot
TIh3skSZpTiVcKQ3LBZaC90X70W22GnRB1ZWC+kHZ5/zqYywbz28OKB5lgtDBRPZ/vnSdBkSIdvR
/uoDYDupSUjRIHg8dWbZ9IdrTL9gFXejV9ZQB7yIs4PhcTEiC8GnnAgmd7JrNfxCfyHUnnPekE8N
DcDKaNTWeVp0tIpQI2f7ycbnZjVniXhEJRsZVvEZEbayJw5YS4m9Z+UR3Zsf2uL9xVPeG7/Pwxxg
kNjYAEWlC3dNKPC8gXqOdCOtgUyc5TXKL2mKlGx1+18i0L/Dwb8pWiciEqMoDMj/DcXwZwYn93wX
6Zr4ACtEIkc2xaq0A7FRvUC3WBevSPcHPS22IhOPRIq/1htg+i+tamjTScZwZM+K5U4ZzHO4p0rB
MsicUuuhUlj44DWQUxM19Hj1xN238GETL5fyzc2FE1ntC5t+ibPZ+4ixfPBPhJP/+CZXr03hjBGZ
w8nw+hLYMxPTs9HndNTet/FRMRz1ywQ78N1DAQ1Vj3ORtYSNGNXaHtzjwP92yoQGIwYZ4eYevhSd
m01rM6/hX1Sq6j6apXQurEVNp8XnxV0rr87RQ2qf5/idElN3l5xe9XEMdqgIiMVkvdiatN8lLsgF
sNDcU/TET41QpzXYg06HzpUPoQJURpFzsSSxBtesF9VgMk4kP0HU1pwQT7kE1jkAN6OT3NsRYp3Z
7b3nHKm8myfJvtvkDtaCCSzUT4TvKwu2svCao/xj8AFAQVF/ZlhhVd6xi5W87+JkcTP9I0ksQqQ8
ijzsl4KqdOXLV3VL+CGi4rBxqr6+06yiC3DHUps9qsP4u66+/zK/wqkdYFbj4MB2GDPlkpcBKMUh
Qb6gYtOparuHQ9Yi1Ya/Z/scQ96kuJPp2Zw1ZVBSg4MLnt4lMi4crFsCcqtfseaNjvUOeR4qf6Cs
yX3hFRmBbjKuzZiTCrmB5jF/M0WpSQPic5aSulXayKB6nxzh4s9DKnwVkSvidSVkBJuJEjp/WaYA
bJ67MGQvFTW6YUrfl3g6tut4okHbR6l51FtYrTioK5GufbBXtxeRAaDFtNtaKPgj388pluqsAKbq
M9dHn0TI9AGbiR3klAA1lZ8lg4I9THS7kWGwhwKzCTbS43Kg2ZgtPFA7Dx8q9SbTjWDf0xPLxDIZ
3LS65Po/LS/BlRvoiO7HdPvXVPajyyQsbbLOLG4hFzKax2BK4mWUyoNzmvSxkz4TjS9gIDscwMke
j11AFIkm34cSZ/Vt/aGCIoOpfRRyOIY7KBUf+CV6DL33Rte+9dN0Y2sE0g4w59Dg+4UgdGQMMUwE
uWXf6YF1CPln8rbj1fZIPDtCpKHnfhy0AnMhyLA2NVuFlVdJdNvcfguc+5RNZF+asBVgQ8UqA4BB
jK9LrlDRWh/YYFvZ9dC2bPbXycFQhtP5kKZchQTPyjfV6LepyMt9Oyyg+FsIULDjU1X4EwrIPbKS
IHu7GCQ1OcVk9vFXK3Ggk07zwkvK5rEGLM4rrEovFueM3rtcu0BAF4QfpHd8/ENe8SDaBdKKB22a
Tpw+wRjPz+gb3xWktK/0j7rBqk6mQSloLW6nCPDr97NDcpsFrDb69vKHJLAzHtir0TivLWvKtq1V
Oow7i2xX7GlDrEf+hHhF00nluvtK7DWHLFHbiOALiWwlzXRH5odEcxaVGWe/63PIAAH6OSNrjPmp
CmalzPShLEjLrYR75aIq3dAe5WsaQXCSe7SM/Sqoe4sH54qyn5L7X32FZ/VJBDH8ZjYPuKU8KWHD
A9b77Am10QrkJIDHN61wsoeQQ6GadgC7/sgLvB9gNZIYb273xbYW7toyQH0oyJgOLrTM+8+T+p0H
XWmzbftdbnhmwbmjI+tLw5SQW9uhX7ZkeJBn9kAupv8E0e2knB1tcNDxsi+V2tj/azUKh3asFzza
Vy4RLkQu/BIlzMJpSjK8XaKh+a9aHz7D+cR0DTiPq9NrPJWQsl8f7pf7MT/LiHnLBLU8IxDz7bD/
+jQ3d/fjeEhpKbcqXLCChW0dqY+jZssG6gdf2O7+ZUa/vbHaWkf1iXJEKibcysX3bDMq7pIP4Zom
bueHwPrmRvLpAaDrL6g/VcT+HYkfBWOl2u1OVxh16Abiq2FVnhXtLqi1hiUNQOEoOXWchc7Vbb6I
S253mLUlAKh5Nzra4AcDUIr3hVbpa6lWX5e0eCsX+eCmToV+Ofp1I/0HcK7/lQ7QpZXLyz6hLdXr
ha49khIGiALWErU69KYSrvXhE/gEdf0e6Nr/H0lojyYuwJr1P7vHvDAGjT+BbOdnErgd68y1S0VA
LNGY2y8OU0gpGL+VThgprdlYR7nl8rKImzl+/lM6uvxUeRN+0v6WDJApvFVt/vIeSUIEwA2zRN3D
v9jPXgXZo2Zs0b16F4XePy5+9wO0fW13IVFESVCSGl9Y9KIhYg2JBsccNIoGxGgAlamdztd9vTsA
d518Q+tgs9qPNYkpTL9AGyT8P5wHup1Sh1HlCwYcMLPuH+FuV6PWnY3xPsKS6HkJTlgMQE12dJl/
9CW7jP2TmUriYnLkIIfdVyblRtm3xTFWpHUFZUyl3LoYus47z6moqddiN4cT2mThAj6aMmQ2AHBq
ylyKWgCAY+XdtULzz1YSGxkmVXnCg6W4P8cTiKeYpgIDKVJ889xffQn7zUfiiqkotT4uZwOpNpoX
AWqTMZ7WWlV4kjtWxNJLniyoc6hU3cgkZ7FtN9lUGAVIRBCGTMO6XtgzOOrlJpM25wrqbfEOco5j
vJl9VfWq62Qzrr0wBfMMtppn2Ki+B7Grc7Z1rBUZP371/Lqf8S19tHPfPWimoMQf9HFeNnbxgaom
VdEVaIfMFtQWuGAyS10eWwNmQg9c8cK8wXAmyke5yFr/haiXIYPP0KTU+lvIu7O65e9yAkzpHex1
3oH9u7jbqF2c/AvJHw5bShmGMLNj/Sms0w8PjjtXWtct93iiwJRHhFPV6SRT1ol6uEwY9zt2xyd4
C400vESLCYtGwvDzLgpi0iLSj0uPMcdKI1EIWTA72mAUcUK7yu4q6XCQyvj5k7zux6OcsdgkV1FV
qSHy9aPXKE1OL9Konqocxg1ZcMmcY/KGTKyiyFFmVfDir8KdkfSyytkkYFBHkPuKE80pKKItKv+a
IZ/+20weeY428RJu55trcpaxtbw8cl8/cGOR3APlmxailZQQRvPCASyxEPZP1O8FKZHoGwujLcvU
g+kIX2oQNQAvnx5A3cSCOGnW5oVuDzDF1EM6/YYT5bljvEKupzlMRWe2QliT9UqEQl9yPbtvn4cO
4TKnUf5BVaf/ZzjiP6StTL/hkXhiAfte7sXe4J7vurqzLqM07BoqNxAfXrwmayRZi0tHQnDDHAXi
/8mY6YhdIz0VB5jtNjaXQR3C81oaOMmKewMHWSAbiWkSG4JcfkEpwhP5N1OTio8ONbLYVdBDSEee
9hSBClGu4H5EoDooUCreEhOTSE/f0Nab5UIrDoLbK/kUDKfpPPMWO86t8KtXx2A+fjGX1KYa0XN3
oJ3kQ6dZanfi1dky7wb1m7Mn8AcJYq118Cdq+mU5XmLvrsXP6LGcZ3NrTPDs4KwFNnVytFQyMkgv
seIWWhFvs5Bmr3mn/QiT4Mp3agPvi4Va8reatZyg+o+z4rpnYm0jysYeWcM6luEPSyRq4NUhbgOs
grOtumPcyvmOGdLjirMMIo+wXz0k8EDW8Nb3K8X1Jy0tjATxIl7N07nRdTJn5imKBWq3nwMa5mFx
N4th09TahYIAtLvZyVvtlT6hG4pTkCpTQlYFbl72qtf5p801bkWlV5qJ39uQSNQySa5T6gUMiQLg
wp3zlgwvCTTGvZM4HcoXFD52cGSTdebNEGwe9R9ID9SZqFh6dlWbVbhtZ0nv1Im2+CadRCjQFy24
V7pO0oIFXI4vL5QJBgyVnKQz8SvKbUqz7f4KUBk6isSA29DqlLndPWOIe1PlfD/KO41pHEGeRJF4
tH/aRO3Br3PB+Qu2v5ur3cJEFRYR23XiWS/rQaObk7m9lLT0RkhtxtXiakcQ8WquEj8JXXbI8T4b
gC7P3b27KdwMBrwoMlqUkqZmBLq8pL6OeZCjYiLqhUFWRMxNmutw18P+6QiYAN8F6Bcrv+a1+Jp7
bez0SUdh0BSw8n7C+dbnV97GD4Sgn0+yhWJWYtxwR++WKUWyhS932LR4f6l8ytIYozINYErhtqOZ
J5Zg6Ie9oks2knKPnTm+o/S/RElFcXg86E8rEKQXRbayI6MVjxtWUPv6MfuXYEW2ZHr1JonerFEW
qc78QPG6wcMgwUpXX5kOf/KYclm3mX1Ssw2bKOU3AxfnXbT9vIaJ+BsX8bORoNImiyNpJWvv9HUY
vQLQ0jaWSaofxxA5A0Ua/T0uJLJpufLpjBZFHx3zTWxDigemVB85/WXprM0DuDKU4nvI77c9zaR1
BZAUwZvTqOmt0FhQ9LavL0o6zSdjIloDoEKXCCPaOk8hYXjiigtjQcwWS2a8sqkTnh+b8bI9EseQ
aqI+/D+A2wDVO5qGdZpo4iazhin/D2kk6kayhQZV1XQ3zkfLd6Dsf8xlbaNCbcCozD5MJaV+kOkH
o86AUxveAfRyQ/G5lfJVOGFEGcfrqM5vypkCSLvXaK7yA4rm3oiChB/gjI/5sSxWYothHBhCLJ7v
hBnrkkxwRV6Y+sBIKC37H+CfzXNueGuyAGKyMLXHtC7CTW0x8YHTDQm86LkFlFxt2LkINjFhGXWZ
G2CPym5b+2mDp1SEbFw/KPba5DRJGEeYyq31gJOzChxIcvouUJ8OYFCuIYL9LkcbzU3VLL/mZrgD
hXoVW73Lb4/G8CZylC/1n9GMskrzVCq6cVLyB0pNbTdVpe08d4W8t55JyFPtn1D2ZKLobED0mDO9
q7G81tYIPFRHKpEaZHz8Uylex19/GzyvmO5EqZJ2ZWDuFVILLc7wiKI4vdMwUgnALvp/hOcnFtKY
j8NF4/PBIbkBcrORSBqBg60qFhCwAoipEX+HR5bvW08FHQH9h+i0WYEKeRGU8S7umbHm1EoLpmEI
7X6VxFRaa66zLlH6kmpfcHgAmvEVys6LxOUMh/jFWC2GL6ftL0ZVt7Wj0JaqMXj7C8zakh0MhVlG
s6uvOMJ2LW5yYxgnCv+5YtoME8OjOjHjSCPlEpF3J+2PZyea/6PozzstpwwenmPLOgMamDJp7EMX
/vyb4J1xKpsGUI7XC2ferJSBrlCzNUuLKBfCaOkQjiwEU49UzDpmENp1dcchMtboCVX3jsxkuOXE
1Br/OtYWzBfzin2QaplkPg1t2Bmxo3hkv0dbj0zUnsTABdLbyMcyT0BgB223H9Jz34uUboJbP95e
kwnMv8IqXzOu3iLUx37tcQ9GK9KWh9FnTWvedVaQ7werJvM7EjqA+kBAALy87j7R8Syq7C5Jf5P0
S6NEKASVwevyh/usv3WiuT6I0J5fQ48ftTy4qrp8CRjrV8m63u0s/Zb5SjE8+vvSkSMKjKAzO/XJ
a+xMxIhBlH3ZhX9ADRZj1BHIebEG9TyveIi/p0VrFAO5k4ADqON4PP+xgBc4COqQLaUhCea2FpAW
CwPzD0+cCeo7Od0SN61WoCEzEO3L3rztJ+pGOg8k2rFeeLmce1LormKMqO1PSMpN37sqd01NJ+wy
LFu7nugs6kDHYqTMcPva5NVcEnwpjmT7bXL5v6bhe+/w63EfLLn0iuGYjWN3+dRgSmlyqlRPYrDW
1/vosV9NRMdvjYVIFpsYhElTphbmf9EGu15bxjBy49PlmL7u1XNYSigyDmvFfASu/3gxJdceGTkf
bzpPkRIgAH7NpYuLrj+UUew4j7QgFMzxykQ8/EO5+SRPyNlo3ZwnAE7MHCASygj0O7HpKBtk4mfW
jamr5fjURkcXPEpwhTbBcC9qi72iMdqcP2Cn4y1NH7gvqNDijAPwkUZUG3FzGjdOnFvQ/wDakQl/
A/t8NgYOSrJ+9LO7gkNSlKO/bT7ngVu5zCDdYz4bUIbxzoGSLWgKfleZfi7bCQ6Z6idbW+GG/WDE
9DYBr9XuypKxyXGrFZuVxQB9tD9bI5HnNgDMHmm1hPug4T8WFnyjk0crYwOPditogwzAZ0tmCcEO
CiZSC3SU8bVXJIw93TkVYkvj+xC53omxzHblPfH7YV1eqZZWABb7JUm6IVolXY8hfdhRaS8BGyza
4PDEZanmFSlPw6oOSs+S+9GfzRB6nOgjgPMUgDpp/iWRiK6juKHFpjZcc3OBNuxYefzhsNYmgMEk
tzsSwyHAINjdE9NOZbLIvVNlNKjEiHOanKzWjqlEiLR9YMyRQZRu6PzGL2fWnD4uDxPf05bvu3HP
PNzMwhIJDHf35zMcTKZirgpda5QoswmoPM+b+JwwANTMZbLmrbmY7d4BumWDxdnGYmEh96x7HRwf
cMZD/Hv30nJT8iEKeRdc2vKh16quOcasMYmpxXGrFwfMd2sCTZt/yYZsjRtkL4K9RdWCz9GpuG9E
3FxBkx6HQjY5fkspQTG1y9P/USqLTvw6bhNeus8XVTorGUewgsZkAjbjk+I2g3K+OJDfhwQwfDwh
zuamd6rjkmpxv5ieP+EcimdFuPPNZfHwrc+J40QriN08FfnXbthPUREjuqrik4db8pJwgMaScu8u
2mmNg6YJ+54q+CKzq48XLqu/nNSVyxjC8emI1OM1qzG68SZnx7tZetW0MgOEFdV3rVDR0/xwGCgb
e3GwJbQluSPJYo5+9SK/G2zfjrG1UH6g/w3so8ETV3v59+FLwxYbp8ygHEooXDWLgceLhcrREcrN
/BmCVWdyB5IRSGL5LpJ2gSys/oz0Dn2ShX0ItMCMML9feOigCb2WL9r0F1777W3lnMFafvYEFagF
768G9jAVf/VFcmUBpa7uqT/Gyjq2PFvDlO8cjlIveexoAjLvTfM1Xlc2Yzvp2l5beBuLLEQtjMPB
h4KUDpeIAwBKwORuXiEOyH6KCNUmZJ5ckU9A1IYOOjurTk3VtMKElaszk3WdiyiPvkmV7Z9tLJY3
4Uz2cXA9xSacoJNML9GxNOvLhr9Q7QcGzP9r02DZebzv2ujHd/NkqOzXcNQQAwvxkrrMBwR5UcZ1
mmX6rtVenpHjb6Jgk1l6di6BoftN5qYAoa+8X6HS8Ozvdv5DhchqBdRRSIhipeSbbc7I6PvZoHXk
p0J8tdg3aPHmY2ou9Epj506+TTOgT0JzNmOQlHtnj7NXYuVMGZjFtDV1D7eM/wIlVlyjwyaxWjDf
VjS9H5m/bmSa2mCNMfdPW7IT3eBHBQ2i87RnaUT66SjCl5dsmR1JTV1NF5yZz45qFcQTUF24BPPG
VEGhdV6j+fciDvTWohda49qcsSUW3DPhTZfp31fwduutf0Kg/wvp07n3X96/GKMKLZ0NiWE1ESGL
+U4NgLdPV788nZ6YwpMRLUoxrr825necgbZtnKELCU/CPYFtn9Ks4T98sOr91p+HDzp8rzdsev+k
KE1lUv1JUEDCNONWaouUiSGzyHKgEh6OhOiDy1+Y9QLwruCKlXE3kvzXpEWfrLf7Vr0zRf3V4s9J
uy8Uf9RAWKGrGhzm7/DF/p9X3N7UF5HFU44b62XDKyNTVVX0oc6SdVd33Jf/byRUu6jsMQiIwuXj
9W2emohcTGiIJOkO0mDPTsspcqvGaBO9uQjaUbVVtwpWvoZIQQET36428iYa60F/0rE8snL0gx90
Uk3MOeGLxyaxiEbWerPXYS+ujcEhO955g1UHslZDoQZQsvVkhvwzweOlBDRycR37jy0N1Ew5Kuni
NJkB+5fYF9dSycE8YeGrKE/hKJCmsZCrIespEnmGGubeJCJJ6/60MWn3qMAcdpx1kbFFgnTQQhG8
bVW5GLWoCpsT3pv0T9JbE6n9+UcqWYdgjS/qDv7VFhXhRaati0FheooFOojqoAAkNzelCZkjktXv
O9U/Mtut4Lo60b4pPKcOGoDQYVQxn6TxXHirfZH3ACPa8giE/rl1OPrmKauk6LBA081xco4d3FAN
XGjX9bMgto7LQKeYpCsNTQO793Ue1A8TJv713KAzfXrXkjCiOS3x71D8jIu9XZAkhPPAbRK/f0hB
m8OzfXnwW48uZD68M5AokWhoF0QxWs1sW+OyV5e9HeDaDv7I/r1g3yuf20kzcd0nJOUvAxAJDJ8u
SL6mU24JXFJ2/ASiQFtPiryj9EPhTuMhDNrgS/2YwTSP5nwxyH/Eou4SQkMD65aPfmO3PJxinoHs
trF5gA8oA5kbp/HRk2jK+egeeBFU5K9/1mH+9mjnZ3B1VCzOC1ePKrmZGhSnaf8Q72dSVKXR3gFi
s+QhO18dirwNKzlzGxy3zaNihAyV12hBqrrj9n5SqT3D7dFbCl9RTi/r2jcgv6r4IDahRE9dHHOs
ZrTBRLdMAYoAIy4rjQ7ZiXwgm72eM7YRN9Zj1CvjxIPdkcgDQzLjGp/CfhHJtVd/ajdXmk68e/ye
ceS+gxybzwlEyv3IbMO14F4v0WhYG71bVudxrErRVQjygLXof1aYz7+50DNJ6SChdcvgr+Vc8AgM
e3cd53eVmJUPv4gz9L7Okwwy+Z0lDr1ds1Fwk3YSFmRvOWlktawwWD1bokfS7I1CPYrIWBAnw2Bw
5fsfiJ7peJi7FhU6EfAQeJ05kgvqdrd4wsctHvPQqX6hzUQ1DYLaKUKq7MrVIN2TuCjl5fDMVt8Q
adc5aAEy5dxuUUMc6U51olblMix7pej9n+BSatoLGyTD2w+S4UfWB5MqI6CKu3hWLwy33Wr6mwoV
BcXA7l0BOpqyNY5XJXfGhEaCaqo1mr3Un3FviJm/iYOzk/bl8UVwi8XYI14Ch14KD+vphyJLlbLc
fUug+c/wwTWJVy4WFaV+yutvTHfEzZNeaFUPwVi+bkYAwUjYnhlQboU2sAjF62kt7SlPmaUt+C1l
lcry8vRdwpPQEKEf/oui1SNv7vBoURvzS1yr9v94CbCapu43p9IjIooYDKvz3EhpBCr2nKT52jzA
YoDDXCiQJhrc5naizXaBqPoiOvH9HUhdx4QON/UHioNtbY9BkMeNG9yVdkjaaqPIPChsPf19qz/v
m56dm3MRfoA7xr/NSr+bcUTw9Hf4t0VpNCeA9rO1fykOwVzaFDLte4qBtE7iW8+WqgoKH8QLCkCU
AqbWijIaSzgZDpBjJAuSbtU5Uw4Wm1QJ6b8w1dPzB6pAnhveMWS30zXwZew0i/5vVApFeNg1pLtW
Bbd+JUjv81TPgjdaW8vWZ7x9Q1t0XdJW+Rh2yhBM3RtR3FiKkAcSmSR8YKLaF0Yh0Ff8NTTyb6eQ
UkoyE36OZCz86wApFkHDgwgdg/V9mZO8OnSjHHweJp8rUa2EHkiReYPgRyZMx6uZ5nzMzwdYqyBu
91HIaDa+DB9V9dtUCvKVHD+ftMO/HNEt1Y+475qGrjL1aPSzrQ5fCkiNN1Pz6jUScJXEcBgesPUz
A+ys5CEtt5NHLxt/1DnOsIuiqz+JnXm3fpBrV7eqU9VcdHVjUuAaEjtMK+4KMHFks9xkyTuK29TY
XvVx2gC6eXBU87Kqbi7B67vfnOzSTobhpvIgp94zkDE8LEHFbe04aSZjIUmQsz7w4RhbWu/DsOWy
Vw2CyOKMTzUSJeV92qS0MNyKrNZzrHdlC3Xg5MOWuFARdHVBkGKgz2Iy+FCpk+X05a2U9hLBGrpl
uh/zLhfwqid3+r1CjEKGfPvxZu/c3/zE5ZSUesCjRAF8EkujHi8siFReIMJ5RwX1ylZIMWZyVoBx
B0ty9EvZ9fecywtG7XrukR5jR9Jnbzu0o31eaqT+QGyUAcPyyT0SZZ9JO9PlU8FEWsOLDk1rp9F7
Swoe5KAeVgKh690wwJu54pjw3I2wjs9BZTi59ZI15miJ9dFRf/c950nWx9hh8EwM3FZOPb6dV35t
FywAOnTMtgC2gdz/JJPN8Tme1DPOLDIMrZd7kE3hgKMtx95KAtsUULWP1w8MU5WVSug3y2op2iM6
q+R80BL32lWGc58bKFciFhIOGJN8azUPQ7lnuBEitzXkSxhsR9466haln0wHHrx4UMqFQdbzXDYN
+XCbALu+4UPaOAtk0lGxxcwNZ5eP+HFyttOnmIH9utK0A3CmropXMcbUJag3Rvcd2AuGlNBzLPhW
fxVzPRGPcWdMZxCiEyLJxbVrtxdMLoHYqPTYFCxQKmQijYt3Bj5Wtk8sndhC/RmkV5jI93koymBa
9PvlDfB7dMFeOelNRrmARhKjvbhLu/QbFwjytYDLjGTlUWPI8k59GzGUGXZf3FrJBEqB1I0cnt1K
qUiBvn/eYOM8vnTRNNcD/22CDC1Y4vlZaBwHARJf0LX/yPczEyk4cbLD5Sy08c9EdFApuFhtT73C
GnRCS/W7mnCgndcR4CwgDpqjRhVAAVbjN7v1hktIzrm73clCXAN1FibdHz+/9TieKPJkq0ggwkq8
7U1U/ho7iFto0j0dlH8BVJOQ7uViSlpJemSiAyqZv74mLs8HAGAhC3SAjfpNMUp+LR7GYjjZr2BF
3eZNxzr5CVr2z9mgSdMtFZYy50R2nYZ1pxEQZakr+jSEECuyVSCReMAxNqGiUiiDpgWFZferJ9aG
t1WKSuQuQPgBj2BAB9TGKZHSEJGGM55HmqeNHjz5HhOVEie2diAblT/QxgtNg2Auemw2vUL6DY3l
fTkS58ZCA4877199WVwZHbxs0nL4gMcfBWiaJI41oefuBV+cpw9I0cRS6DmT0tfeReNPoLIU1MXC
6g+XXdaNp72ZQnRuK9npWZ2gojJVj3W5PLBSrNIxhVN4Eu6zOYKZQcQwAxOtwyeCkmlqpa9kojgE
YHVQllydsOSpAjyeOhtFGCtgoofanY3hbC4cARZwXsnxWcYXOnckRZp39bOvrt2P3Pw40bETl+Ym
jEyBv0EJQ8wuUI7jaAn760szcC8lw3kqfOQrCON0Wh8UBNeCEfZ1bSMlHfRVT60diZVnFCWwH2d2
sVJWI2tjJRDK/MizDoczPZUJ4I1NV8Cq8MpbAn12RxFZBfqqnwDL0NXHnTdvbu2ulg1DeL+B+lmv
EI47aM8K3BZJYpoTsnQWb15kYzsjGYpBh41Z7e7Tp8Fd3c6/7qk6annwHIlcMVOSqEfmrijjPx7R
8wBUtSP76tC7Plbddy9ksB8vX0AI3FZ0qx6DDKfoeYRtBnJKWSTJ7eIMBtrV64Ku74yUf7Fv9lLi
bowJvVNuYZ/Uv45hrdcL7J3tI0RwzwcJ2WXOXyD6FnLW5tIWuCBsTo9R45leeKQD6Q9bP/DHCGVU
xK5zxP+/Kof/jNv+DCuQP8+iP3+Qc4RQnMY7Uhn9rHjcD6i0kGOulT47O7sDxxd96lw3Hgoh0B2N
LLKMbVaUhEDpHOB4LiNjUlng7eSfTDlu1E1FyUyJ0BqQJmbm7OsT2UKPD3Npmpgpag7AeYIoVoFs
kU2zg/Jia0c8eo10wFKXBUjf0TgUfzoRseYBhmhdJ1DXB40JxKejrXlObHFk0gRfOKzSlaInN11H
NEWQff7yeVuAptOe6hw2qosQ7ksx2HgqgjEEBInjJSc268U3WJ/GbkzS07DqBnz0NTO+eUsmUW/Q
j1GVl49dZy5W6rlXXYrfAmrtwiKuFIX67NuMifFbzKbfXT1tMdh4sFgfdHssxausxi2a2HdC2KB4
db9lepHQsI0kmADERZUdfvgxh2tQT7O6nrMLrrzTINhzlgqoa2e2ANC8Xub5Vnl+7Z9erpTWIl+k
YuwyDm6Oaviztus22rz3Ds5/IIJc8xLEly9F/S//eR2+5tnL5xX0U4UV/pkcjwOwEAXIEMcD4xs6
9cZpu+1p7SpH3v/Q5l08f32K+0rAYnMrDVWbv2S58RJK5ejYFBG/fxVH+O9cxHEA7N2GKQUlJSNE
vUbA6iWy8hG/ZtQKFU0PMoVH/wPAcXIkOUIFwcSSRprNycGjKkV5gpJ/YmRVVrbMQxdr/6sUKL7q
pIVHx3dtQA0UyT/jo4+gbutKL8flzNw2k2q8uYORtz8b6vPxQJ5KEXom7v3s9TvsF2LoEVaBJR4m
jOhIRn+7HeQRDHV1jy5XEj+HvEZVZ3UokSfWUZ5oObjwmaxayX49snWHFDBMH4wzBqDrM6Cjukd8
KGuowYuzU/wFFqT0UIC36EWArfH6wYqypKt1iBm2FHL+7H2mREqIzc8yDIvDrZgNPQSoMx+u3HHG
EyWBV4IJQO5cXbUuhgx9e7woTjkaDucmcDTIvQ5GzT/5szxbZ9nAa9deSHMSBzPrYQAqu86oa5ub
tNX/VW/eIsHpR3U2FX/a0tNtFV26lURkRl3Z8WLb88j5OmZIwhsnYQifUAOzpgFee15Vj54/m5+j
UM+jtngEyyIfJTBHqaN5nA644vBsH7jirHqNEbo/yMDBhTRG7+VlTsWgPYyFN0UGWKJPFxbBAdee
TMv7Yr8pvowsNcdPna9ADlSrSDv230SZbcngSTSdsb8kUXnojWuAXWxGOq5C0IE29g/xZbF0Q8mq
2sWGPIwBUmslOFftuQrLSl12ErngmX4pQYdI2Iq8DL/gi1XwHqPwSxHtkoV/ubsxdW5/hD6gabO2
/xcIJTaQT1eNNxeuL20cYeiTIlD3DOl6L7LQyinALpMitICmR67KU/qS/ub8kPmfzPgDEpA4R8fl
QESYT/iD4tnmBBp43pMi8brfchqhTVlpd7SO1n/77sppK/JzMIAOYTBPzkMA9/KJH/t38jZO4g8S
hFFrLPMriEfu7dcfboYJKh4PkM7otf4vaavkKZyr2uTet1Zxe4z2kXGaRKOp+Jx/64JzXNttRxpU
GTPR5RVWbUZVq34EYZ4QW1hQ7h9E/v0jiEUy5vJ7oULG/O2Oh9dD425DJzJknEZVIBOOHDyRl9sP
BgJZWokcEMCCOcrb6t7UwO9awRZma/Nhv0tlW9Gm/pmFXFVYtzbQ6o64rLC2Dt6252hc/lcG/ESt
uFYK653gIUoZMUPQWuzSiTQ6nWHQ7Fl9TaAP5Vlnu6fB+k0Bh7VtHj7VIUlHgqpsiJViDvSiuQpI
EiI6RXcpQ/zQ/iTvzS8u0/ydjXwavtT82fCjND6MkxwCyt3r8EvXgP6ciVcBW/TG+7OmYXFzcHxr
p0Y4xYWX1LsryT7hyKhlrVXUP3AHY7O+JDB2AgO0f8OrWQyuzNjTtKVc6F2CTJOmLi0omecI8bNv
vZmbPdO3HwR9bKF4TZGWpgFAG6YWXBODVzqBAAKGw+ZcMvOtpWsIAHKHPZ37IykuLceiSItOskjZ
yiAG+e2GLB/ALggvUITLr3xfS6Bx6U4LBxO5wJNBB8lazLmDAugLuMydf6nIMuTjZ8zUyhqXJAH9
2ql9LAvbgDSHURwb6T+vHeVFowgw+rB2XbMaCIoxn6YKrE6pJPdUCWfq+ZkXWOpIXqWy+bpAxtRg
I1w9sXBV6s7bwMcWBHRSBAk+HlWmFMu6ScfWS7rVVbv91pxnwuiG0hviFG3FrAD1QzvTuoEGSGZ7
nrLeihbNmfilL3dU31XgtTsnYE60mje9GrgVhfwHQU0yQElgbk+644Pg0Cjau9IryKfGMMhzIjnH
sv3Zb4lTdEn06Z7IhKuWsaV6kZ2AC9fBQqhTG8ERLz4Xk+t2FN4Bqt6r8ogYwKGLQsv4LaEFXIl8
Vci9CCauIg32yr3LU3rH8pRDxbRCE5yOpKkds1nLFPI4v2oP8URrw9v31/sjcchhNYjqdevmTbQL
s2SNsS2pH3ZzaS+UWpyRiMINbGbt9RyT+2OMQIxoPJFLIF+W6XZo7GGOKwcKC8/T00n3+YaNXA8B
vsC07tpqcsZoVWGx9DxG5lSnWPW01lqOIBEWPg9pUq/voj4hVL25qNZj60lF7g4aK9OVQs7cYlwV
Ew3/jpKMet6xDkfiXkRssoPHryYjYgEdDZAvUcxLYD89t3VCSfSxtLuTxqX/yUyV4A+SzHSgk1aq
ZqvHJkQtpUj1ctmT+NwP7YSFVrqVIgrOi3xZAZr9hhTfAydZgbVX1h8a3gUDnzlwRspQbOTHQYFu
pjBkOBkqW7RqKS4Yrw4Es3sPJjjUM2X3fhWSiMUqdhEO1C/TWSB1zP/mzJ00G1Ve/9QXz0ThYRb6
cmgZhjaX1SX6KygrnjEed6Q9gsalkVSW0wrF3Gsyxf70gMUGp3OmI2KU6J6AjIncB0p+Eg0ZbZMy
84epFUV2dXY0BUHEfUSrb0DKJNlRf1OWhlC7vKO/rHMSP27sZOF9zwOubMolTga0CQPIK3xLQwkV
LN68u+EFkdYOXP1GkImBJU9GnhotdVKbcT5VBT7H+pU7YDWj34tdjt6ITpIqyy6TpT4BglEXbSIr
Is9XH1NDLNqRVnR/brsxKkEMd8asYCP93cXi9JBybEuC82cOpcl0RNcOW1ESW2qksnxZJuFUAP7K
pV1oxkCUmGEtcajIdQNlbcUXPzWF+Izb/9M08GZT2HcAjYTisrbdin5lGhKLAwfdYdSvYGcVID+H
dPReP1sPq3mWA+CVqFZQr6Wpk0mefXnskpZqqDzH8Vu8s+/D2nfemYpps4bNIAzp4CCehqZiv93y
A9nJ82oChWVou+T55948SiS052LAfitJiypp2Q2XWybGG2/J1s+x17CP0NRepriwaZWlLrYi9+to
7PQxuY9CQJaIs/s659tgMNbtzOM5oBnOFcN02WS5EO4eCiS9LlVEf7hBf5HU2SsKfoMK7h979711
bb/Q5dZr5tvnGwVhqU8DidG+CkfxW365G5qQWztU0vqKgsj+yBNVmweyV3kwR3Qi10tkqZ8t+pTl
wqu7Ro7GEHOs47v6JVMbpnE5ECTCPXbma7Uj95Bp5xe0PBtMRUVA3fxyMuz388FDayLj9N5CdmM+
6eLeU8JzfhgVioRsaQMFFCMAPhgu5Tbo8173ooOzK8YJBUKQVckQJO+Ha7Txvz/Nl4UtRBjLDGyf
C09hZ4vsuJ/DNjEuV+FfzKdeNcalWkXcBoeGKlKL/ZNehESVzeNT66vPfTm99jnyc6vNhbEReZDx
EPLUqzUnp7cuqYv5WSHYWG4PpPltwE7NW6bUTqUxjk/dIU2qz7AxOkLXu5monpQU80So4G/zv6lQ
Xw6tLtzKN2pctEHILzPBysHW4cfP2AocbUsMK9Aj01LAxOeJssqicU4J4Sq2q9ARtVcvcCQHaPPX
XANHwAZj2jY4DctzsKlYuuXI0nEX0c5lOu2sl1kdx/qxahbJtWx0q4zzX3czn+Hyaacv/aGF/ry8
xHcskFQWYrrGi/Wsd3TbEvcFxXMEeBDB3yGKdp6SJfpHD82o5vYHT7u0DaLjFArfxsDlTGtRpH6d
yDLH9Aq07B9Lb3Tdy6dsaPFLqVD+FfLQCt3+/TPQPgTiHkQS+J+LrBBs3CmJSLgZGDEoPdFN4LJD
g6fl7BfVH1DQAg2aJfNHR9e4x4sUOjhnlMjewHvVyEUQmCifzaiatIYInbDPrfIBslK4sHQ52U/C
FR7AE7CxaaxhNKHMs3mjND3fjWShrerB/1/ZpmKuwXXcQMYHkCdPAGc2Sh10v1RiEW/rNOPxkcSM
6WlPk2tamcOF3jbYBCVJafYUczWcUgJLiRaq83NzG0UXaQDtusrP/B8Tx0V+w4+y9XCcyvV8A6qL
8d+4rw1sag785Bxxh08lkX+4FlKaYdPSvDa+PyeoAoNSFbMw62dN2EmVqVdjp0tAnLuvX8EdG9eh
0KvBohwiei4XIvYU0v+co/GoVaz5wFVKdwLF5lEa7jZZuwe4Y7cS1YkF8YE05myCHYNAikFnGuVU
7jxQ4Q+QOyOQpt3KkPXRozxxcDQh1GFkt6tCTVb1ziqAqss4x0YfpZbV+nyip/mQSSII04+ffrS8
+fg2S15Uk2rcms1R81lUykWY3BSb4ZTF0UDYWNsMEunYmWd/KVY1WccsnpRipgjbNGFC+wGrgf5/
TBoib3ugu9f5mWh2MQJFwfTtBuPzlN2FUa17zo0jWPn+2zjHaGUrP0JfX+ZlF9G3cOJLwav2S0xq
BnAQSCY5EP+OOqKdLyb0O1dA8TfDHZ4g0S57yCzxWYG8m9O5vdN1bWyCQkVSXlJEt/PMo4HC9FQP
1v67sFhckEjL6hn6O2TUvdoPKe8W2uZy7QV1Mwn+PhcqpxBn2Fn89cdzpUISc9SrJBCRLLpPFhzg
th1edrtVjzzMRCfTj60+g0f08drWObGVNBLTs1hXyyhSKDyYrM/gWJj6tlGNAoLW914rrdN5n+uz
GDeJkDrgJvJJqtJQ8vAdRAWWnimb+zQ4Qj9x160JMjie605ouxQufv5HE4As2nrWyCJq1S1JOV4a
O7VTyCINnH3ooMjEFbEEpQe49IF+1LvedGGfDTdwLHOdcF/rWtH2KuOZSO6H2ZF43ucMpLptDcYL
nU1vFbIP52HyWeHVWu2wqH2foKXV6dk7PAWqhI4aaSuJJUlc21LLjn+ezwjV/PzBLAvAIj8In+sh
iXldK/dS8F/pEcK3fq/zKRZmXCdqNupyd6f3GCZNlt07gESg5TlUrVIUj6KaN4p8wxxulTgeOf94
5JuEUB5Fb4yeYXM1vPGeeuRvfzpHKAkdtLtgBh9l/8Q8QePR+Lmqu3mhfa1v1agb0WgiG3ITJYqk
rD8PFRTts+i/JTA9St8PCniCObXgrXh5VzyyKkkhOmR3fOiOSnrGyV6GE+lRP9EZ+vVEiJdCXUc+
yYW/Ss0iqVHmX46wviMCRvvMn9EAlucFC+lYPP5scqe3AF5dIMlyInjFU/9ClOFhuYp9uM/MGu/G
Z5PksSFx76QVX8a4lZ3uXj5ITj/bH05K8H2YPRsqaLmDNdQrduJuBbr4xICpu940//+5486SPlVy
drNTSfxQ5mst/VRuqADzfx3lly0+Skls851oja0olEkLrH8+w42AqVFdr32/t8VcNwf64ryyu4JO
IV11lIMwf9dNvucEw0XKmLW15kPgryS7gPzl+PWTUXL+utI4RjaYrcMmmvBlNKVMms/bLGwzdTS9
0aEGo8Pr0B0lNmCnGzHX8q79MNo1u9mzCYp29XoHAFPG0ax0KV2NyzKo2L9rm/UAJiykeQ1Ev6+q
jKr8ASZOSB32pWQwxGeCWNFY9hu98X2SC2mNWrdF78S7+/v94ycT39WKA58AcD0uI7JyDJL8Pf8j
t4Ht07mP1mIYmbYxdQ1JyfWUwrTRaNDCtNyRaB18KyfAgwL3ZZHTtwEgI/W4+Q6tFpgdtVwXG0Kz
FLoWEIc0nQybHBHegIONS3JCl3eKimfj1ZfwhRwGTOhOb6KeMlMoE0DdowE94kMyAAhIssrk9Knm
ph3xPbU/BBxZNuH2rbrVLJbOJ1YhGyHY/Bv6CwaSwBnIx2GGvpHBQ4vfY1AyxbhX9RJ90KMqJjGX
Wk3MXzLVz+QuAhT2Wa0A6NzRdg51VUYzmwa+KRJVXDNP6KAnpjOJDZWUBxBRlkwA0HZue4L1fPrX
sDp+8UZSzBZScDn1Xi8LM8DF9tCg9SpkcH7kFePV4v/pWAlj73LuPsQ4lO4XaNZSK4Umzbpau3ZP
cUxjYDdE/gtRw33IkP9vjQm6OIx5da+G7wsTwJUtzBDFqbLgRBJYNSl7Eju8bZvt49RhRkQx/CFE
PzmmGTPB3kEp2DqT2heftxqcRveLLL+qhmQEDmKreSwU8p3FBBObO2eEEkr0zPILmjVaLIZ4CiAD
fP5Q+sbRYySrQm2Cr2TLLm3i7Sp0kRKooeUWylTixY1l57OozM64/w3QGg1lu5kvf1w/n2lsgMiZ
Df2kkWr+5ZWllwIYEayz7TKvdgTfW9TqWqMHbT3ctnf32qSg+3EnUGIZlbpq5m/fJc+51gGPOgeK
MQkjVssdnnc7OZxfpFwvaptLWplhkPKyQvKQZI5F/jGrWR9zcM3awOyUasnz4YZN4q+D3cC4ZQuQ
Wx6z76VW3vpAuAlNXXD+3fEDcDKXyTZ+KuWunBlciAarZjIG/HnLp0s6QeCK1Utsv8MlQ+KHqDJm
pv8u23EXLo7wCkdnJu9zC5M1YdX2sRzVXJQSea7izDgiazeCornyQxwYEcj2aJUq3KM4Mh1HvOGr
plDzpBpB/2IxyLMzCeW58DKAsFO1LsMsB+zOWLMKsWDkSzxEMHWB6Hs75Po4ImqEdFYSCC9XvNmg
BX6kyIOGw68qs0N0rIbTxbBrZVEp6TrcAOFl/N08pMFzAtsihwM8YA2RPChq5l/Gd2YIMnslnKwE
iBeM1snnlUAo5tkcVLsNdUB0+AfiIeKtUHPfnCQ4lfvEUNvwFBSiuD+fYNx7dpFshv+O3P+j45zv
lZOcQ5BDA6Zc3aloTtTnisXozGCXEZ8RgfYniePb/wFEFFJ04yg0EkF3pGK8uxCLtVw90rnxrVz+
5Ez/BvOofF5VQFl3BdN73MlAT2AYEQQke14xLOECeCptbppZ+RDVT3vUokIa2Htf+M+NOvyRyZok
MQ8iPnMXI/g/KLgDInzqfZUN7fK77GB2MfcWs8Knid8pFqPpjqVHXuWtKTX1OqvZRmxZwKVlrvzo
j12+kY+BW5CI3c49M64+ojE62RuScrd+ohZtsIT2ir/E5Y+NYLkTxDOjaGQxM5PA1gbyFeXMu/We
FhthqhgAaejtv3/sPgB/blP8ZsgmPsfoqk23PIODQL1r3oV24v1lIZfbl5B31iNRCEIu0z61EY9R
qeLlaRJkwSTwRM5ZhHsWyL079KahzmMFE1tHswCeWsrwK7J/wDKDmP3Lx1urwFVfJMLsKNyBcpCE
enpYE+Avws4mrDavvI3UgTm8dVeDG3jPBRQkDeooxR8uA5X3i3C/9w7s6hwGNmY6zpW48vDajeV1
3QvlQRHgPiNcxP2kZ2n5iYjjqagwsArPKfrd54p1ICSg8V5HKvw3M6DkcJnJSChAfesqnu5sPFjT
jp3rnNev8RpLOlvuy/xrLPg0ER3mGZQA/HoU0fHUoZK5+SwyJ5pA/KZDC4aTXNeE5cjEOVWfAqn1
hcYX8dsLRFH4PI1P+RrPNrPkiQtu/ry69Ri/TrjBZ5mSxrLXp/Qp5fUwotek7hAsTsY3/QrnEd+q
DrdUXo9kf6bTdsRfD16DS1QG62XxWtVONK2Q3DGY9LsZh3z2Bc8IfSYUQfgxmw7TYoSaRzUjQxsu
EEPIDMslqKPwfBimNTap2nBv3eHglbqr5KP115J5d1kjLjpaaIRwDEaEnNeP7e77wgw7dRcQwuAS
OyG4hYPoX0rSocXsrksXdyVQO0bQ4FUmFy45fnrtWWcSTSBol/v4X1N59b/TFHwPnzDCEMb82Uom
N0yNbvXnqI4REF8rp3JpO1TKjLgA1BeJB2f7XfmyIIMYH7vB6NTo6+WulU78s9IlJf+UI8LjT6Lz
9WQV4kqDRz4IZf0d+quDKc2hO5TVIeB3j0kydPCia67YbvdPr8B6KTpe2r0aQJEeo6J+6iPEeU8r
2X8tuO+ccwesqNducoe0YbcU4GxQPW9NxsIed9bn5W6GlUXOd3NdEI9SsTFsSu87/JphIvjoGemy
vnEpab+/2nIHxXQn5DBMlYHlWwRvp1dNtOWcnAsV4Q6ImiMcs49TsR9yOPm4Wg9hk5Pa1WECQYah
mtGNpDSjyTTEInQ0lWKgvwMisO5Sj0qVe4RZOotZkB80tySIviIlzB3SOk8xhr/d8JjCsDUQho9+
c8BqUfqG53w8rTD/4yOJrFlAeJOEAaGaHkpH8sFH5kOj779z8bp9MY1LMnWARpVOP7ggIYLFjGlY
jCZ4cNOMBaXCmWZFJ/P7j/B22t6ivpo2ShlrGXFarvESIg2ItjA4tlVShfcx2eE7RhQ9r5qE5xPY
vI8Y51huzW1UEVhn5/YMJ8h1XwpsY9FwTpXVKtmBEUpsWY1ZNwWu4tfqOj7snAk6CUd/+3EMBIBh
sleZ23Bxt0MxeZrBsEYk4xMYQyFyMVbmadT+cqLF9vVb2PYhKUHOqoZae4Xwyd7uNCJsm+gOQafL
99OXszslc8CMFC3s/5LO/ymX8X63z4Cp+jwghLYT92Hs0gBzWG2UWAlNACZ2zxFJhxnqLvgFhq35
6/0an7NmkNt/lgvqErDs4QrriIfKHABRldO2i3WYWFTpGjng6RpQ/hsNVBdXQbI8an2EcJmc0SAq
j1c3lV2UGaKjDAq0CxBvswJEaonk5qdfYEaZLUs4A5vmNgpbbGdQiXkGgt3xZQ9b17ytfjtp193C
HZgfgGRsKZhR0cLRFQvwl3sl/KPLYynVnKzfzc3Ig0f+/fUxzFTwNWPo7ybGNxqDixfoep/kVwwB
YGfqFy2OXcYw7ENE+7IDePfZTyK5mLmwiSC5oMcMjlU+4BFtC5lBnEqQIjunRrZSQunvPnqgQzmp
+8anD9kb15I33I+XfgFqazjNMcvXOgrhVbr7+n1h+Wav0xnYP1x5k6GkZ9ZXn831DxPidhh7IvZz
aVRBjIYV+I5TNi4kfx61s12IQpnW0NDA0ZnqF3qpTYvJ40wB2qL/TLMEsX/78FmhNTNMSIlpZ2Z0
8P95ESVnl8Bxlnj6v/AV6Bdw5x0V6fX6t2JurfgVXVqAJm5UY+Ns459lV4QJ5/pbY1MPR1YwAq5z
hJZMlFmBix5hLQmdWmsAE4IZZKILFqw9E53KeKBU5JM2JiI20NNLYFgUoVImFw5AvyTrg5dIaXo7
rm7K2HC0GbEcnHML0QhQ+Yyf159P8AuS1jLIOpsmQu8E57TLSrqPyiOt5xWQBbKYJ1yqejFf/wac
k8LiU10gNtQfGry4IQFt/DEPPGljG5AscamgCfV+T4EHiCa8j15l2bFmWVQAGJtYBoLbEIlhDPX+
+WoJ/nAui8VmJMJfw3Jb/3fN3w3EQjek8nETPoNHoM9nfKLQuVm5Apm/Hx1U9fDxjmFggyXzL32S
0PHaar1Mk1Eu0dQLAg9ynA+S4fxO551TGSO8jxuS1RNZ+9mPuetB8hOEpnn7mp69MzoEOlvu+97G
WLpsNNJ1X6UwKX0hlUuweh4AfpI+6AshecBMESUgIY+NVMKF+zwOrBGcJzBcM9SJ8LjsLzQ4l9d0
nC5UuB5oc5vpaQVM8zTWdgI7uk1gSHqANBDNJuYmaoPCXPK92z7groDdlZo//wjKutLoVgTjAPIB
2na0SDuuSKXWaAZEXdGmFnPdplgrQ+qfEqE3Tn6aYDApenRzt7B6kO4loAZpPsJ6pbYqaYLmQD+E
zgjvD/DJNPSGyBriQiiPn13qzC6q3HfoRki65+mNsyeDi9z1fD1c/KKsb2RU6OJO3QH72x9olntL
idLTxhK7NgjBS60pdLW9xjUFqRldg3ifvF5EaHV8ax55qtciA8JAo6jumMktrqBeZ+eeg8pwJEEl
kAp1PlUwsU21DJvQ4x1IfE1zpAXF2v70+7R0lFkV+J16n7+SVQLIs/0qhcyaH0eUtB3hcQ1FKBJN
WRn0bFkWfKLi+mBsT9GMQ9cBpBKccqsylmiRae2RMS5rfQ++9RdF92ZA5ODatbhKz3FqSfkJTSsc
xAotnKh009Hngn2Y62Elk4xEXXOvxVTQQelXzJeTsCslNzKB+tZmqtECc6EF5yh++AqQQHdA2icJ
RWZiOeayqwl905Aj0FSOhkclAf1pwRxCqPYk/cVkYLAYX7RQjz0guyN816kS2cVfQ7j6IJyQf8pa
uYqSEdFvqdt3I0zXSoV4tJDiXtVa3U/m8j/fMgC/novjZyrh1OuZz7OdliYnsMHIbpSsD6wwUVdf
gNW4mUzES8/sM62jyMdQUebK246EXkbwpZUCQpEKJ90PARzHmbiuLYTW6SkCHCwdkuiQA/Yd6/L+
XmC1jitb7BfYiSEASj8yN2hH9Tnxs3lz3EZbX7FeXO5SSkjc2dwTiOPo67mEQfeKhbhxBdSkkkbc
DyboiucU/LPMqCaY3KMUOeDNzr0ob0X9pQbYVMIkGn8Mb/SkcybkbfWRiaE8YVf5iDMWkFcmMsJY
9chNFbSaKATbPuWNfPQUMQ8LUIV/MX4WSYMqTY4mSwAuMQ74qsXLjhlDQLscpp/S68n2T4dKMy9U
gu7QqE9veOKAn+yHudGtR3WP1ywlEwpSgX9G4sSxKHmnLr/W88+QJhDBPgbg/LQxA5uwpsqahFXe
sOnY0p9B0pCcj2F6Nrd2eTbTNdVAaZ4bZ9vo6NdWVtkjXNiGJEeDekIPbZDHiKnn8unNx8Z3/RrB
4MnYyiELLAuFzyg5QAqXBeaISVdOfzXQDyyAxVbihUPqRCW2WGm8cCKgHDbabwcNZzNUq7rxLW+o
fdnmScxGmY+H53Dxx3eB1MLkxR7Jdf8J7w7lbHwTCESH2h8P0A6Uo/6hh82wlaOqoibvG3VjqdJ/
ZIqE1s3AffnkrIuTHLECFW7Q/DnYlwiRSHggZk18UG2KtaR1fZislUmLR+iXSHj47ewjbjIU3lxH
gbLHk9pJ6tPQ9clgzkldYy1V5Xy7lYzvebEHBuNCMBgOEKI1ctJVWQthMVJyghaKwuJORYZ99Mr4
FQ5E/yGVL6RKiTQoSEedoC9sREZ0nLbfHb3iya5N7fvwGHatztdYa8qs5dyVfsCLpoNjpy17nm8g
DLvMMmPrcvrSgz9vERVa0ZN9GrvsvXpVIKqxKyxA8kT3tdnvG65kdlr1/ePPonQdiYbWKFam3Alx
DDWe87+rOVWQUl66BWgbaOYVHb0KW9JBzijDPMz1Nx1g1wXM7UK20IKa5fmZpunu+wa/nb9gFu1Z
azh2IUviHtv9p1YnA8UgTOd5IaUPeY/YGimIX2q0+S9eYyYGC7zkwmfn6BYV3hQJx2gQ6zflkZ/O
Q9m5NiBxt9dN2sauSa5LgYQJfXZ0/eTsenNXHZ+pbrVxuvpcxBD3yH47oYte0NEVm5jcALXBAw/K
LH37KI2EljMKzTvmHAPhvdsarcZCLG34vbkjzGL6tN3KfcYA0e8QBhOyxzcgu5E2PCr/qpslOcyd
18LwcUQaUSmbpCX5VNEV326/rnnHh6cABHVT8SHHqG/MkGSsN6p4aizQ/HbDrYQ8KAS+Jug8tCql
PtaB9FhgrfF09FsbbbAW1Ifbi6vUTwCmP9YfsiXbakLx1AhYWPLDa+8M+/EUJhJ0InVdnMQ6JtX6
4WXWx6Hn5vzcaRJZkz76lnUXFTY82WOrtu33VGF9q6jY+BKXdkwgJ5jG1Isx+G6vp1YhwJ4oy0+b
0LiTUecPbqneSl2KEc8ZsXtvujDywj1B91682zTAt4Q5ql8m3bLtadzQ4WJtAdE4YjZ1z1z1mexq
9AOx6zb3Zlh5UczpTwJ3pz0zvAToWUyB6bc9PEBi2evIU3wpFqytxdcl3ZtgkEIw4DPT9vMcnt6+
dfx2uxnzyZKt52DhBnokLu7VIdtIGIDN9us05x3iIo9C9mDqPKOpxE/VrRFIFHZ6vt/lP1Tw6ZTY
i7viN/SLZj4v5aPVqVI+4mDbN20MUv9DJvaiydT0/VBvymAQe/b7Z/Gptk4RKKjPbqiQMvHLeS2v
Io5TnQeOnmbYqU8WX0v1VeAOgbnmCkJz5T/odAVrDEXI/CAVLut/1bcvwpUCJmihdtHk5M401+uJ
o+XDKwnzXPWW9wAJdC+2RO3Kib70did0V0psB0AVHH9L2Ghxn7tMMv1wNHmPG4SD2Z3BgxsRvcbK
w8tpQzfk7YmJr2yaqTkZLYoejlnOuPgR7UECUCQU+Ky5xHv4P5m1uTyvzXQhXbdrBBKy0EWBqBPX
t7NYmCNa//JJ6CzDqpJ1pwpstaQ29Ag/DS2vfB7Svf8ofIr4qajK6d3OgNRjMrEiWCCSocqZhbAv
Ovrda7qXnNLlRTXqc7Bo8Oqm3OiO2Si/eyaW4Q1x2wRPjagX2pFHktOq3VXQ5aGsqw64HG1XlrCR
qBKFSWn66JYAf9LZr3h4RjkJis1k1wkkViabqQbn1QfVcV4LpsNuUTvfy/DQ8z0ESjVrqNGqoAZP
c2HiGaLKMfk76xAPjKBcaEaB90pZwPeJwFoeZzZM4cZ39bQZcJZ5LQ6C78I5keZ9CXFYuXiCKO5L
uXOWARxa0+O+vb4ZymrvMYM2ZBwbqM3JNGXaUuwQYJgU7TThioHqEr6UOwol/QSo9pRdBV5ZxmQc
1I1TdQ1RB4iFAglPfUMybKhEjO+88+FP8pQcaxMUj+ioXEhfvoeVjWTNWPTlID7Hf06G0xc51PVt
ZfleTD6ChsplyTmqlcs/oJHnn4n4bJ8KUb6pOTu75zD6zi1RhRTkC/eVVAz/6f5PSyhBe58s4z04
9njNphS8B+XxGTOrvgoyI34JHJVHvfUs2x36mWhaIce65DpFQfYO+wi/CQ9Y6VU+y2/Fyn0fmucF
FrAi4GBNw3lgCyenUH9u9PV7UkRqDDFK9fq8VlRREcjxr580I0uBLzDX0nKWF0FqsZqolqlY2q2F
omWuLNf0LC76DGAiHkqc2PfYGVLR3lnsVAXDRv7kalrVz7cDei7mNSKqrCjvbFlhVGF6jIh2kXJR
aNIkUyKnSdieBCpilfZZb6JE4Q6iLMs5dLhbIJ73+Bof3Z3IK2bzxokgU7m4UBq7nW6+w205m9vr
xTJ5M9Rn2tccU+I9uPe/fhlwmJQaflfDxntAIhGmlK3A+UXREph3F12bqm0GRO3INSngq/U3Jopg
Qtzd+sk5HYU/+WtDO/N3HeMIM7CZGx2F3yCrrn7aQHn47hN+/ozYTnQoU2XHztUkVhXrh5eo2H84
QtEuIkrbqq3uFXlViexyVyCj2uvoEiNynyOx17niH0jcH8Cq04Z+bC0atuNkchzvsAqBSvbGmVDP
xFiOZFg8iui3X2hV3+9jPfBGARKuSfarxDOyFOVBFJo8a2KIAfXOnXbQ7AlHNFpQjjc0EUUy5Bes
Wgu0BcsIlN0Wx1nYs9V5HSql0IowgtFMfCyTPHJyB9qLRoox3Z1qRsglOsefe0mNcSgGZaItmpMK
Fljhd/MfaYDIazYa9Iie+MpyIUXKsPQTLhdUXNe80+2sut0VbqDACO4byCh9SBmCtdWtJEXqA/8g
iIjY8OUNEwdytGODhWa40aiRP7nUYqdTqpkfFwpKB89XWh0KgPwbzpuYqUC6D6We5KI9rX84QG23
Vm9DDhNf9C/OEGxo0I2SQy0Tz/cfZRRCNavpzLK0GOnsuZwQXtwshQqe96FFdaJoEgb9mhMZE+GA
sotsMotavYymX8qUZQWNey88mdmVF/vZ3hqbALeTFSOeT1uKAk/al/BVhAqVs1TLQpMOOsC7b6v1
hbzSqY5eQAJulnFxyHpbOl5v03QM7NlPsVu5lkXTmKeo+to0aAh8R+XuMPQ5ZcCPQhRbWwHlU7nB
Uh4Zmufzi/dALi5WgMi4+A42MQpJgLI8Rs14GjRHQd7AAXJbscgdBrtH3eWVlqcjCFr123C3+mLu
p+SD4zKjn1yt7N97AflHbnCXi0cSilT08IfYrxfG6nvQAjAg0jGOhTyXDmBeMyzWH1VZw+jZyzxL
tXpZ6MnoNUarlut6AnS2Fl5dWZiTodLhaFMqwD1spRuEYXoRmWGk7F3KWBjkON+BZJhs9U+h73Mu
MwuDCKafowzmPysBmoLwq2mvZhpQU7pi6cc849RTFpmYVSc6Cj607nmhlpHosFxrNVvjGtr/nnXX
79GShd3raz9lvA3q27amH6c15inaAakNKPVAYMe0hexCcAV//dFmgmb8AWLhX89mlbwXsSWOJ1V3
8NGqRYWwck+9fTQHxG6lE/bJ2FIMUThhRoRuDB9ZuUehhaK74lxWL79GgJhaOuvZFpdIopSpXiL/
/4zrrXNb04kPU5aietPpnGtmcdJ4YtNF7ks65Is0Eanny57OP1J8UrEE/FYfdSbz+MX5omTmz3l0
cTJJuXIuZyl/7SjKfN1TdfeLl95wdUz+tS+SR4UHLPw9nLpBPOKHiGvnbvTLp5vVxVboU0AagmTy
Wzc9XHIc8TpD5SmEC6LKm1g7q3HZo1Zlu40gX0SygfEWVjlfZ5BHKGGqdy/5xkWsAmxbuXMC2/4F
bH2rRJc+r0W6CW3eJlQS+7TZ47OEHY1Rc4mtC2TUtVWMNAgUqK1yB+/pCXG8sTYq0RtlLIK3F5bC
fVRohZOwvP4TN+glZGJ/4qc8a7V9RvfAQ8GjPOUpr4WTWLOh6CQeq70lSWXtdULAVWnz0HdI23oH
y/4ve287FBV3kidzYd4foyX0tBxRanjei2tkQw5U/pddpEoTngsS6sOqsJ79EWP/4fl5Q7wfnctf
n9WsPjKtwwZNxKIK/Xx9n8YqMwRTv2FPGhNRGtw33q0MPvMqEJkPMFza5dAhPXWLTu1bcx0cLekj
zrRDpIyUJjCQ9Rj2wp7HQc0aS8jq8tL0uzMNOBEQeAi3ruJYIMCOYQ2/OGtjwNQlhUEWSsVSeMZ0
0dRUCkW2A+QknhZykpAO95k841gYnkRts0NYJuoAxUkLpvN5m0j7NTlsab+mFaiYSZZcjuQbtT2B
daVrMmqLK70Fc2yWFCZbCVNTHb+CVY4XQTs62//4yRZL4+Qn2EiN2vOi2gIM3m5RYXodWz8LyxAu
EqIfutu3UsQvcie1ymbwaqMuKs/mXQ/xvTq+92oB1eKXQyBye9BruNqCjrAr8/ytogJh99T90GM+
zJCHMvN/AZ7kLFCpuxO+eL/bLIutRRBuDqAf7jty5CqBycR+4WxrsER09D4fUSO7DxdbuSNjR2oO
kg9xWiGwVi8Z8uVyBGUBfW6DCzyKeslm7hK1/qQeNvmCpp9cYWv1vBjExM7MjfuRQ+k7UYbunsr6
/bTNQ4Ro9sbN66kFpJvjcd30iaIffu3HfePZ6V9aZvrR2l6ZUQjJ635nTcbYEgcLOkXgmQeA6QAg
UwS25kjUHgoXHdlav5HCHSie+QH2bo3E7Px1Gt8iWpNPYdve8zK3NvnC5pW5B+ooXGVRl4Q0vKFy
TjjiYXcFxRoVlB/UHlpIfq7n0AFuCB/jxIQzQ8CVuzLqS7SKwgLBffBmIcvlTbWXpI8tClNBJZpu
gvzpyx4QEkWRDBWTBM/Wqe4k/nrmYtUoFQmlmn3huSjUDbjIlgIb7WM/DgF0jklVbHgEapArSiad
0cIL2tbzU8Efnpeem00ZZPj4W/j8Y1zS5n2gUxKqsWPoUVzMPMFrl5RI8nmdpsOaGYIjtbHL2pRx
XuwVjVcQRaIDqTahYbkHEi9dEIO2dCpTDJQGQhS7MEYdnhruLzscMzuZ3++wFRez4bOpGnpdBS8G
I5gouCg42QzlDwjM06YgLJQuSp2q18bDPklH4+TSvMTQXlvUt8IwMjcZ47ldRS1dpQkYwTbsjnye
7OSURRRw4zbBWPfikzv/XSffh51j/jFaUSaQPjUuQ9e5df/WJ31oXXhDViy26g6Bm+hs9EiFO+qf
KTESCEDmCAoO4I2/4xTPdipsWY/x/yf1YeQ8tcRIgiiAbopshYVlJWZubhtryzMp4+27Z7r8dgLJ
pLAQcS8B3J77kA6BODieCzrgjOQf5JbXjhSdKWWyoeEIp4yUBsSJFrOxv0v+OmNz426xjHrUpB9l
s3ni1TE6HfC6sx5ehkPhUocsvUobMKQAORPivSY+oivKhEK76wRFJ526+zhr+BYHzW5Id4dqLZyT
Kd8ibRWxlS5fpFA4WUqX5mWdjHGV0sV578mL1e7Fu52/fzgIEohXe5GuYh0jmRfu2M/1oNACRF2O
FCbLbPLt5yH0uPnX/eOJYSzUWJ2QQl8SEOoiawQHyws33xlbvbKQTiGW9ILT8MxImAQyCZ9bbEEs
uZm1jgzs4NkOXfCRuc1BlFl/ZqtJ7fO7sdXJfSysz0EninOVNeHxGvuXuDLjprkFgI/sIwR1f28n
fF4f60Wu+4pJKrxnf40kRgOzIsji0x0aaVZW5cvQnRczkbZ2/jLqiGifQHOydIVl8cu2trsaRfDS
V137g/CyOC0fEYf/xW5lya16kdfomIidFbZmOD/vkixgNJV/Rah5rconO86YDm7oDBbGvev7HmJR
jaPUT+dHYN8rRh2e3qvbEwEMe95m/noA3BsmKMiG2JmhhybzUv5dqZdpmtBHyrXz6xvIxBPMT6bL
p2HEMnbTYxhQ3nPnPY+EFC/5j850a0kE/qUHRPZSQEMDtBTX5I9iTuylC0Kh6KQXCmSd5zIHINMW
SIGhS08QScC4EtextRPv/WWw5g1YCnsddPKQqyNENcPxe0LcePvI2Ex0yMsWsv1kwACJN0TE9OuU
pDmex3HniNV9PGRNP4E60cYJ/aR5Km/pJzg13G1amH2uvS82XU7VuAgglDgtIZvOs4/1zyHvDCnY
VkO3k6lOXgTIwfJcXYqcMZ06U98HjDidDTsAcZCntUYUkBmRCAz4/s/tk43snoSH/EYjLvcHV5kY
4BmLitmV4Nd6ehuqUhyshjzXrWRJVuZeykIeohOurHmV3MXjy/gMNpntqZYI+8A8gG6rbGL4uvuK
TzcoaH/XZY8BYe0XLRVWWApVsoT9b0JpRC4NW0TlBfLAFR3Yhb004VLuDZ41s9KpZU41Iu94UIMQ
H1hENWGDoRHUx+vBhjyepwzxvPq8KKotmp9vmhnk6wD1oeehtoXYtUHbJ6DzgEcPaR+YCiqE6u+/
6iZ/XRkUH70XJ2yY0FGEOg5mfD2cSM1CRHgFcWnjXeRcetnSZaZxMwWQGO2kdv2i6aVpjQDqmOKD
RcDypt0eVjq3L1wVrLZ3sxgMscDNaNnn/IznuJYliON9QAKttQq8XNDrEmj7YwVrodLSCwRHd3NA
vCFQDUNiLgcoUyAG7yjg9/uCNdKRu6rfsvl8UXJeRdnmW6oLiK9/UemtHDsh6Ut159vCaZaYePl2
U87R8XX9MPOp3JI97fLEPOFHxnpASryWz+B7Rc6GdNGjSQl/lN2elFXBwy88yKF0/KO6IwpW5aX6
CQQVAWKC/b6sSNMiYH0HeY+6Yca/NE85hXTW856rBf6QTaN0mzjpmj64LD/GFDVYZN8dsBYGWERN
WHGRYn8UJJjAQ2yMrPOe2WYh9u04w1dgbSE4bfsvKTrSgj63+d16wYP98o4OD3qoi6XA90u9buMj
ftgxSL4MDbzmSHsa2V9NsjCdWIhif0IwzZ/ZPCo12HDMIeLUDaNxjUrjYU71dzq4n1bVH7q9m+7S
dc5eZrhAD2KdA4suUrpBmlOSqNX+b31kfewksl2Zp0RNo59hg0G4Sn1IkXUPS3whZk8sN6zDBa/H
1kVEZbFE5RhGCdEudzcZfjphimZqc4h/sgKbvx2BXA3VsWyaElQx1HpKTN0Mlnxmp9gde5VnQV0U
O9eEv4Cj/Ofo5ieGvRapoMneYX5ltcY05ER8KGB/95/etEdtKR/Ne/EiuyXijrEBRd1GuWxmkMpz
Io39eF2Fx8/bUX6+VYijgO4j8z2lvSwd4xosDs2olS9Sy8gzUWEibGoHgXLPOUA5ZS6YGcvcO2LX
q+2WADZn6gQ0DcMLLphCa8NO+0zmxHZSEiV9Wx1wEPxO+G4uDsjM36mHIVhFwf3gO6V/mzQEPpAh
ndWFoG8aS4UKbya+3gk07JeHlmFsEeUs95rbrQfWuge0fdlKJM72eLk1LJLgPQB9VHwqhTTH8u6i
Iv+zOGizKqNj4IU8MVIYuM037FrKr9+SVGgen6lc4ZdZgvgtRO7lFm0gPXnc7eTq6kdwXaq7NBOG
FKqySzZVbJdajkSCCWSABylml3i9AcIACVLhKWTk0Deth0u1A+MwiC/VbwCs7XuAPtojpauMMcPs
x5y5gAgrum1EB6OTSj+PKdSfh/oE2BZwzxSwJlU0HzlObzjTjJonMfBX6u9IvUgyCpV6+wZbCyfL
Ww+W4UEErunBPvf91dZE+gwfghFQUuV7b6aspN4YSk8AOqAW+nmZWG0iLVvoyvZ1m7h1juYIF8Mk
ZYY95AZEv8OWfsCa9sEgmBdLK1ACCSmvUfwH5RzxRZius9FvFJWx049P0WoNxZ4/TvSbLQQv7ypc
F4Pu0duvZqajbg1vSqmnpdjf5XPI/1vOdtOoTGS5zNk6jA+pK3RkU4QzitOgPfTlsShM1yRDMtAn
1If3Q/yV4VgDBy9zvhX7xT6VVPiXMIUVH1yUNdAZF0h5dI26zBQLO+eAv0V7cCZUbfmsbomjZ4gF
toRbhx4XbN4MaRTejgs3uzLKjYxRBClKBYL4/qzMrvG4L6o2KWezQTOXZZV4NaRaRqgilrQoAE8Y
jMMkz3gqgmHQvUKA71YsVbfDQWnhqVxTEBKktwPEIOkbNYMxeG/cfRCNohfJ3JA4mV4ravxYkvm0
o5XN+PR0joVxKmBb2vUrWpZpqvv2YOTC0ieN57qOtP6wv7X3xDxqS5FzHJe+rg7/fCMZ/ZMDiZ5t
mCuK9o/0Pvew14blbnI8JkSgbRLLrep5c13bG58aS5F+skP0g3SZsK9Ju/h7AtFtUVN6pZVdWFW/
FQ9suRvA4dM3lWf4CPgtslASNwJPizsCCUg6QjB+5cUytcBxAeS1QtDCDklL9nrqzxHAs1Xw8+e2
DQFEsKfdwdn9LgNrFUyRsP/fZ8jlGuFTrGmTdC0MN8T29OY0IvAiH3jb/ImuzXEB4IXmxiuaHvO4
LXY7Ssfus/3AAVuwDXH07I9c1IG//zvS+I2CxwjVRm1kiUtGZYjEMJTlcr+pSup+tlaUQax/s6WU
EDmfgzfhBNCJkgwzsdISEY/3ffg8feRTkvSJfYhDULb9HqCFDSXdXe6HQRjLKlyduYoNW95a2/cH
FWx46lsYwn8kJdcPd0+N+QXbEuYHcbCWe/DQSeUFx5YNQCM1vVP5Ty8sEaqZ0aj1jjqx8B5DmHxF
Ntkl9JvfskTSL5rHRKwBvOEbCvbEX5bgexzUZg2Mzy2/IqFWvbbltOHx8yMTC6yojxKDV1clTyeF
In9MQK2hTuow9CFC2V+63lzsLqjzO0EclazyIJx+MuIkHOQ0qs4W4NadcA29zB2BG9/B0ULhSp0o
Y/up9+He5j3Q4tYtGHvbUvG/qbE6GR8YG434KRfVtzLr4ACgp/aD4SzDwMrAFl6qHeEA30RBoLfo
IRIKmivYhM8ZsFa4ZEzcdH2lcixOX14WmfX7sT6JqktbX2csLnw7anRgvO82TMFFsuLVubWosDpL
Np85k2xA6/6Zw9N6qv7M9CgD+ZA1tFlLDWPDI1OwaIkuLg7wXYUDqTxLIMKDun6y2sprlyXyXvUQ
HLqTddrBySfl6hhpb8itlLkEPoExMraCYUdgFFOv1lghE4LqdE251sBhLExv/AjRba7J77PCKM9f
V57XwzrIBfMukd0kWTfoxtOLtuT3AFQyHKEEF+YsUUV/KpkSoiJbCl7yJwZJCGq50TNZi9YlT+Pb
rRPiU0JzosXZ1nP/6dAOvBTTG96xBaHhlvu1J+JlEdFhS9owghBPWqOSV83Z1QL0SOga8llAVW71
FAoB9oMCrdNbujuMp1aX+HaqMKQysWVqjXYUKhW4IczPvCQ2kDOOjn45RjVjQgvtI3LlbZC+yXqR
j5Y7U9ozAeZvkPZYLlKFJ6sYvrKmG8Z6mh8DSMQLM4AETdZwJvWQmyAI56tUWI31r/pTm/iLwNcd
0ACVj5LOtv7rV1tRRTP8U3FHIDd9r2HGSvyn7i4+mGR0o5u38dGpDezAX53G0wW5vjmTc74pqy6G
/eE08/0mGMviH7J3VXsv3+EWf22vDj4dD/oZTIvRwJZtBPfeMW8zeYZMv9n1PNU/SI2JWCy04ZS1
SO0HjKaZ/F4r9B2jxZJjkxvbKtiDH0oZmoeK6flvLjp/rDBmXl1DFmVG+8gXVtZj4AtmrEN7OTTc
ST9la2gpyAgbzt/XKhaPRBw3PTNtSw2kOtzbXriRtnBhfxVpqaPGzF783Jk5prfgK9JBwk0UB7hJ
nWVvNg/btccpfXCQUmV47xm29vXbgRTPj61h4I7KqduJUlYxXsHKih26LYKZMKJBFcXDx3+vKQaF
FpoiSGOWq7cyt17oOgQ7Ch+V32GXVkV2BZpPrD0WUuWT+cU/XWvHHxPiS98BtRFhGQ4xtIGYH0yY
5/WVae+ukaj7I5DTlEDaJoAz441jNts7bCchp0I6w9g3So3c0iq1dl8IWxMw6d9DHUEnv0gJP083
PyrPF2NCMv5yY8HJa3ijuKqyQjPmay8Db7GqWoWWth96uQ7UNqXjecj/fuGPlCFcslVahV2tNmvg
qvTll/9PEK4SKtlRAQ5Eiy2t+IFeJ9xJZ7Pw1tnCWNsm1JJ2NQBYDiVMwUlynB5HzvD3N7jsvj85
hE6KosYmITx9r7Jhdi7eQodMAeU8X9xbe+7JEQqC4TVw9YLVBAn3gLP7+y9m9B/z+QQjnNnbsAIw
iP0v2hVMg0/bMPw2ivULItWTd+K59SFGU1nPoAmwVr/kkzNFW4aBnXEDYWQQPhsOfhX2rkOQ8rMa
6T5S81eRG+nC+0g/kWyQnlDgr+S1VHiN+7JdepJLDp9OBFj0TAdZ29ZQPLVHyZ8lYk+e2C15irS3
EkQsqrCUkBDksp9D7M7qu6w5gc0qNTI8nBNi92v5eubJL+AvFy4elolnsGkasKlaD4bs1Q5Th65W
i9ZOA+Ja+S2MxXaU70YD6G78GO4+KC8jpHoFIouUMnEKzWK8zIIIxKfSb9qUcxFInyl3D7cleIb3
ckCNhR/veJ7gOXOEFk5L5tR92+0j3zv77mTyFwqQkp9+axMO/OGHLAC5KNh1R4AkuTbREWqUoJNp
ee5EQKuDJOglFbWALGa1ZHBjubtBf8D6scuCTxu1Lr7KWlUyv6KgC1grSoyM4HWEu8ZV1xzd/BPW
yymhHNtV7w/Rq6fyem7ygDeNWlJX3vDZTqkvWOQTa97vwmnUpIzP5+vKSswVEO1MJQTp0KNHoL3B
la4ffyuAmgqykWlhpVaXw5c869fAa3YBXIx8LPg0sstvT3JTWOs/aSIWzUxYT/WjKF6jMHHUnpw+
BpmnKOheUPCNp95vBnuwKyBuYzOzT4RUjuzyqOHigb++S8LoyqU8ml6lUXTh64SiudpXqtIeBZcX
ydEfTCL2iKPFlq+lEq9kq6dfifGh5WlGNyRrSRTd1xWjOxPX2VYT0uBmgyfcvCCrsCzQEXDeUJo0
W9CpHUw6AxxR89Qg0P8+yfiwrS2Xxu27FgFPQPQXOHC7RVI+gNu0IRJFP1POxBBip/T1GguEdK2E
0PFBfk00fi1j0uRL8gxS1l8cPEBO1wxdG80BaAMEa67A5BLHSdiG/OnCpiJkh2NE1EyeBaMJ+Gtj
7veDL9EssysbepS6Rz7VEwe0jH0TZPKwIpQgPJy4qZyZw5LVPDrujTNN4mpDpbOMN9IBgzO79/di
vr4Io7vRjP73BoPdJZu9tBspx8V/JY9JAGkLCZE8huLbD+kuZlN/Cv+xcyaCcz3cLfB0FGEY1Xyg
ZSIqTtDn2xDTRsMyp7u/sY7S3JfRaNjY8vS/ddg8K0ut0boXhW6iIlrLeSIeE87irx7i5rQ2A3uS
tofTXTkyw+YcP93V/VwHvYRXVDIT14BmdV5eTvW97+R8/X8zDtZNt0Hhd1LzLgYZcKHM3uaWel5R
IxQ5S2gSnSLKY85qjSbXRZcSHrOMJDcgVILm6fQdtic43xH+K2DKMcGJF34XFtEdqH13W/+PijI8
uKK7pb8jbtXzgtIShdtADJw9gpoSFrNAHO0h6A73MJu/kPbMaPBQCLp8qg3xxifhSGAdaL7jfuLg
S1rTXmQ/ksspQLyv2UpNoawPWGy9i/rdraV4YuhWYhqsbMbS9oAUq8Q+oUNyBFY3G0biGCYxZx8T
Cb0Pum+2wUdOMVo1EbSY3ZWELH/6tZjNG1YiCf7eyt8YBg7OjhcyXeZIqrpa4ZHi2bOW/c5sQukA
Dpcs6iER8UYLmg1UcgBJjFO3nmLYjSmc+oypVKc10CD1m6LOSJxXXvTuG+amMbVmfIO4YF5SX/6g
epkRsOHcVmFGH3Sn/dHUxQ/yUuS9C+qgOClSO35AyhHp2Morl1U1IDltlMaefjMDZ60YUEqqc9f2
vLLtHrOhTdS/PlQIzfOB0nPeXWhjbWB5V+P4Uiiy0VZqXqneUjZI0FyMuekwb3uTM1It+1OqPohP
zxAd9SBJ11xwo/2cOF/fxggNiw/iQqL07xakVj3RIri9gKUlCgjD/P/Cu4XTopp3gFJ8h/Gjc7Sr
CDA84BrA6t3HJUaRmFJc4OVjvP/KRg0aXNPBSmogXVtcH8I/Y4wolqscDkR0zAaDXPsLl6CxIugR
EK8oH+KtG8zZ51RPg/uzL68t2x1xwjbZMKwuh4Rl9OkxCnGvYjYHUGtA9zv/EOhP61oPMCG5Hyl1
JdwJd15PFRsoPuqcfMSDmJYZG+E/PCPaVLqDkyqDGgeR8d1tOxMpzzthZosa8eo/VmOmRTBQP9QM
D/5aWjUj2RayFmUX49lLicrNmNYa87hR2qT9Hht5ll+12n5neauLjC7fnWPfUBrvRb51VyGuniFI
RpaSBvv7hzWf7rxe05kOHAivn7/PSv91BdQOAOizbZ5ZbsvIHRbeIUj0gZuwgaUQHMMQfXnQolyB
dt6ztmeFdHraFR0TjgPm7Q9VICWnOfe2VrhkcURm4ZkTq4EflGfBUf+KgDY8gMS27WZUstgoVK2i
EmtJsf2g1OIVZHh58onWx1x0FW/hIFB4mn4gqHZMsEExGWqhiQxxqFBQK5TBhEAlfIPhvePpbDu+
dzNMaMOAT7CNBIjDr2i2Avf4Qyav6PqX6LQ96twx9CmXcMM3Je4O9snSh4q/9Zf2uXrwdz8rkekq
d25QFzDxGXUk29ptMbZxFDlJ0dvjnbkySPmcmtCtzIRheMZqG9PrcvMOOPqc+e7y8Mf3aHaicOzB
WsUkNLfhF24fHI+/nm49J9CsrKvr1+ZXijSBuznSVkkvA84oXPSTdURipJFIp/vEvaqrUnO7S3OP
XdUXRHjxsHPN3h/yN/o+JRL69yBAO2/sXoUTqycMVaO0mYtwjQXQqkucnc4vd+tYQEIFYmMNIsMc
FJsU196U0lc/Me04n/P3b3BX38GMCHr+x/6GMT7VkKxTpEvLWi5yt2z/qL7MnGom5qEjbgtSKD2q
b4tAS/57Lj+VC2fn6GTZ68Q6tnGCIFM+JuCdxDLXEDecsapfsnO585Wd7v6LeCvLiS24Up3ycqNn
RpOOv15HkTA0mf2fsddFZlj8Dq5073KM64aD8nI6YOrJioy1xmRgiCdz5VFFvxADspPXpd0lQymJ
dTVlQrELEb0kFpZopb9p6XNWWk5mpR2rOC1vNQn8PNj9JS6xYyUiHEERPvHV/O0TTmWWDDzxn5bA
VqZqmX7jGHrvlChRHG9FpjjbpUlnATfjQuAheNkGG3EOP0yuqOlblvXPyuxOI6jHkLdOMwwSrufo
k79BF/yZRvVG7DCRAfCXpjQjlRiB7xqC6T+FGYY2JaTZXE+OobRua4Zn3gyqICbX+JFQbhekP7ky
36GEKMzFthsdJGC9vbx6MBIuJg4IWuOLwGQtFTPzNcpV83ZMkpsGhJQ05ZynI7iZyb94Lz2HYykF
tZbEqJmJESevrjS1NM0K2dlIMdqf1Jcnj7inPYl8l1wt0frwimpKMbYxj2Bq/dQD2s3DPN4Npu6Y
RxacM2qtjGfLe0oXCPAGAeF+U3tNwIPU5WYnvMCt52e0Optj5uCp7YnhNM43/LGb5iMTlQ35RL0n
zmhcIM6udU9FnVAcKoKSg8vQ7nTTjlD+NEY1K759VsInyyX6KS4uolhoGiGTGnLxfNbidDpw31Z1
2byYkvyZk7fuSj9UJqKQYMWcPyj11iXC0s2oTlKRwg1GeGgrL30tQJrZO1JO8ewp3e7nQT8xmcrY
Y8SV1UwgH9HKvcNgcdONS45x6r4+juKzV6Qjpd+3wTm0BRQtO17N9aoJfyCvJI9jhg4AZLGUcCWU
2rPvPF6z5W33UsGyEtas/vVqKvpm+V5A//V8iH6H0hU+jJ8E0Ma3/PKXZ6tbjQgE1UtwsOhsNRkc
41ISm6ESDkHa/Yh7T6eW1tZOeIGVEVnLnPIZUDnzHN7X4Q6iVKA0cVBqUVx/FsVTZdfEHf3SsPgM
awIO7cywSA/amlq5mb5hcImzroy2nVii2iSxr5md+v6RhPyQQ/iO6Wx1EYLfPqDRtt9y1DNb+k3e
QT7ubeUaJtotvGpmzjNf3CIXLKIVRfXovOftaXzivoq2oZ/sRRn1lcZdBWgRf5W4Tvb6CtBPdv2i
EV3A+bXerhZfejHrynkdEDtxzMl2Rj+1xq4yp0VxftY4FZ5IjwNy/g/cIBWuIWleV1vHiUHD+/PY
MzKzl9Nl835Tcl8wlaicwv246Vpy1202qdo0R6h0y4ejqwYdPi6yKe8O4Tk5oBOzjLT71TrEPSQi
9UWW3aIq7l1bh9A5EPJEvBJQNZrZQ+PZKHlVmu+S9gckHjrQSn8wH1ezwTuXFqCv+PCCjJz5hX+e
czJRBsKuGJPK4HaWEHsNXrftzhLPvVivR+kA8Wrx7PGaxqDybWbvLb/bSj/hcbnOzV9a7lng5zPf
P/bJIs17meDcBIZj7O5xe8RlAI9V+ylP0Z3mnLWL+i6rbqP9qT68AdUrSXmi3BAHm8ai9SqAeblM
jvxB1RyEINfcEVNIr7DLNCX1XoT2OuZ7G0XemzN/AkQRsx2e7NbDJBH+2vX3i//LO9+krqGwfWP5
+wefMBFYF0fj1WWwBZFz1gmEXTnGpn1YLeYdmUDmXFkGT6zSyn3J8YnEQAp5XJowyrioY/rVCnij
Cl2OLtjwg4T97pZ+RUBbvB6xhRzOF2YPGui49F/C7wND7f35MX2wHdHxr+M1Wtud+FoGwtQBR5Io
JixxaDS/3SbGCZPaZMQlPgE0VCpGcda7fNgF0lMOPe5w1kD6o32iJ2o/zVEoPN+FbyCoA7ylN+pB
M9ciD5mZ6q566dOKIk6snYQUgYipEK1OO+ShLzdKmdAwMuwg1GsfIgs2VGdWCe2FeEfv7xYnq/sr
GycUwYwCQv91DyhIGOnRnrPgvh5bzHJ2LnIn99k4QEgzyvY42TzkHrGzpjNi8iuVRIImwTSckgSp
EqvQki0LhKWdngqC6xKa8och3+HsPgqgd+9L8TfyCCdEJncovBkh2hf15rDOdOlb2DLI8H4pAG33
LqhQbPe0sigAEQ32gmiBgp/bMRc9HHsBZCiHG6GNItaNzW7sebq9fSeza77JDspZaWOQUIK8Z+YD
uk31jImsgKw1qJDo5y5k0x7C77Pjea2s9b7QfJevRWdGvU7F+HoD86hxLDfTDMncekqMMAe5jBGe
tENK2whuSR0pWLYFCxphDa33b1Pvrj2j56KVjmTH1Y5dweMo65ICvPZdGQ9/eye30zvx7lGqhE2z
dMr5KdBgQJorPNW0zmskrGsaAynQw7GPLiYsMwqGah86oHYYC9GIdJo19IpoecAIvyLlBPfLb0/C
QcaoW9qj4iamIGZd795qWDg2Lo/xn7xfSDdKjApIXzlHFC+dWdyKL4pidhTjVNlEymconPXJnBE6
fbLTi5jiSiImgRGjt/hcxBm0IbDQlkHbfDK4IqPp+0ezDkWe/yRQAannSn7mOAxAVA0GLI/dXU8k
HWPnCugFrGT1SUehZOiBeeR/HU2yQ5EqZyba5QGmOe1vfrBNl9G1P4ajhhbgjOF5mkasskioHfBu
+31ZgsIPlJy8XIlHoB/f+b68mO63u9Njs7mTkrQioRrYk6Cm2uNnpr/dTUPMZFb4RbuAbiuqu/O1
2w8fVTmKu/6nuV5hvxAa7tVujJujiUt6HdvLYLtGh/JC/1Jqr4GsVObRIN+zLzCzQl3R4NJx5gfS
xRmpDouKDnLybt4fJgn7yV+YYOZHQs/JVWofmbnbIGGTt7T4o01wSJqkNe7UtjV9k9citOL/KUmc
ssAvad/AL/+HWBHFfUmy++DWjyTCJCmMBYr/w60NM+tIz8OSK76pYOPgaYDA9Zuqe3Yi7jXfPqEL
i4WxcBlhMxxCu+3yHqyIgwH0H1U6EV9fg/ZatFmSKXSNxoypZCMYOMdWa1qBp6UEa2fDM6h/g4MX
+E1fipTDJXgvgdUZNSQKNsfqepY7OcGtcs2AJ46BZv54kFuYEF+Z/v5/NnLBOBovgAXalL6trhf8
3OU5PtaNe1aqz8+j61PpDyQx/IUXAkYRaxgRhb2WK0uNbikpyL2EAde7yUkuG+zmlzhpQRgq4zPm
IcYg9UWcu88J09AANjBdbGAoOYvHDk5I855AnvVmli5I8ca9UGq4+6jhCEK0Uew+BmH97L0xPVcT
os9K63ub39jc+y6x+JfcL0gt/M98RBsQuDDP8ZCRsb+QL0kPg8NlVuSvIOIZIEIokzwvj/J1YYYY
32ix3idQMMtMkF6XRji99qjVU3pJfsFf9Amvywa1PlOsjZXU2hevdPO+FqE/1BvnXPDWglC4+INd
zHX6WiluCeCg2zgLnoMvIb3uGvyWxL+vKkyZJ8o5ANNcH0vU7UKZUO7oh8seV42joMzTp3h8014x
2E5hYGkqxidg11vDjnlg34i6XvKdHffYysgfd2JARL6Pvt6aS+7gTRXS6QgTcuFaetaBjFlFR2sF
8usyZ1QhJtWeu3R1z+1ZKVj9cURTccPR8NOo9TfK5jvKqYCSCSjstE7RY6zr3c2Of2Uemf5t41V+
Kl4HZU0KtKJiCD1DYoY4jUGU8nngfsvZb+7hTyrl0vKbhHFZSRbc0UyAQEjitYXYwLS3DVPa63N5
YRmbm7xPFY/hsD/ugkDBvjDftE7T9W1pLiHdFmfqLPDcB579wETXQ+nRRolPj9NmRqZr37LXZTAl
XvaWBkgb2/Rw6iUVj6qnMCVpMa+7B3MrtpA8hbnbYbUz77RKM1VEZCR9Bn822Ptm8ZgAVVb8hEsl
32NS075zfv0qqu0NPuy14lrPNSQyYJTH9dqAv7V9KqfaaT2JJ/4ERP/CSGPwbLflhiB4QveScbJK
Tl/ubioi/jMweoPERq6Uoq1xjN2UjxPSYI1Q4E72X6B7LJJEciBpiX135AU5bWTRbSz4mNLSFu0J
OUJJa9zgkS9DzWuBnclZyD3KvMzoid1i0uY9aj6HLOnqjDSi/IB3LPiGgCbQhPH8uTkHQFhbJ2Ci
YQ8WQ1w6QftQHsatCs96ZRfyOvoIvM09dWsp4UZThOKGU1K9pSehZq/k9oRzRa0aQBdIZC9x8sJa
QyM1ivVye3DW/htvJcouTFbx6yRNHCjnxaZdvdiU67xXd/AEwu7TElOy7UEKSJMkzNzDPx2loOZw
FWQ5cy6HuqtUgfFK3W+035AwAY9uhXtnZ5FaTmGS7ASAzjltYqTu32Y7k3ihjeoIsZCf1O+FyYlb
YjItVrfgLLb6AyT6FKHwKDyfh9uwkbRexKrGUVxvHivCZJ/koXHoDufl/BzXBaOGGaMUy5Q8/BFQ
B1jFXiu4x0yP0XSlloF10tEAtBZFhg8Mu5Nm9aOFZGvJ94Pov3DDowHhunOow7qAkynvZfXokaCq
UzuBwEKXpCpEY2bAD/yD/t+wS/gDwpYL1GyuZJs7Xfx++exGbdK52jy4obEYMEWK5ug648Vc+gLK
hZCz5q/vz0Razb5zB0ul6RJLohEhlyBPvU1A9y/jvz7MX61hr6RTXihpprACeVJ7emsBVmqKS/lH
SN/hoZNEFzOMuCadBLZUcHr9iZTF5ljWfrs4F8wF9lJjlqeLpHtPBJfXtTtFqmX+RQ5kMDJKMXRh
51fPmaLDfR9pFVwClJziCqdrs8YNZB2M4BhseZcKtsUZnaxRFNcdjFh/UJH++U6PMMOVC9JE9nOG
6idOQhQ1O7Bl92KSXHGe3nRtwpVjeyawNZOuKdm8ZkWkNzzdWilGUnKFbhbISrsZJVLg1lZvTnCJ
wR3hHItt1q1zJjfChzIttV64pRhNxJQxR3nQop4i+8erKXtl3gsVZIdcg51B/hvo+gN/oAzXQ3Sa
FsgVJMBk9esx0W76cUmF9MSHuFtUM2BuIecI6gQ/pRUrHHwj38XEYn+AvaxxjkYq+JPt2S5nG7jW
nNNEggnePlzW3w25cD6PlOAnzdXrDXHrTRnzRYvHCn4gxpqdTKyjGetfoIckrv9sn2+aP8InRPuR
nxfN1SrEJCud3poo5bN6x5SES39j55twpCfKQQf75vFKpB2vxtNA9y+x2yQIcxoyqGjx+gZoQzns
KHHWpSMYjAH3O7Po3cy81kLKi8dUiXRIq0IE4a7da76ejqTx3V04O9cvQ1E3JIv78w8IMg+yA2Oc
3x3y7+A7cOMXZxewPX4ECmTdc/1MDK8Z0eZzJyRHh86zWyQ1w6eUl6/ADaQWnq9N4JmVx1wxW2Rt
jLbsznmVPOW2wa2FlWTUS/5s+0TtAhVKFXM5Z+lSLeFKi77enpRTRbZSP/jXrH5co3mv9g6i96kg
T1iiPf+jD0J4QnNymmUz491QPG6/rd6Wx24irfOj7lS73Ag6PezwZCm54Hf3Xt0t7d/ml64tOZLK
7nTX0b/XtagWPpctaWJFuEG5l9tpbz32tX/e3RjHv/11sJDZQrlTGxo/dSiNS0ovLWQQ0FoYBPdN
RANNfyfBNqI1iJK5d8sz4P15RUEmNmbG3MZrtKe+rtQn/r8eyhwjRKZaNvpC3rb3IVDPVfRsHFfc
0ieo6EkuroWwlCkd5cVb2aPU3u5U1Lo8IxMjNlic8O5vxDJy+q82ULarnIaXH+8KtLO3zHF0wexS
WBLSOy54MxeDAgDWbQLXWMf6HxerXErkMwnsQywd5Lwd8QaT50+dBWSxYxGqKQ6+g/1Cwcd6bOLj
UV12pgfHOA472ToPMJFn20abqXo95x1XsFRd05hnrQgAkpanJI3yzpdRJ6nuDBAl8hh2bBnD7p5U
SDMo8KDvAKj9zoPJUV0P71Jwi7H0a85ubsqT4eyjarbRmj3wkdJwbor8nEBzFj32QdH88TLD338B
Bn4p1W8u5XQzLk38H6uLdAr/Ocr0Bs8Z2ORQZeExz7ifmm9/N3u3RgLDWiB8J2Vj+SPGZJnsnaOB
Vsq/dH2LXvYxO11br/wMZc/daFoFCp7H+p5rblC5wukLWEXEOf5+WKXchcCT/EEcqwti2XyJoVpo
oSorqp7FeElX9FZDxYfo0zKXdqArLpBYGGkL8PyaL0RmC06xQiJJjqW2FZEzJvrY0TIhrhWlHAgy
zDC9wYHO2gCRVYmZbx9b+PbCtffPnaw1ZHOdw1+27lpZ1jr5k7KWyoDVXnvNABAgamFGr7cpf04i
DpFoWf1wQPROpLONWhxWNUTcLq0LcaIuTS/Y57G960I/m3N9zD/nxJONbdm7oXKM9Ohl8jy7UweI
CRKoDWtyRNSJs0HDvDRr0JCB8C4CEPdc5Pwzi48RfCHLB3zNYXnQaYcI9MPMAP2e1MQIG/YRKFXT
Y1HDztQlNy91/9kPffAbvluLQnr8Foc/RsD7zzXjPG2A8ooqHI1DVvRgQgJODyqDU/Cu5f4uwZlk
UBYkecwfdSEP8kLsLaZTkG0/3LGv8UOHC2Jx7IIquGU2cvq3iM13vCZGNU9DqDKOhvTtd16uER6t
xqJyvUsgq9iBk0DLMM9uORv/GZkMLRrmQouyEkNCMv8AW6QLpSKB78Sd4wQAo1PwFIOxtXDesAlz
R/0Z6fnjkxPKjGTyrbxpjXxVCWqiZObxpAGd+YbYSxEuQdjAg8TXRAp1gox4QBrqTLWMO0PeANJA
AH6BfBPIe+fFiKiJAhJw4Fn4Aicdv/ftQUyO6mDyBnq5WL8UtREChg6kgwIp5xAFkiGlYa/QH2Ml
607+ROlgDlf7wMXyMhp4Fj6qEznkfBr/3X0yiD1T2v2UQCu87Bhabrn2A0kL9GNzC5Q51HEjyKwD
euRKG7Oi6DZIjpedDNLtEIL+5p79zr0m88zvy1tX/hkCvHKr1w/a6rAXt8vG9DM4fa6v7v9kG43b
91SLYLEOtxwiMOtygZ6bhBcpWnbtZq8U1PkbNUVe3lS+BLHURzDxqBBw+0CVMtuFKH96Q9Qn2K1M
uZ+jrkksfbGwDyL1uhY0oJ+evXV1P5B1TcdzK/hOGu56sY6LGpNlS95YcuWFsvP6k46sQvYo5ltk
vRnzlaLf6rboyDK0hcCT5h8bUg5aMsPwUcpqfMPG6femEpveUfHXtioKhZ13U/0ke1e7C8YKkGoW
OrZUhECkASJfMJUs+60GYSNu/dI6UaCGS6YI0TvT/JmEavkvVFWPlvraYj7oKxZsCt7SsYeXe0gt
UtGoWX7jMCFIu84nJq7OBCKhQjs9WiIMJbuRyYBtuFy6SRYA1uYkZe2i3QkrVULVB6YQuiiB8anJ
kz1f+dOTQITVwJS83Nug3sJ3VCCLaTwq3Sjrd3RMIShmiNy+4cRZDgkurl5Of8pEuJsRZ2FU8GRH
zIpat3ltrgagrXhs1seWM+sZCcYD9YD6nh2BY/ul4+eO6kkIpAxrNHgPqOvHpUjsfn3YZ6MMSa4k
8NXhkZhlyVFbG77wsTIl/S+n7KVPT6rsunHkGET/PrlbXc5VlmAD8FkmeBG4eJa3rwrCKmmEiwX8
THrKxritN58CNNFJByvG6F6p/iKSjb5G81rDZC7tBrUSBDUJ9romaivbBLupqad6rLxeOJLn6MC4
3RsAUqfjkIZe/Jo1hvKddC7orEVh8Xo8tWv3TvVdmzZu/By4rB8sUV7u6B6KmSlh16esAYB1Fri6
ctj7uDhRC6bVQ8oGtuwfgU27wbHfCncgcGjmXIn1KhTEfBmr1YPKBj8/RtYh+InngbexUR9YzZHH
Z0JHEcE2/QAR9eDSbwrCJiLgl5Xf6Xu1Jn+IasLPdw0xY39qIpNi579nycpSKi1Y5ebu8EIINHTI
ZzlJ7wvca9uWPfbQF/s8tVzttqafaMyO7Wi/J9gUyZKipoZsp2sySpNAEOWlIb3fRwuyqaX6Ciow
8MZ9Gyc+YfyKedOJSdtptrKruR3cQj0hdF7JgGJwWO1ONR/YuViRaPQpZvePuGFWGW9KEisLP728
PGFtgmftY+PBUPcuSJf03XJ8cINsq3LL4lCx4FiFtRMD0uKy+WdyGL0qWziqfbD+/kaUdCS+VKSd
SzKMdrM5x+5Z9LQ1hbKc2m8igKBPNyIZ6nKxb9DZxctF9ahRtN3wUrb13tV953mrHvm81eu5GYWN
IpqZC3mwpkN+OpSUCw0TFfZUwX4vmVmxJuXQX3qSDOFOAMpmRIm9iJloX/d536MbgM7I2TUnZBRH
KwHz9nFPUWqFNO/OqX2jRbAxIxvFkBG06SnYZbmJaKB5ucGQwAcqBPkL5RmGsBUtkexIngUjRTay
wflZ3bao/+6bgPpZ64RsqPWUXmlCbs8T6wGyMmzea+WIAuJfQpMfUV3lKS8YYu7dJG6LrZFe5qXo
1n9Re85ACob0iaVW+v61x0mzMbM0lxKYihfpT7s5jCBif3V5RsSHGDlVBsYlxzovnhy2PnOFk2ik
qVAHf2xS9wfMmDaKRN2Jg2cI69zWF/PYua3DPhGrB4ANS/JIbrIZcc9J8sJ6j3YwyQn1TqbQf9CD
Pw0sSYtHPx0M62MbrJ1MpUyu0w+yC2R6td5LkViLC2f4h7V2sv6s+pRdwEUJO05xu/GVeAaNRBCC
8bvlI0XCXBLwolPnlo+W/okRcegMXZItyZKDltnmOLNN8vretxTwJ11aydaA/g+A5GUME+wZql9d
HD6rRfUT7PHGHH5VsHmV0xljfY9A05QXtmFgvCkO21yM21+qKEAjaBbtrn4wOegjWLrEtmgK522k
ANB09XvCpRcr5Rh521UZEIpzSnAKN6rrkStVKnwhdfwyF/anE1ciyLX4EGDOWozluQNDlkfpQyBo
QcIj52kWjVqEvZhNNDnbC666wCb1Wt8IKxTpdH320NtsrZTFhMwPSJH/2XdHb3aWvNaWMl8f+ie2
niA44dLXEXHl21tE/h4K3bmIy4+ZHEW4jTz0SYHhc6KL0IgdP25YHZMyeD8R06cRMzYlUfAfeJLC
lGejhoX4ys39h2QkWmmeJDfdImVwdHgUoNxDS3nwOSmkIMbwbTF8GIvEzn+KXwxQXtpe1KwdruZP
t9F+eggdNI9inRf5z0mfiaxSzR9b6vEwbS6TY+2x3TjkExU85ZPVRQzhbZt9hMfehNo7iuG/6V7M
EVxEWS5NsyhUZeK6/YckyE71QgFx5Umu/0SKIPtB8XTwLV8LVUZeTbMIwSHD8AnE0zUXYnk6gdIJ
1JxX72Py04umv4lvrxW/PfQZsjsVtHypX7RCb/FDuHk4dkjwNhZqKEGmpXN7HneiNkTPbBLuEkMb
pA/ztREd7vXZdAT4FuCZqDxPgM9KRQQKdxD8drNJ5wqrRp7+Fovxhoo8hCVHk8qt69v1YlOphn1M
xAtVt4Q0xw58JkhgngYuE//2KqpIRf2zRC6dX/UrwVo2Yig311uxNp044OXyU06swbAAPRHAM2GL
FMafQtLiEa0s9ghy54VgKNExN7eNRg7lTqHwfFcanAxlZzju5NZWy8B+xQbnY1qP5bHXL67tcsAL
/wrokrfSEi7BppGjh8+vZP/Ufksgb/1cqxS5F7z3Ye3u4V3kYe5N9226DIK47gKfu3iobp8miatN
+nK0JhfvkNU2CIEFz0rlItwa5OJfD7PHQ0By3BuxXIf2ZdThnYNI5f5ws+EdiF/SeKphdrBk0ARK
cgbQ5865mwwfxFsXEoZr59to2sF6wtrzmoKQgCkMIJc6RgmN6RU1UGA6ceD34H/Fpe0D4n2TSiRJ
fUU+Mo1P5v82NDIn+jAyzKcGDqyvkgg77t2mt2erN8+4PVP0zVd1VQrh90Iucw5oV6d2/kh5Y73o
emwj6Gq3/+ifQHLHFb5Bs584F+AwHzcwQE/2z0w1N1PW//kjwGdQ4BMWgcFTH72MQHWFpDUiFbW2
Cl9EQQXK7OINEO1UB1ikGC0uUw2ZCtJ7kw2fHE2KqxjxF6kjlAlJTwH+nfebLNTW8fBXAvlhBIZm
76gspYRkHU7697ROCmaqkP3OOx22gsCZhEmGMxB7naHqDhigyTJ/H0nMcKTWNu7xyaL5ABz2r8JI
vdqNwTzQlRkJZ3UorNs8qN+ECMlinIu0P8NktGe+6DFtqMgzpeYVR2BJIY2RdpymNC2KxBtQe9nI
MLH60A9TP7Z9W4tzK73zqXJ9MzuMNJp/CIZZ1Ud26zycsTWPOV8Gr3Pw6ep+oYu5IJYSS/Of3Goa
FRk8Um+qkudsavokusSrFUxYlmoR84ZKwA9pLGAy2g7yAxOs5grEoeSg5qOYG9pbH3wvsNPpC4aF
hL+ksDMsi3O1w8vv4uybHmfPnIO5XaJP4LWA1IdPtDDbSqNK002FNJ7pVLpH4igoXDBWFRkL3wk+
9drSoithH248+zIszThS5kdfQV9GNuadFjJzpSVee4fcKBrJgi7SgLjYR1cpjvC1WJnxNywIxH/Q
xuXmJW1pBi6G0cRmwY6pBGVphy7KdM5dT1T4i/L9o2DKFuG3Uz6dbbwDjxlxn86eon/Mbijuw23V
1YTCkDza3lijEKRta8HAqR1i/vTLohhwVCOFAFmJfU3+qxf4DTmV3ZiecYR5pe0wb+IC3prFzBUj
GA+QhnzkzttIs/xN5wyVwSvxYDw1jZInZhHnkfi/AGtoWhttL2hObmsVWSXLlyF/SomCGEMpvho0
8KdXChYuMdRiZvsvHHsBG/OtOiaS1XO+9HWSmRBiUYH9fJGHNi6G4JwtmYMjOy4uzwBHMQtW4ouH
h9OQXBj6drg6mdSLy2n24qnTnLa0I++Zidhq4iDOrGArAU8/esnF1/yEcPhbb6BCYLorqidVWGK1
tnhmCse0YSmLEf9Cbm3pzrzVKXBRmVGQKpRtdLFEEYlxxKqL07ztsMuPLMNae00TLhvABGU8wfRr
3tO+m+qe6KQ67CAddkC/6SVVy4fx9vDQAGy6yOTXLFrgZ+rShqa9SVT/FboSrzpMi6HFcN8cd+h/
CX0lhbGvHhQ3kFj0CDReacbbk0WTNHCA6cBnZ745F2mOLdpaqR9MDsxLEH9jhMcNHAHsWRm5Ipzo
I8bnXhkzXXq70B4TUBvMeOc2gsuYXFAkKh2uJ/MAFtc9+xy8oHofVLx4Nt2wGTqwhql1PGvcBqpw
5siNW6xSLAD/U+ob+one6UwhfI7+PD5aQGyIQFO1SbHBm3oVVbDx0WNKM5l/bblv4v6tI8vHiNA4
6W0W4NujBxx3dZ6heCSP/AqK01fYEv/o+AgEDK4iCNXjlpdO0bfZrIPXtJIGli2sNp6hMa/pXXHB
RmoSgKb0IxWFvGQG59+CqcW/uht7jrcE44pTUEfyTFjMKP1qLfJv5ADA87jCeXtwYl0ckJY+ykVd
2NLPcJAIFKes5lXJD9Q1NKI/0TWIB9HTvf/v9JBRxG7HVSOR6cwpi7DmSk9Ndqg/LAeiQFaRvNdU
Kyx8erhvhpYSVHL+B8UC9RdnkzAUHYv3Y6YFKa4sCkPIUdFqMWsrGwnrg1KkIF6Wu8tHFyC/oOgk
mdCqO9xc2nGqTqJTIbGqT4Ya1zx/C6gYo1jtXX5yNr63cXo5sRpJHh9PAnD7DDkwjtB+dnDA2fxo
1fGzIk3QutcuslTiHAhxdWJku3cBB0BYt73mR435WuyAdz+6X4tjO1KKUkD3V1CI5Q37kse1rjRo
hu5k5G5osV4ifYgx/Xm+XkbGswNrsmC0Z7h/EGjcejIw8CYyaouHdx2O/fH4LSsxAIM+dZveDAHO
efgglWIXTZJfpW58IwGPMKcwAaS0sdhaqaatDStra1XUnALDMOQvuOE6ZTypXcpOICNTUt5tUmZ4
Va3C8t9hZx6IF7lLY6hL+/Ew9v1g4LbunWrvduig/v+DsdgKwrA5GAqQ3zFphrXwhohazOeQpKNo
R8sMG/PYKzxWCGZjpfPYoKyJDyN3WWy3LvANj7O6Ko5yxwWg2EBXS1U441eQQqefTdgQCaOLeA/Q
dRNvGmGdkolubww4w3QPkTDxSuoH7mTJdvItVUelpr/+0flgd708L1kJubViHMn0H3Tut1f98kFu
69mJ+LL+MVo1htfJUj7dRfx1krZeGDbxwN50DRnkcUi3oM3hTdWIuSsle5MVeIifSxVLm9GYxQmw
+GAulbXy4IcXxZ3qxBCYybQSBk7mifYUCNndytG9XpTzma9NU9g5xZ7YSfj/Y4LMs1EAORQUWsVM
PMg/v6ivLMzFt1roRGruQEfVBGPyWVuevhrpejya0mDGzhF8UDhuJ7Ij9AkUQOtnnboosql9acbD
+HZb//c2q9N8ve97SUvt6Kaeci35cssXvQucgx9JtPoKltfPy6ps7k6a5RnQZXiuoP8Mx6Ad+h0G
ADBsOQr0CCNJuD9b2eAVLlpjUSJBJnoZ8yypwW4FXzxpob+D0yHyO4zs68iGSABjwXTgCN29ljdY
VnE75bONHVhr16z7ipwqgqZ8qB9FVdWALWfn3+nv13+cCOiE/jDTbqKv/Ap1bMquhQEq4ad44ei5
r2LTXhErH2zl4YRm2hBi1C6wieANjFypvDTHddcsn1g1499UKIThFGUrnJyxZutdzPe0paoowoEO
fxhnabBF2B67uw1YCR5a0Xv6RvIhauk7+WtPl/wtj6aQ6wRxR5ki96QcRW2ANMxOD2q/zk6pkN1u
tG52uejsn5TziAYuQx/5OJf8K8wgu0jbiqG3qQ+4VvsrWyreensmKGHwZVti5fh67TlL5DWIBlOO
u/hyDrNnBuDfoqaDuwqO54kewVrqpbjCMI62E5rwa/fgNKaApO3Ke2Cg/NNzpHZS2aMVFfezOcTb
S2CmT1LXkQkzB9IxU41L6fR7Pl9uEgi/QVj+MD16nvbMDg6Wjnxvd7PWzZvDreDrIX+MI21xm/Ig
YmQ89Y6WKjXyI4GPVH7oF7VasKzv+yzv1d3wusBVTURE8cvkETsdf+Doo6+IyiFsXMsxcDgK7O2C
UZzNqq7TFO+Mb36DPmVrfEUK///kSqyCcFv/dfGWsbXw22YoM2z+mlRAAb09pveMvGidpNhtSVsB
J+UjPFYzVCxpx8CDPJZlo0sWqNcpRiPYgJDK9QfKx0gp9CA7vMdcb+6Oqumf2BTDMMFks3JLVmLq
R55trtFugnHy8aPmCrLA5bBYiy28gy76rTrGnLyuQknzuWNsZ2h5Q8rW31haiHk7H9Gg+Sjf6oJS
4RYbx9w0wdn6mzH5rcVbztbvmUw1tyYFF/Za2SBxy0s2jhOwcJzhdW6m7fEUTKsDYijns7YL64gI
Of308wI9e+eWaUdsKoJKxLBXD50hwJHEqK0ZZbUNDFxyxfT9YDb4yV/87U14ajJLrj7Qxkl2NjeH
JVXw29zQKIctMP4FI2nWUfLWprSMBIdU9SEosKMVjoSNuElUMqVlqPOnTIBtP00QmCP3GMCEGfpS
eojivpwDSabxv2kW7+ty4KERGsXyXSB2gaPq2wp+XI1XcXS45f1jlngFe6KgWI0Zr9Ma5rt9B44u
vVuZQ02VnRhQHDRj/+U9fjk1l5tU5C4Imc5HVo5HhBYSOTE+ATdHYRlEl+8aYy8T5Xt06O8Z2Cnp
g5rEpmDwBKxXrzWC1ze4nnUCdj4qLZ9x8pftYLvq7gX2IC4FK5P7ouF5OdUl53LJwllSWbnTGaSc
LOfadU9dtPJFtjPaOoc71iYgj572xgF6hqAw0Cf8BLBpgkH4VYB2T8SvxjLsliOscwuQpyTCgyIf
TXswarpbPObwutJl8pZeVviGXrfHyb2GVoEPV48dYVwNK8LZ6yhCJQrrXQUncbUoFijI90atKWYQ
D/G2k+qTEXeuMrD0zuoGbztEJUx/nuZC2QRBpQ47vJdLyfmAbKsJAwrfAV2HsN56X416AUPjKHK7
TMOd+x9cYtWfysqYN2uLxduQ99IQ4yRTJcLRE9Ey08OnmPYxtwInHu0ktHzc0yAJAAPRI0SEYhG2
NjbxGEYH7SMlz8dEeHPeHXLLCo2lkBLR5JKiXZXFcWXoYF6O+WVorgWKVrvIHDy0JSqS2p+1DvvR
l3MAJKtPDiKyAPNyzOucQRNwoxUk/chkZR9IF0CS/cFXBJSOxjeuaLH3pE5nn0/qw5klPVShoyXE
Psdxdzalahx6Z4qvHJieWldguZu7vFi58nSqkSzBrHyP9CwleWgCI9C2HgUBSAiszjtn9HopOWnQ
rvbX9AMM2/5XaaJiT55/MHKv3sF9rfkOVkN9gFN2S62uK/Jw5KxbCO05Y1L9hpvD/yRp3AxH+0gr
+HCLxEy6sd6v7tNGjdTZ5vM9ysJ4Mxm/Y3ruWQGa+vjVL43OCgc3TNRBWju/Z49nSIoqOgsSINbt
wFkHQIR8ZJf35fdzU+QM57t0P9Q+KM5561UfV6fB1EcRm9M5orkv5uXGwccd7P+04Ch02S1LAvh7
wr5zy6SEX5e8Kve311kjdeeAwtcz2Ga6yYbvFtJEj03irdqYaBdQ2Ng5YLTZl2yIpFO5UtKGpral
Z23q60Y9IbkP67Y5Ufe6moctRFsKmKCxQ6kjSPeelm2t6pLzeICYffK3N14N1oWX4VXHKk3t3/Ft
2Heq0UkyLbQbXx6SuME2miyZpewxSPX8zcyQ41ZELkJUl2q63JkstayjMi162CcPcWupfJA5w2AK
4Who3/pyCw6haT+/jATlPCbI9/6za7E/1/5iuMZnX5BoZQZ03A3VPltMVsSPbmKZpoQyMWqPStMz
7j+L6QunyPQG/wLSQEm1DE8MH22Kc3GBO1EmVtRhTRNe4BgXGxKft/PiDJFiMURKxI2xDd93eRFQ
OOoZ+0i4NyBB9T9elytThVggYtQEN8hIuAUGPVYVdgIX1NyYa3pqBdbtc+XxU5Py6d2VLE5Rwfeo
7/al7mr2yiFIsI1pYOIaZF00YEOuWG4YLWBXK2KtCLHb6SbLGSXOvIC8KPPBttZ0MClJd9GXp1wj
EeKE0YpERx3iiPYJfvjfYY/s6OmgAyXDCxvV/nD5C3pSzcuHOxYsA8VNkokyLficO5MsWzBUF4Zs
52uAI8Mb9Zmu5SL2ufkguDUqbE44CbiIihVfBo499JEUBrlZThMZat+Fd83sPE2M8q2nHIsgFQkr
ce8vRNhlmx2yHo1LMpXNzGuBRxmHc+Up/hEZf10RZoCMj1ENYqn7OCCW6TlYdLoZfRJPr7OykF90
fvN85aXBrqLUDScbakdpmHRZmhYERZr2aTV7/BShGaxawBpM39hPOw1wgHSdCqFqd0QyBb+YspyJ
F+BepAfEzZ/oCqxVrcIiQYNEDCzPCfYSpW1CLY+tHcq9EU4KtrM27o6NJ78HzkUDApJPu67DcAgf
3MIhCbsGM15CX8kK7Z37cTdcqpS9/XUimcr1OI131JuSy51Ji5opVGxoALhFf6ht8ImGqc/qJSQ2
qD48AQOb0toc4W2BVEU2iWMQt0dl8D3JF6NHNqXdG0ACf0O+8tWKJXBYGUUY1HDkdnxbU/M3ITpz
ofYAQ/xeEhp4E6SpCagF8pst9/PjdgijcWMhASENKgEKvQ4pJSBOXoPjVF35qjaztOBZx8CsTg7r
t91UgA2kw9z0vmleVGiFo9fVCmZgPFL861c7y18mcn3aDErMebT3UOwsosR2LFIpw1/fXTbOICi0
SNQuHsdGYjZBOvLoMITHmJGaXKqKVQfyuCtD1K0yhItnpSn9m8M/kutjDiexKu9qfVrmRzsrY1aW
tVYwc+TbQ7tu7nGb30+SzYyi4S8I4O2x7x9x78W+xTfxiLjxLCEktgJWMwiCZh3m6Fjb/5wh1i2e
rZY88+qK+UALMOJnwjOHupoqG7F4OHziXZdaDAgFG0Pnc2pLiH7HVDXCzRgurDn+VgR81IQfbDH3
BgMCirNk8BMnrp/ya1XUxzkli4bN3m2FrJ6nU08T0AbF0XNoAEaBjoAP3A65HDpE5KZ88O3Uhm3y
yNp0ZfDx6FdVu/5q0fXqHOGIvSNBhJws6m1jN5KnuG0KvaVGTFG5/AtvsEo1ENjPJ26oAtdI3YPL
S65rnWqWNFx2YGeC8MdUmPBp/gilIlHuVI6fP+3ISsZS1hSegzufbmUDWXLRE690nC4JCTzlBmg+
QixDdi5sUAxEfX2ZFChQxjwD3uBuYWluhNVKwCpySNVO3l9QKnal6n+Xjxz7PAypRVRflxAw+58D
hqaKcQxdvYE+KoO7GJgwsm7ZjXYR9cU5mziY3eBOGZXsdQR5FTU7fv4YeL+q5F7EAAW+dI4EAAQD
G6NF9nAMGpCD+FNbzgRjrcXHaqR5F/U+QcwBS4yD7eZjppT5IPvWpoJwJZ0UwZ3Db3f+xyX8fgNU
9FAV0VGOKfaI9olqXMbXHIZd0A/Z8eHD+qJEjPnBZ7dw9RjbvuqxGFz/J/SW+vgpT+z1LHQVmP5o
YQrRQIbjVB+HVX4rb04ChE686/9DGabSRGF8Xy6oMT8RvnF3QQrpW07t6RGCcEdiGaOUzMH/E+8k
CliTdneD0LvGr59h1lrunf3BaEnsRY6fdvMfWv1WVUyUiQXd6M0MkPyQzX6xWnwdUrLQTa7Irhsa
CVWO1RUa3ZCjuZQa4W9pWydlNWRkHIsbQ0V+SiFdkEagXi/ww10SYD8QxLooklO9lWeKTNX7Zt/g
/AxxEITRBbNHofJlXrEFRT4S6rxFoobV0DHjVQbM6EsQijUYcybUUQ8UH00WUc7i3QBLqV7CdbDk
deTSOuj+0FRr7T4R1FdPc7YSUWxOqVsgHCvyTtZXy98kbFHwyO0r3OJ0L8gGORBwMl+/GTCsnh+7
iUveeC6BuqYMkpaVXNE/APxJioyuQMrQ9h2MMUdMBtt91t5eRLqT16Ce1vp+pln3fkv+RsH05z/m
pF7nPrMuo5BgwxzlL8241QkvE6weCZYBp488/CF7S05RpT6a3pOIWT3V0wh0adPTMMzj/5JvyACM
abNKRtKrYttCRZSC0PMuTMDlrB6gBAvHiaLjbblCCe0lqWfRNzyU3z9ZyjjVsw0hLXGtS1zJN8V5
YORrsS0FHlcWEUo0yFS4TwbLPM3GCaxOIzziZXRLUQQXVw+8Xp6VmgotNsjSy3loPt2yZi+KxyGG
pXLHSANWkg0dMMgRr0Irb8ziZX1fIdKeJRw2nng7a5czhHHeLuvtEAHiRcY4nPA7i+qtf5RWh+9l
JBgnZOB9R3ScrVjuWZ3AByUc6bpmsMRH3t2b8Q4o7hS52CoG4AnVZJvBf7IQop0YVk/FYKRkqcda
KwxTCCDoOF0DrL/UmW7ElrJnbDnYyXM3lF+mHuwzGaVNHEgVW0amFgjQZ7bjZlrBkeP3+ydA4x+/
NRQryv5qE2+r9PCE97NPGARRh4Vw6mPAIn5FNHL8x5kkKJQP7qFFtxOvrETRfwOHmeST09EUa8sk
J71F5ti5YUSKdEHBC5MNg1RFyL105gwZDPZmzGgmMf4Et7dbwG7WrpVLt9Gl440CQ9UumAaXP4Xn
+lF9rhuj7Pv3IDm/LxtEdfndwTxawoVoy2RKGgzG9RwYUJmfNlNwdwpy+9OnkEywXNxFiPrvBkzy
l/ToGWULTBZi7ghdj+waNUDcZryd2j150Jv5wRmRd0lbhOd6uS41ZDZYe4i3DHdoKD9pTrSu2H4k
VWn4kNddSieBp9pBePSJ+N1Rx104Occq1zG+uqQOXSpLAOoYtEIXUIEkOQ+wAzENJWOWE4aq/BTN
SxsWSqhls4J/+lRTmwiktiR2kOEXQuMrR2rAv7qaISZSDYrAIMm3S6OqtOx1rpg9rs7nMyjhaLB4
3vgiNOOqJ4EJ+/ugpJPFav/ntDvXc5FL7y4qCuHbhJNuRN+c36QAmC6kwO+aqyQf1YFrvEzCEzcu
+iRx6/qkarnGLM3UKfW1mkPv2Cj8xRJCreMpT4yjZdFqueNrSQTukR2HvgWWWvnBK6JhEMCe270l
pOS81j9aEO15NOUAg4vxu4y+virEa94UqOldcsRkq64JoEuefXgV3y99kgwQkMq622APEZK8HTok
bbZbF4aXKOxDmdF0TTWHFHcKDmSDIrhJEywGmnIjEtfgb6HO3Joc/kKv4xYeamkWU6QXCsxPcRcJ
5thFKFw3PElCt1pUcys6yZT0QI5gLHJQLRgQX31zRvdGqlWFN24B2UJjQ5hEbifMam5+C+7yha2y
TMgwEnSbdVMRS2I2TRezb2vHT6U/3fg9LqIcpRPUUkubp5Ji2pBZCUC0Ds8UXwPXjnsO9kb04Tyz
IZf8ZCVpb9MicRU3iyZTTWEJZl6OE3meYSHxfB5EdP8bt14lllqbHhcsV94woju2Q+rozQKbvxUZ
R7hHndkwpXAq9axqwFkD1L+034EZODgMZZALZNAylzGQiTyTRcQl5/1mDbV5/QmYqwGU/F2WJ2yr
01pFBI2TBe2UxsLaSW2FXs1Nqu91dOLLXA47ldcGmrQyCNUQJlkvk40e6I9rzAOKaZcrEDQejrg9
QuBaQxwy43afPK1MRhBat6LtfRIiX5N7C3Oyma8hNQ+Psxwefs+hpeQqIDa+aVUDWuA/pYwIc1tj
7jYmFR0PcbbTLCdEVwlrlSnJRNVxcHeNa1rsncaqXDYGE4JjLMx0xhuLcgg0pFzgGGXppqrVMOdF
+CqhaFesNHDTOkFwCi5EtG9Hv6UYhQpPSFz3MBBIiae5dXQY6+enc5xJNbQKR3nYtyF4J5200rTS
IghH6NTsOO5367+jL2qZULCUVSU/zckm5zwLxOHPIIceUwfjVkRA9xEX+unuiG9yYbmmWxX5jMTN
aOQksLx9SdXmTYa3ZlbGHAPmeLt9W0G3bbKi+UQhGgfmR3aWxPH56J1Q+Zobk1ztiyWI5vwCYHxk
r6NpUd7oC0OgklWu583pAi3/9xP+LbiWPlBLHoB9Org9HxGgdH/FO+QlmQiLzXolvxknM0vJPYzh
pOVIoMagqgZKekB2ek6DKDH7juY1+qhZO+PQ+3QbuAcPKUztEPGgxhMIbfDFkQhUwnVIUz4+D2Qd
s76P6QpHYG9m7zIJQUoN+0jk3uKw/3PY0e492C+aJd2oFV+ml5A9DxGLVxIfTOUjgAiLsRHQqEtt
csM0t0KJU9Nm12nE5hBwezg1OviIZaQaHXaOwCgWPHuCobiU+liLAYO6V2MayyiLBbz2ttDou4X/
ma1oGZ3ZXa+aaW4fYaVPd5JTfLE1IKGoW+GoCBDNml0iA6gOUdXsy0bofwawOrK/9h8O9sBreDIE
Z8ppcD2QtbDulB5RSbarMoVita0UsxpJFvRif2qjzxr2p8nQbDslFdJch7K9W9byanJmnTK45jce
rqzXMRYUQHxfelsdb9QXFp2kYdr9LUL4NJoXJT/Inf7+Zi/SEhu9bNXktPCJFGAUja2QASgUXmUH
1RdnjLFo/nasBDl6nX+JZvtVxqlYHDfXv6fC5UEtbYvszZAS46oL5zqLoNX8R6WtDohe3dOPuC3O
ateuPXjUVCpIKII+TARwt+GVrX46BMwr2lcUyZ8QSSqK5IfDZ7cnG4sjYzQUCQdTng6+20ImKopc
y1bVjjg5b7/iZbV7n/CT7+lz4YfhjlY4+AjNG0kMe+QFLKCYqGenOttRT8vP3aK+JetS3xB2Gk1F
SHw9wz5eeyUJwcxYtAiaIMXf3raydSb+lkFwPyKVPj7BlwTYBOXi1v+0jIWOwp4pMBuSTMMesd0p
jnBB4bmiNjk2YS5rHfs7kCTktY4fDxUEc6KLh0v5DwpIQx/TerR226PE8hlKjRPNUqZutoE0ARP0
wpp5N1K9EdS3OaWXRPC8lIo2JSAJgZ+Gzdz0La5JPEyjVejnU6NdMcoHQntIGDc5zF+8u190dYrH
j+hzCjdQdjoU94KRTzs0kCIacPTDZyDH/Gdn+J/l47oNYLLS5htkbaDjTY8XwQlN/Akrs1Y5OSO0
U6HqIUxVQ9KPxIY6KTFI9cbs/PjYjgwb7CtwbVQ2BUWwNI/TrUeypa9xFANoQQVkaDNxyQqF4DX+
jwz1dbw2qS9V7b0ujs+jEE/iBVZZBPLK9xkWXyVOCLi9c91LQ8wD5BUQ+OTZI8tvEQFpgs4aV9xA
jac1vpXd5PwoXMWC8w0FESNx4+1knj4FG1H3B9Pdxdnb6esyyVlybs0j70u/aWhM2W5IArEOej66
UPhz2vCyRfWDjtNmsjnvjmtT6HnQISaVCYMGwfr3IjxdfNM8QpnC2vECQ67psxYZ75x9Gxoe9cbu
hAkvhwbBH9WCXGclJcVY7tVDjC4iaIibqY10SNv3HACNVOJ4sveScHMJLP+z3e9EeXB6Pmi60GuX
d4pmE6ZpQZP/d5dHoC7ufgk20CWAYdGyNvsDo38ie+PWnXsVzNuaPFvMDfbZhvpmxsjVAHLn+yuz
B2mgHxNeWSf0vwZ49YPbBg56EjZP/O9OpakFz+sj6Ae8sVB81tMKApdnoH9Dg0zNHx8oZ62aCiMQ
pwJbM7vK33yTYs67K5rVE654k2YomoKO+R1oVHjIedj3BC2eUzHjJHDFk4IS+h1aa/qugnMhci5v
Gp0Ee5nlC/FWFIRODq5VjwjzfS2stGn4qj7C0pqJwXeIgBtOtprvdWFU9hrD5wdgj4fUY+78hjXU
pygt5VdiEbmggZ1WqUQ5VpcY0odWIqS9qQMGE38S6DpY/64+3zPOIdqwJzLCZAZK8vt9OPb02nJn
Ex+DhQGeOZsZAbCXcY0Fm5r3NpbI4zd9pUV1kfyCiVrHO2Oe+/E3mbi7Ziqsm3XjqqKKnBa2r+Pc
LZv+Pld/SLTmSv+3lEEfBAyR7L9FEtWyWyyy6L0zmu6+igfWJBDDt7oI0mRYy8ouRrY+9W/ibF3X
nvjtWcTSCMzWo288uPGrLNRtNmInxp2LPjE0puZXh3NEciuSF21JOq0K4Wkj9Nq0R3WVzrYnlG9F
eFux/hacYKD6/0Cjw2UsLJYFG6z+3GjEtTbWGLe5f81TLcuE7PE8/A1PxOQ8TLMpN6g6tGUCoeTw
FZTPNoVMViHMjc+qldOtM8mvikMkvMJOv/2MHavvBqKlAah4uDOhISPw9p6ugcHNRcPmD5oCXB41
lqqe+jGevya3NTcWgenTHluUomaWUlpvv2b+6cJVLlqe/+SWXsvIx8qdlPoYsA2a/TtfxxNL0BDX
wWAN2zTCaWqH27bXhPX2EdQpycltcY+/7bRzow9FFM6Ft7TVnPvlO7cTmITgIHgzI6zEeWtrAYX9
EtsPH6+HD4TvAm3Aprrqr41Wwdgq4+7Nl+uP271r73D3k0v6J/yeFpFQc/wIaBud246YbQh6z+QS
PUx0tv9e5A7Jsd3y8reRvCANF5BaXFmkfWdU06FjmoCEwdujI0AuSxb9tPR1LijCns/RytvruvNx
NVnoCYaz2jsiX02wzbs1gl8JAQMf4dxNopp0QPWm6ICQFHAEhJp5r0QuAy8yMR/yphe52Pw/c/R0
Tb1jFD1wUsEZf2KkAXJvY5pXRdgHE+nJlxNaqL+ypTQqvh6FBLCtVrN9i+VN5h1veryRGqvRZiwn
e5KI0/gx241jJi+k9gm+Kh66jhmOadXOPVuT4yV6EKq8imbT/qVg+jQxewX8qWFmmSt0A8Rf5STz
PlvqSlxosk8qu7vxDGrmpO4AeeYvdVvpsvma1IZRxxXRW77aWAI9L6VaOmvReIQsytiQCLPbSCko
9P8X/UXFh0tqSsEhNxNBa1khcqMhd6vq7NhFFcjuIrCyuPdbv13gxhCPghfCvESfxM+YEyOIiTU5
0ExJLmcCwZN+wGOzsK8cfPHCYFxVIuVVfTrW17gNZq6FXzlBSLuQ8XJpNiU1/vMgycD77iTlxTN8
ruqAm7c0afd3XlW7eNWZfegfae+Ti/64/81l6HeXV2jFGY5YQrWYZJsxQUcl0wfMRCr9ettP1loL
GlLekVsWELOLr8enVNAlGKlU6WOKksJWLJGDE6+nwkPNIFDsqRv1Xq6n+xSwk//6/XbZHmFBje29
CjESUR5npHphUjnscqGcjtApCQ1WrcylLXrTF5fZ/4K0gfQRW1Fd22Ky7SlIFUlWpTt/dXCm0VTR
ayXNBD/9mbEjqYrKRz9BJA/FeDu/I2+22SglCbYJAQ7TmkkHbOxaoxz/xp//wTVZnZqDrFJAjEb7
OHXXFyy7YNi1mB3jOLCUSLKXE43G8AYMWr7ocW6a24F6mcps+B8ua4TggoLmxrm69Nmfl7hxQtYd
iO8bkvOILZ/zVnz8tl+jx+Igs5x4fK/x/rQ0gAmzZpv5qoz/NTcaT142q6t+KCk5IvuJIYaKTzG3
2YVFPwc3s03YojpY6juOrNiaGbJ2tkDJHUEfhXBrFidC8qUQ3yNN6lM4+/tZx1lcG9ES2WXhrF1I
dQrkcCEagx3nShuudPni7kgNdoW9Yj/3ExYqzr4VzrSlbiFU5ltAsJKF5yW6+/IQ0Ltbw06V3CAH
x42W/6AxXmJNgzH1Ke0QlA6gxV3Z31uo3X+9gkKaYP9adLWTTpzqw3LtoaFG0PzrXxNlU6kSuZnh
N/emWN62zW7mF+UWXFTBSHi6oCtj1Zu2a6/4UTlHE6wQEVNr0a64SmTA4gaRN7TjnRTFob30nOG1
T5ajh6RUAgGKVOSsq7miscK10qlVaGK1OkaIxVPPhZwHbKpz4y3I9ooEuyEc8VzDNCLMqrwNconR
l2y9trTXReKkElTwBeD73y4rkgCUrKwTXYWaFKPzv0a89iEXA4KTa3Oc98VEi8L7GNrph7XFO5GD
uD8krjqHJZ3bAiUFelQ3+hAxooP8sSgrVW4GVD46qIKJvOtXWN7MjNfVQVlqgjY+z1Av25KOTy7m
ImcvBM8EOUmoBONdcT1Sq4QOdcKpCTinjtiGK4TVrhS7EpYULDkdkymnTI9WiMPKVmJXnIRZPh/5
ZEs1Zl7zDxM/KI2zGwIS/CzAl7CM2St69DOoOSy9Rq55n+ceTKJw3F446D46ZlWDDf+Qf10qghdl
U9UlXhIJsVmfd4u5dXvYCqDKjmolRfdiQxq+3PExfMyFLO3Y5LBvepw9DQjH+CpvO2i1OK/gMYOH
WZPMUwYmk9JGbkpbmBjJF8KYXzS57TL/yPzeYh6ELRCE8ID/3uEYKbygFdwPi/LDmN2IuvFt5WDy
SSx9wq+0WSqk1Qy44scifGqB5OBu3fllpcwy0S8b4U+nc2iFeKCgbgoMsnroITEIK1Fxs2bvJefo
YP5cFwu81dfd1+udo2d6rheAOdylY0Oamx/AsoygDwPsMJyCuFg5EL0OOb9ourLdtGK5wNf1cwqQ
2hIyAXhJ+XUxtN4fNfl2XeVdGAeFuMsPlxBQ+ZCZtUfUuz47UTm09j5Lm+6UqehXnlgFuFTtGAMV
Zco2+ToutcUoj6aY1lyoE9rLpOBBfPndtOfzWNLYfPwb+9eo/CnloxY4bl9CX+iogiFJYmaADlof
t9OFeu1I0s2S8eesgQH6XP2G7afx5w63W68sr5DwtHuIV73Zxid80EjDvMVEcKCF4uaGhViNHBsZ
zfIX4Ve4Mt9oTXAxsnht2B4R+rA4hXECVvVb5L2EEE0DSFb1xRBtVTdiTvsd0jDfyOFTh0U59TVP
m+mBslIXdKSQvTnP4kkzNAkckr/eUkapERMoFp6dx4pRybJIKsijY875e394cf4VlbFFa/f9LzGc
pnhuKy307dtFe4/5w69XUj+lzrPykwhRcydppbcFvlK+DLKmk4pJQsSzttQ77YCeArZX9Wvn6rXj
1DV1wTy7thkYiPvLjI3yMKlXPpgmym5qFpbPD85VZIKgsM9ScVANYM02NOsuZdTUZERiilbHnuNF
93CPk+8PgtU9Tbg7vkSrbk9SMukg9j8VrlIhejET2F3UtOpuUq364PRNAwCmrWEKXdpbeTIiOFMx
rRlUc8XHIqMuoQlvfd7lOfj4J2xuqN6ei8xEonYql77uQYL/oglwwpZE6t0Xnm9nbcuVQ6TDqXyx
9If4RM2R5antY7qGSsATjuJKfGM3zklQ7m9nRHamIrecftyXiPYe+1lkmJ6Vg+88S7/N7fw03tvA
gfSkQ4OVjL72d3JMq9SpFLbd7f7K5D2rubTLFsWYSpAisbDAP04t6/OFrIm7HEWulDcrDl/1eZ+E
mKwMrVkZ6q7n0lZC0QkNAyLkzAf1LaQk/QGru7QDG/n8/0DMiv1BPq4Fp9cR5Vdx5essrF1Tf+i1
QFNQUMjAzrZ7xiQiNXhfwdHfoFYenaCtoXH4gw6mrKu1O5RcAR06L4zoEGAUctv5DddUND1gFbie
PHrJpQQ7+8RCVMNj0lMBdWE0SZnQS1XoTO/oLRlbiXWpOtDRCoQ+CvcqAPP/Ixof2QwvCez8ObUn
UQ3TXNfzPdtM7Cb2S27c6vzE6ClBoSGZdRoedfNCasA0ph/DQkk/Hvpry2ChmsuhDj3t/jnu3EXj
NeY+e5U75Z0ctJz2RjhAC+aFdmBXm/dORjpwKrtZv6w8x2joHbQVpFyn8Ri6OJSyAWhp8A1W6rYK
kw1vs0eVwEJtP7Jk0pBLsHc76ybAx1ThOfN3/IP/Sa7IQogeakln9dvpwOBe51Et8Tup00PCFNfS
eIrAxX+LjZZquWlHMRlelDueTjLEN9JylKeRqeaexgEh6tW/qvXkCKor7gUm8BSpy4tIdKjpDpK1
WeSM+L0mI5HCm5cwTwxnSTJzhf9qqGZvEhvmkgDT5EmIYHTbmBCT9l3TLS1KH1JHfe/oJUtEBAej
VjtusWBVbzss+yJacoRk4MZ00w6OehK7xA6xmPeT/kfLeAUKDkXECdTeqT8HbBISC5kHrDkr+/rB
CgaMBojJSJqD0IJ6LTaKqI1qNQ9L3EI/WxfEH+PGF1aEHs34INKCcC3OufCQNdXhkm+Tj7eAGGiL
Df7QEi5XhN1raUpO6emFG+3UWR97Bdd+m9umqOrmZGr8ondFllYLJHkHhs5ZufmkMiZVDorH4k3/
ArHT1XPpG2isz/PCBwR8caIMrw82jxNYhZyh5t5Bzp/Rx8LNSKZG/v6dJC6uxJ9xC3/SMATc2NFo
ZjjqPIkf9F1dynaSDB82W4yw0VhqV4mLCzmb4bJAhbLJhWorQmBZvkHL/BgWVtk2GjiXGBJHZUcv
7SR+xiDCxFgHazsreDOS8alka6ijgaDPa3l5EjTUlO8dsNS6z9Qg/U1kVGX+56lhILVF7ksa5zYk
09J1InHsCTqRGYgpPRTvEkxO2lO++MHGhKA5dzsKPUy94BMtgyod/ryEbEbS7vEafMlez4b7bYN7
+UiftSqY4ATxTOZVG7XnqF/O4te1ydS4HJ18baAbiXgUNBEc8MNd+7TW5Q/qwkC+oa9fqnEBfTWz
l1gposaqSwdmRRfrk043zrZurNPPpyYAn2L0fOcpRSGTeBaOkIik0Mh8ZFeiMt11o72l/8i9w2b7
2NyPCe/cuHCtXvWtjnlJaQ/A1eMUvGre+4NlSWlgMYJ+3jRzb4InzSyO2x5n/IhBYdg0f2aYXEt1
a85rThzeYzoImEiaPx6AK05rg360pFvKY8r5tJoCZKTKvpndq27IStHCQn4D+JA36E9ract1lFKu
WcmMcC5f2gvw7RosNa2EJzQNuI6QoPd6vAg6ZPxwgta/SnTKode2u6uw7YqJwaxpeDZTPN7ewdkR
dyBHedMz1IFfL7/8FZSluDbzpEFd3k5UUoWdZUUYRDCHFgpdwRcnLmxJWp2Ad07uhKRDj5Bfg8G1
+Mo6p7/JTTEQ7mjEQ/Ub68OTPQkA+1qvp5CXHn9Pprad/3wANlm7Yw4EGN0T2DHs3QsPmgbgzb+v
r4PX2zjmQy/6F10BPyz/n/U6XVKgPOt7M9+vlUrK0zdRoXH2cFpKaj8kGkPfI/R//tzuh2VR4e1v
jznEID2Y3OWkPMstWkoR43JyvioSWmcouDKRNb8D7Cb8aWEi5hu4mOyUnIdlq3jQIcWJ+NHzQ/cC
oNCDXncD1fZkTtfiFEbfG0vZdis3AW+kEtakVsTJbYVTo0gOFhKVVn0PNzFC2TwLoWnzckaVKyDw
GfPx+kJIao8U3koA+nqwmC0DUU+Hc0uGQsbLfEL9kedSpSv1hXOYrA5szsCRABsDUyn0WNs+ubix
DFTGXU6n+t85cX+aLnA1lO1Ac30cfNMgEO1uRD3+809w3N/IuyucOI4yezxNHmbs+I+f4j3QytXQ
RIC0PCwfld1U3Q9NkCmkG1pRvZ7tkk6yzApRcR/F+bzK6CBclAIoQEAws/+eOdR2pLTzqIBsHslw
o7LEKnq9mVrWKaDq95S6ldgCcW5RdFgrfpNveLVQNt6iITvRRxmQPqGrSDQIPnUYXdDboYXrJv3t
RDE27wVzBFeEP81AmXEwGMi/uYp2rQFLu0QbWsYg+2ZV/zuERzVU6OvZaP5NQwsVw1iiw6Im01sv
chOJMi+yN9eONc0Tn8t1gm37YJFbzgsynV4IJeKsK7nfT4p5/5tz8VKfmSu5JBoazGLjc7awNerC
UpRze1c7J5ar2XJKfvLUJSSNsMzuY7HqsogqA4RbqNRFaA3azCWAwkoNx3K9zgs+eXqCaAd0037S
QKa3aC7IognAXJ4U4o1oP8F/t4BtA2Ouc6rWSYslYiB1NFNXje4RKZ37JNY/4nQg7BEAeOXj1yAr
eSPMoMYSOym7CdL7tMjQfllpqARNRBNXYbXawJalczn6JFE96QMedDTvZaVM4Wl8YYQt0foWeERZ
5G5Dvhig80OWLZkQXOg2MKYSmpuBirXlL1e5o7sXSwR6XQNMZ6EYZMfVqskua8COALkxg7IoD76i
0MB7qT7fBfZKTiLChseF1W4ypG9QcDuChyBNK0IBM3Oy1jfk4ghe9637wPzclBspzYmdS7qO1iaR
r6Niyqk/yT4l9lWjtNg7GuOh4zcgJTzJ2V69kQmzobvTB+n3Iea6LKIOUohs6S35Ew9ZCFWRYeSm
nMZ5+x0ibknBxi8v5osuRcrfM72nDGekAEPRwNGerSNWuyhWVZng84AZNQSm55jGwr5GR2M+8d8E
i9WY5FZwQRxeYRV6fK0oo7ns05psZ4c/5rUb7cx4zYGUxoTJrb5p+DWhjxtoRU8fAQzWOw+zk4fc
+cTiyqe1xuuDk4yJTSFMF/Wi8O/qWxHwV74ZGfm/hIRtPvTi9N5WVvJ/iUyjmfhKJJJY1FHfNeEj
jMRnLbDQ3Qg+PcBduBwgxTNzL+DVlP3AW+FTe2chDGkCR4jroLIslZFpEQTmlVwbNZWNxF6EptfN
Ra9/difgzIpBoBjD62krX2m+LJuycRl6vdcFZTtxWvUI5UDhyIp3BhSWWDSB33kgysX1PY2AMilM
9K/pZa/Dmd5YKKGryv+Q6R26ZJTPf7aihu8QZWJkG/RYKio1fvMuNGfUAcU9kTYUPuEBYNk4AeS7
RGeW6fpTeywI74/7VqfKg2rp0XunfDAIJLcBr9tW1FiBNLQWXwsCMMEpv5hIGfMZd8QsDdkv+ldL
n6myKRx1h2Ol6zcd76BWAjbvfYVIzyLS85YyyHMSK6ceF/q0oPUIVptwZSs2eT089o54eF0/CG4U
pUZJiQlSo1cd6iItov6ZpeT0TItlbEw73K+BhTuSo5TDx1tDWUJmPrqYDE2R285p3jKNT8RWjOQn
PvbaeSNcKF/PESOkOna7fTFWJuyYfpNiERl6scT+g2lx6R2MKuca+mMdOLkM3Uc3BgBhtu9IHCyS
fTPo07F2lS3FvGB3CY5sShkb1HB8c4mWttbMMBg9LJ8U6Buuso7SRduV4EIDmMa7azZLkKbeXdHi
R4/EznyGaG/dReLOVJG2FFj/caGvL08hNe8v25l1TlTeSk2TxA6vpOoXvQrsHSeUK+inj6/N8QiX
2ODDKnoFpdzfEVJ0IAI6kB2scool8l3xDsJ3Jo2d3FY0ECll9EkjrYIDPqjefWFjGhsktpF8vkr1
smXxzGBUuf5gsZ+2vCnK7AoizPqAgB+euFKVDEXmm/6MC4xqp/PFTeS6+UnuGWlsFhCfz0EisYhS
tn4kzhjjT7y78nnOUL/kwAXjmmWAFYZG03YRQQMqSSzsjuD2yLKt31OjgZiTNCfPx1Y2USRg6jN1
sJ/RGgaorRTeehw9yq29JiEaWy9Q9XVq7GGlJQ6ntlnuVFiUbKnM2d7Y6FaSS5rBfTmM9Of/0EmU
rlzKzFRnPC9Hs5CDIMXGyft8O4QFBdMeQko2sAd7izrKyekNrLWGlFwUbRklfECDOJyx0SZp+/At
pvltZ8xnpwRJxuKP6sJ7xQc5ATa6stiUjGvQPct/NQ2jrCxTLWHirZWzxBGu37wWOg6CeD9wiCwr
jP7Nu+s+GLTdzlWVcwTlnHoyyOgsmpGvd/4q6die1WqtJEqtn2IHTQx2xsd47rNysKrdK8KWGAEO
2DNyYyC/jP3eJxghXA1K4sFgkyaVfP/onJGoC0Zpj6dPwnRaEkEz5V2RTEvMN16acsP9aUz82hTM
+U5Zl6FQh7P1gNrMoHIfny2dKqb/B5cEWuDpUI1ZZUFyjDKmx0wfdLt8LwofO1O9j+IZC7dHDzsM
2yE0PAls2aChWRrfgWFU11payuuAWIBpEAIbjaksvs7FnNdXcb+BRzwp/YtQJC2nxUQIkoBwmyAd
bFoM1RitG4x1WlrfUn0J5juz+rMss7Up0Nzv/hHykIkwCyheBCKMA9bHUkXy5fOtdJc0rlDnu3LV
tnCYLZo44Kx32/y9aNeln9H3eQlZyuK93qTfYS0QHLHOBspjXlUNIx6C6Z86iSzunKDYw+VbBuC8
LV1KR8EuGr9AUGmvqIaK0FM46Xb9xbJgsjhKDQusqpZg3viBz5lDIZcq68xhNaSdu5uSjBEE/mkq
M8Bk23y9g3p/3jQQmDKKTFgqc2FxUYobJd6LvnD6QGQLqis7pbZlOmqtOVS7mDeHsTHR/cznRvTb
RcemGt6qyMPUBt3nHyIBxP100IAga7eRQzCB96PSaIyIYhgPx6KqtpsOzeispNyrIju5nuN4oKOG
sclGTZ7nSWo3wG5WLNEpvp0ExpAEpPL66numljZtUuiZpmJkpx3hI4lF6uFZjlGkghwLnqvF3Ph/
+lRh3Dgi8Ngvv2T4hzMStl1KPokjVp6pYgt2wk2w8XAl7W7WbkU0PjkEv+AjHRx9w0kOnwn9x5OS
Q0TpUF6iD6OoKYuuEEFDASOoi5AVq8qShc66EvzlxbuyyKYjm/aRRv96FzfTUPNK23h7JRl0PWTh
jtTcFqlfpJKq1QtpSp3M0QuNDklhqfv9ofHu30BA+PYKeprz0iMj8YmEiNUtsoX9g4Ojdom23HR7
iaNMJqTcetkbQg+DcO0T4DIYrmPX9FNTGS6rVpzoXtRV8tQ7+75vYxgFOjIpK6+xjcXdRm+IYqza
nWfCiYgowfS5fS52FTMEICZZncXf5kaYHIgfZ00UrMhfRENrm6iZ/R6Ovz4m8DqjA2jlDjooOysA
fVk74kcRrXUa3VPstcmeYDMZUVFJoM6Nl8YSWiIpe7RuHUkn+g3+m6S7Ch7K36ePuvlCRlfpayfh
N2eDHRG+JBQRABqcuMCnOuvG3Bb9MKO7SZ4dLTzd4zsk2kJK01EX++rPJCyi50qser+LRbL6///u
ND21nuyEmwnZ0tX5OHfMQHOLFbND8j6utsFkiNNiR0VeQ00XcGRaC7n9R/31+3GM7hgFZkmGE89m
1ayAYjpM+BmLgsiSJgAUyfey6zAEFB/nKX36dDa/0qELyaPMw6k5R8eIKafOjXrBNmdjVYGDfdRy
1zT/YhMK5n2Teta+4mwSCGjcj205rJrPXRVP71AbL/1QppcvXt3GqbU6khGnBEDlwV8ZrYGmfvVM
ujRapEZ5vQUIwvaTnb6OKEHwJMzmUrjMcFOTpRSrmWD8uTVICK9i1Ai+3EqzkcHg7OmP77DjhMqo
G9cGZKDN1C8JpfHsvoSpzgWTmvtGNu288AsruP30WwO8hQNASEyMNK4x9pEJGuNNVc0AhqmxNaPT
COnGS61DPyb3J01ZNf3CULGOeTTef8Lkl4MYzcsrIVvhzaLrGZT5s2JJwhJB4SRI9gkDd+F/4ykJ
h8UgpbezaipGAIo/vfhOR0MVpXDQ6EkSdzbuP8yHpo9dRj7vGE/QtQVh5I1yrGlRK420lLKx4L6u
zzRcOWIoNym53i0u1TyVNBMx+0v4VCqPNhCXfOP7vZE9IfZeJgqH/HFn0SVQP6KzHzeacgYCZ8Ah
Bv/zT30bUP9yVR+gtFIZahlwOoTk1v7X2LSVhl2MNCffC29aSYyuVcEKxJu6S41X2vuGVVkvTyl6
I2KWEdxF3Cu/1K/45PWvM6SWIsGVcGfIZ5KeLk+PPKQbei0kADzkmc07ZbhxYft34GDRZX5ygyzn
veg7Tp6qA2iZD3DeEU00xigQc1M/6PCwO94kjF2iySzgRLUGu2YAzgL9GQji6Gng4SP+QG5cZzFV
iAxJIxjk7bSV/SQyX+ZHLHeAdc7sfdlD+eYs0W5+O8KRSAeyrEd0RmHEoRl0iQnuwb0xwqMRt/EL
SgeZ7FRnE9+VOLTNmPoPjCxY/ljawvMRQLX+cQkyfAaLiAe3eAdgOnzmRPUhcUYmQiKGZ/cmmqJ5
TVUS06rt7nJfdrfV451hfnyB5OQn/esSXXbNajg0ci3iUtc9ZnXkN17MZU9UN5oiUIORKEQMru5u
nIgIAZro15f89qM31Y8F9wJGoaA3CDfXBbzONmd6z134E4DWMmwY/mBuFFzRnNq5ZaJVI04z6xG2
+kkGluETg6ydNwavcGFfPJ3mGwg8YfQBYr0clVWK9bIYyLgVyTTHtH+Cdp0dWbyo0up/GaJaw6HZ
EwO88Fxgxnyie//FgHv3gUCtlmTcHO/HtxkyPUYltqkuPh75XQI9WdlvkaizZW2UEWQbi/CEmWhT
fS84oBUJHJH96OO5jHaWsmQiS8ATVgBMn0OcHF0Eg2f05+vhNpzIW8I7LlJTxtx+n1IqDBF2AExO
ibJJH5ppPpgqlyuzWbXn5wvXXWf5VPNVv69l7cbSE3wFjEWaWWsUAg0eaNlV5HtsWHT0QcKgFAj7
wS/TNfh62OMQdtNotHBYqs9vMBPutCy4En/qWXBInXsFQv04Ebgsu2t6aorjNdm+xYDPljACc+Mv
UoqK1Hszq1U1ZZpKM7+EPWvLKoTzSrNQgDi18BFGTOZcEIl87yY+g9IcMA4FuyZ+aifvOXz+kTxa
pgI4RYqJWRUhlh4XLUmdPX7vyDDW/w3MisZhefmVQlpcI5G2UjBTGoOD7tB3nLR42Tk0X9DMWzuv
66F7qlNFulYlbXZPzn7k8HGE/MxMHpWKFkUIrPFfQrSpmaUUfFyo4GhSEUTEuj75J171iKLgBxab
/kR+NFI8+Qnyl+iKPC1sfPZJeiU1Wnb1V/dAntL1rZsF7FH3e1T21CZTX3i2Jg9OcGFe9BFpuOM/
EjazIk9RuB98VG6xXnNiaJFji94+x344BcKbR9h/R+j5D7zChBi/QAMqxs9Dl4pbRYoyymvcEZ++
mGv3cXoWtJ27EcRRHwjgDmsS/t+4rQx3kJ1/YR8op/4KBgO1daCd1vuVn9vpREPkERoSK0PPzAKO
vuBrNPjU/OcS8xudTHK52Pi2uQO91bIkuyEWhO4q6yiV7LUDo0AjxbrsxEinNAaLrHCrNokawejQ
pUT7ipTkVjDPKmlfK06ETTJsGBhXVZPiPoQMfTn+ShPN7cP0RS52x6s0YktH0YxisfNZgkPhZSwt
H3sPj1OvbMUzHAE6C38H7FatN0oIcUfXhWLoooHSIbdQ3lWbGFwMw0EVZuVZDnZ7KNSpjJNJqcZ2
/IXYPY3VOFD3mwGGT5EhR7XjzxccIFJrE28FY501j+JxaG9PQ3oxi4o+HCYoIcou8Z2u0bhtlukO
mhBNvsSA0Ftj7KJefsunke9e/bSsByPfnlXLyROEfM1vm1dSSAyldowKfTJDpDDfQC6gr7IwOpak
+4sThGPfu13xuubyJGEvpi/SOleERka5knWLDY+1Xn0+7kX4w72zybP+78OosGaYZve7Gliqx9Ka
L2+p+S8hkHGIEdRdnQrIeyG10nQxyyJYmUuReL/AYJwc6hl7zjkrhgvtJvMi4WLGdwJW9uBLTLJf
+oWYtDNHi+xDmuvcWgpJRZuSuLmoUz9eWG2WlbOtOMxNWYz6yCY66PwsEU7JFRBzRn0EWms4UuZ+
tyAApeSDYkG/OFiV8EsCF5yF+YZb5IHSdnKf6Ph7kQZYhN7pvH+EgU0vKG+0GDql9NmhkEoFgFbg
lyyO1XflmwVvHuHV5rW6Si/C0JQZPqSbNzkf0kCPWb7hu4XY6xEerXW6Twfah55tGntSz8npqzcS
oDiRlT3FyLwYBMAdb5TNRXh04dd6IPjfpU8+7RRb/Rlkbpa+eeJt5XsBxRmyW6xmN5C08lqUBL6R
DRoJfvyHsyYEZQ0lKjpQsF/mMJ5KDcDFk1KauAtm4TUGu/AvejSFveeNZvKHuLgq63/0t6WdplyL
j8r6wud+ILIIHwmkFz6kV5MnKhFxpNXbrmKmFk4ezMTnSQ5yzZXzUF1AYSylkxWqmSTE+bSz0wLj
ZHdUTAns8Zdehv/GvrgmQb8BBg9LcWKjvJoVOFUqwLnz42/8kcK2tvjdPVkZj2Co8to2V06PREZP
WC2WlRDvn77LtCEsd//QF5OAAYU3o65c8wgFnxs+4VTJEQdI5tTMQah/oJZjWMPWf7PDjiiEUn46
O25A6h89ns/Kh9R4AeXIih8sDYaaYghQki0xltRHpvShps88Fg+rfU5+tHCtnU18oTqqJxlcNbYI
TOy8Y9f8QTSSWnBkXiANcNcU7SmHzqtc1kZts9jTXw0t0sUDaFz0mI2FNudVt8NV9SEB5KTPlWUy
jiLst93Mp0L3x8ER/+t+OtBaVLZWPyw7lj7QvdigrL4fjH36CVl76nf0ciZPB/vZQYaLvz1vwiE1
kPoAfJzWfotGvmGGZigfOWiEqj1AC7vN4Iiw9P0hnbkpM8J9GzpyO9al9zziAO3D258sBRkSs6S0
YU6GD0BaHX17jEf5XIN8tVbVt+Iua2Um5qo7qCk40nWROZMiopgVV4ire1sQXDaMX9w/ObXgSVIU
f5zCAfcWlrYQffYij4VRAAIi32U5mwr+RClvZEq+w6C9m2ROTeB3NBaZKmiZBD+b2dkdD9BIqOTb
F7PQCssxQRKuPJG/CFa/OuxQODRCkFRrNrtF8jswjYL3xJ3242/fLpb9Sc/x6hLzOAPhZ0uqWDnm
AYxBi/DNYcX9SeGUQxiNMfUNDC9qek+LoH+7+A1PBAgbhGC6M0hy7LfeWJ5zi9a/u5Zs/W4JcnuA
5xWMN26ca4LLlEaIyQpfs7DGewEbylZ9oHMTnGR+97FoHsns8/cOraSGonBC0T7dtj2FyiGg+eI/
/rSSW0UxR3LRIk0TaWCnBXjbF9SjU6tz0MejdPsEAKtCfyjYZ4jHqUA9cayjjPrKcApRkaEgIlzp
WT2J4Czd6d27MyGRzmRD70mKM7PkFdyQJU73SsvPXN6oMuZn8ZWnjMCObDceBR+VOoRwmLEUCWNy
9NwqAWCpBBqWvYGGyIS5bxqzn4mCqZPeANySk61TTa1RWPhAeA==
`protect end_protected

