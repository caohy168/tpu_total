

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kPMKaDOi2kQXuMCKSdPBKatSDEqsZbq8dJQr4x1jAazoyE/zREc1R5J/FG8XDiEZQa8nw9j1ix5C
oQvQGXZKrg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qLeApUbY8ZXxl+1uDLQ1NsEgbqOrFXLgNDRZCtdy+tuQcsXM0AJiWUKY75eR+midgoNqD6w7EInO
ie3/tp8VrUrbZ004xy4XoAS9xgxtpDK7zidDI9umrl7fJtjyo9eyTv2JnFiF3g+9pTZrylMG9cyL
Jqdjnq4+UcuchR7QuMU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xnQyIQHzqLl8QgvKsIJHNSu65sa3bd65FP8/+jBDrvhjpx3AFd+fwTGyhqEGg0LLO02WqW6Apap4
SZrmb9BVlAXKAX2FpWv8ZQS2DyptBZUqKJelwSN1W0GK4SL3Aypfzg2EBF5/q/OFQ6+flxptDiNG
EnKZiLXMdX/1J4Tj+1tjCxDXDYaw07o/YKctzqbqesbUOb1O9e5Pzhq+fA4LTgW/YQfuObYcctm3
liRmYnsg0glfs40T1YlZuMnsG3VLcf6TA8Qd5w9qhSCFabAAalfNy1QkOkm6l1gqJnS7k4Du1tkw
MlgEyUV09+sefXYVTQAkq54DH5v2E4QzMjJFjw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
USCdJYK3gibHILCG3SZ3rb4rlPe1EhirdeqNsVg9b6Mgq3qJKWqbBaAuKwIjo+Tn4o1pD2pgrckC
cOQ5ofiFQuZJojzr4wwMCwaBuvhfgI/ph4zv8ccFi5qVRkYlJ3TIQmkJumbPP2t+QDoJJvghELjB
psgLGLrk1uXjPvrZ+AwGtIKiK3PQ+76zch26VX2KNbVfzFf+zQYvdp5Ucf0updVTApLbEt61HHIS
IEPPXDO5Oi73S0kZCDAXxHz4AGX/EQlNMwb+ddqAkYTcqY9FaWy3GrnMD3fuB8LtD3O9he0eZtEy
n+YGhLUj+NxpBXpKOMPjHH2MeRRn+cJVH4/Qzw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fw2Ueu/tNez3Yov9HXY5IljhQKemjDQX3jbPt9ijSgyTaMBDw5Kw9OGOvX/39JbYv7R2dcGbAP1P
/kWEmSQMBA89GmYeaTGGt+Y83GnY/mt6zlTgS8D/ZCCbHHXw+qlNNrVhfSARjlSKhj6VppGZWZl0
Z/9z38jibEwD7vn6lrW+ir//DI6BfUjYTBLXmYfppC3D2/3udy24bIFP0hfmY9zgR3bc2D1Rl5r/
6waaZQkK4WwH5lKNGqHdDOUvySiNCfY2eI6+parBeBu09U84j3/aBmgL4A31Hh+KVxmFG2CmPiSo
lrYFDLXO73zRYbDZ8IBU+S8cPzXrNNuT1Th2xg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b2uOQkA0sbcvZoGixYW/raDVvukcDKw22dxp5j7Mw3my0is9Uc9JMBTxHWTVCo54sL9pMpsNrr+1
9P2QNefar7dewJDfc6VsUYsuwZvpLkPtPyKJdFmhbq0tfQ2vaHAr51xPIRE8hjeIhAqGu+hpa34T
PFAblWc4afnyp+kRycw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nRBwi3FFmJ/6tXhRn1YPnZ+j7GNxvO548dGI8tBZq7sGV2oYbdspjCmXgEAGFMB6Gn7qV66rW8HW
i+8pOmwhY0+xr14RuwYVh1ued31kJp71+NEFBpoQTta7c+m1PwuinGxE1dVA30y6W5BpysFvceHu
kjixM0ey4iqe65QrViOc3aFMoQkyNG1jDnNPVU++7Gz4W2wPb/sQxTeN2+p9uYz/OZtk3mEbAXeT
wLx8I93uc83hkZCsbBWkiLx5skHPnhGWD3izNSDLaScE+bSw8hwv91RMtLF/x/xcSN5xZmWuZvHg
m5Lvl+vMZFztzpt6D06wDkAlLioGDe9TeEzkiA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SvCVHEI+mCgtjsQ6p8gRD5V9avjftzeQS4O0q+g/VoNHuvya7RUs9btiXNIkrRJFV5Aj1b2G4lYB
F8F4jkkU3JCdC9kJt5bAYq61b/I1sy47P+BrX4VfWtcwv0ZU1u+hliYNLweMc4nBjnMLai9JMFHi
tq1VxNnMGx3tC82dfRlYCXwZt9H9Gzr4QFVY0NH6dgHUeIr09XKALiJq2xoTckJ4cEosT4gQrjwh
JzehJm3/WLtM+ga7ihKtNttmvr4EuWqJV5Ts3CwI8No1ulolCG0+PaZjXyXaAPYs6b6+HJS8xB/B
JnUQ/C6VU4hJXwTNp30KrUn5Zx3ag5/n/nKodw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121872)
`protect data_block
0+P8s6ygqpUp3gv3VKJ0nnHNHDkqCgjBiVyoEyzSwbf5+rOAuMAA/b9Fh+xBNA0IRFEkQP3musei
UVJPMFnyBG5iTYH0ZLo9wQSDmuMxnBAfCEt6t5jKJRxZKh45CrfkOw56PTqW9RdyywjKJp0zE0Xb
CuixKaQdORxG+AvaasceI1Z9iurjKA+9SSosoQcf3DVYRgRyyvL4mme20zBbyuTrigNae/MZHhhS
AOAxk7ekISv820Oipu8oe/Eq0vzBre6+9jUESGka0Gc/zKJVSJqERxG5lT9Z8z0CbFlbldtTHWrX
QcY6PdTVuhYAIpstAYj63jrkuguurYi8KrvLd+wdUqJcFV2QSfztE6jwQIe1CVu91Z9LgthXyj9w
Yzh+ooJ0axdFerOixXF1RLhX/5zCw8H0TYhMr0QLpd95UiSX5pyVoi8nsKWd+Ma2sgD7X1SKVjBi
NkElmiJ5MBEBkYqtdPPHqc/iAHNAsUc/F4DGs5dLsSLIIEr5F6xWbQEaFuHXLUEIdUPSZHADPrY3
I1EOsWWNcCxKMmpLFIFOdW3JXNDe1xWbaZzK6ESW5CEuy0pBA7f7cz7srqonnJOYpqrY8F4bGUJy
Mz2gQCWFduYMyhnI2LY3p3RnRZ6aH0H4ryxhZ26s9A/cDw6JNPxcj8/wfQ75fmmBl1o94h7pD0TP
oI+qSnewpOc7YzOumezTsdDKTnVvjO7gc/INzmQMnp92OheDAsYT8ckFfjn/IhO5cdcMokNF4iMO
09qhGdl5oDDxMKWs0YjeyFnXIdIe3ZKRP3eGN3ns/ZVU9LkSd2huzXNTEseeJIcPfmOm5JUNnsxV
CkokKddcyF0xf3/BVO61feC2ux92UxYP4Mz2nZ2knVoDpzrUekS3DGv0QG9OLblc78Z8/1rm/smY
wVDiW8nTyCbkIY7DAYa7i+ol7oCSncqViNVn6SL07QmpHAaCPPvYB9aK0bKr5EmRaMJIwgUV+OKU
i0cuPOtA2RsiMR8/AC+fn4Xq8FhK6A7bLAB2uF5r39jvFPvQN6DrrQkjM3Rf638K4lFaBwJ93BUf
IWcCPc27EX3IgdCS6hV9wrHJYsv4pMwIiV6tYnPCzWDzf+6VU0sEK7bv7Sa+IvblyQb4zuaJdA0j
As6BkkmAp8NyMDleGDd6QhtKNlcE7T7P/NcSkVURiGdjg+f904jfcC5r9dXlfX6KbMN8hCGizx3O
3SuQrQ57wKHdmhbRmZSpRy2vXUSFB4KIIEmEHb+jJ8iqUHzn7zQby9oECJOb35bI7Jq4Tbby4tdH
cHTfXTn6rSYPQTSQL6R8hEXqGJfomFIPd0hf1a4jFmKvSKG6/Wgca7TPaAjSHeqCj0+et1jMpMN9
/HWaKW6O/wf33Ij5HPgj1PVTElrSDqgOZ8LG4e4e02iKDgzPXS9j09RYupMplEMq9LQd/m0j8yyK
MzH8ZYOMEPbCWCVt8o+U7KRit0Azbn/jzxJX08Xmmve1fv1BUlkj7CDn5WvL3eHpTV9aDQoEnNka
TrDfU7LY8QJGtaKhdIk9QnlzE4w49jjfJX5wfTAVFDBgGg/n6pagZjCaOQZYToxdQswA4JLEd8YU
4v2xSs1+7Wi1BiT/ODkRoMh8YK+mUDQNi9mcnDjp1hHWdMWavfyP1fV7cLtlAQvZQJYYDeeio/3F
iBUL+n4kDe15f84JtGL5ODfu92hkwvJuntdJO7RXwzt5+jej8BxBNV1PifwVY/X5moN80VMURHvo
WC4jJJg6Tg9foakYwHEPjm28bgc4xqVHO2MJLbHK+BseCQLfCcqm0V5Pc25jLPiNP1We88IdGLrB
6qL4pYHQ2ry4EHC3S9WP8X0QMW0pHE5CPgOad9BCYjxuQ5duAitPKNa1HvZdVVltQyY92kBHgJOm
my60fGuDwBpn8J2/uu9w4O46TNn9YIde3Tci6jqYy56yP94FBVdDqmhKyl3sSkBSFa9sId4vE6gf
XWkseJ41EXJLpygg3LIv/okyhtrQ7ZVitJcyhHcrM3vvwj2lo8F2suSKShkP9mUUm/4sn23jbLDl
5fWGSqfVK8iEIi2Eg+qBQ5AYhHEmq4AixBCF0Ux81NZrz+ag31tMkTYCh/YbJhJiycHSkXmx2tGP
B9fQ+uH5hI0BEr3K/YNQqYVQjlT1kntQlivV+TyjvQHLLmV/14tu+R4o9cwSKIIKwtz0DA5y5KUQ
1uh838apSU6L/xorRiA4mSgAZl7lrIaRGqbwrByzrtShiuqBdnSJyhHWr8fs2T2n0JzBE3vy2OsV
dZ+E9VwdhkCm2gXM3EojLOdUAxz3qIBNPrvbG2ac3wYW2zjZAoxT5iB/Ke2RSNxxliKGYSZkSgrF
gzQk5AtxD4/sVXvkNmFhbzNkro1XGee51o6aYrbq3ud8Ptz276m0fPlnduazYcVJaF2GMXZCIcKB
E+FXIYKxF9STx+urAuZi6HrWwbe6V2NS8xezQ1JL/SimZr8fAFNPInyizzPmVKVfEWbPJRA7oyNw
k6ug734PKS4cyOjTkOgHkJYndFCbONPUXefVXguiPo0W9+cYIOnLq5bwAeKiR4aW1xYHyCwDrsD6
m8nEgS3465xuKuZI2AOgiioa3Q7LiOLaDbXkrlYjpAJwfXraPHMRErJlRPiqCJ5LfUsvzBVfTmhb
e5qLTIqMJHJiptiHH1ALj+10cJFovctNHmH04fGb0Qb4uURqf7nyj91G11+elgLsxZP4eY2kQZA+
m4tyMyqBG8cpD8kvowvAAsVG42yODiTZvw+IFuB3VJY9c1IXL4DnUetr8qYIlTjN4xrrm9XtZQHr
tNz3QlPo8QBEQ+mnXtDhgyc2QHDxEzvCP70NmiRDXboHCTWiDBeFaZV79yrVAQUal7Td0R0D7/qN
8MxPT6Pu8EShgWnkAXiwQCF09pvXmqbtfm4JsNwzRiw1oQB1jAbwffNq/grECglZGI5I+cXXGBEW
YQQ6xqhePsZUMFY8NQQTQJm0s9K9XKaCV0tVLhNAbWecc6+s4l8YHR9G8IQ6qWtff1VsXB5IMlOA
9fcOgBfQr3XsCcEHZzyXDgt5NIVISKUYDztzxnKxsoDXDRk+NnCZXW/fC0CK0VxoRVGy2xGMqQLP
+2fJkxvt/Am7x7K7iGt3yeAtwveyHYSizA/n8Ju9kxoOwXMBty1RBNcYu299vXJ1NhHHd+ADYdP9
y5LrD6IKdZLhQGrdSsH1MsZLsfcjx+BITJwXezhPuNArx4JETDTNPcKply4imSNEJ8uDKIxzS1zG
sQqyWKuJEHnhZQg+2SgBnfjFGgpdfpkZEHNmKfcBtfvbSEBrwh377DkKIJFKgXxphUr+OO5IhaIp
MHUcNnDqMgQCK2ZlEOvhE5H0DAil+a04jJFdrtOmhz4zzZB+QtDn0FHzIoWLc8e0mh6I0ODViWam
XZcvrNQzScqepC06/k91w3IGeqPJUS9maoJwOu7/FJz8gt84FhW6JJGYS+E2ISzTHugLh/8FH3Yo
HOi+yJWOPtJzbCx/BtLden/zxasiERs3yXf5sUDCDGNFbb9kFbQbawVN8FLVT+PV4hmlxRhsazGh
6It0b7bbBjYbAMmjk0krvfDy/eAl7QCNjE+nmO+0xX9kdsFXXuuDDSh467Fx7mIHhDtfzGN3pgtU
IrA4stxikq4dF9YsNaCRO6Yo/s2nDKroGDF5tEdOhXNF9orV6Z9rD3atGns2Qhci/2p/0mdjeJ8D
7Hz1GD9+yuiLlFFD6stvyYYdCUzJrNlPcPd7Rc/H+/wHqZ2inZYp7YQRQ5U6gcMIwgGphSQ/JLZJ
KaBN6owxMSN3g4opVElOug7fveU59jOgDELEfKZlaLxHCid7O1RkXIx5FTjWMRVNZMPP3anelsSz
Pprr4uRwtDLVGNU9PtkkM5Zx1DNt0HHeG8U6nFA4/imyViWz/4u5h8zyWEC9kGw2P6ixAUdd175r
Yx5Os9Hq/Mg+jJMtE/pHIZasaxAd9l3Vh4teS5Iah6BtjEPZ4Duvhml6N5vwLIS8T4d8o9w0E7oP
YTunQlYNEdUTcf/Csl/dL1nvk4gBvQw+4tC9leGEPTB5F/K9bLzJpdyJVY3TYFcyX2+6V4E+4DMo
5ozV0W3Y8Qhxk5U1u/Pan2sTJe/w57L5C1dF2KUqDuaiOwJfA1hO63Yp2PGJnHScKTerprnxeNs0
mx58lCIYo6h+DnCWVQmrYPlnwYOoDe+VqYXusTmUmpJTnhDlLKYYTgPpqVTscJSowR7TvE3APvOc
JdSnMLy83mbD0iJ4pYccCIpAW6iY0Xl+p5js/I3dukJY84wMSKaunZTafKR0sZ/B35/e/sYYCULi
XwVrwCbaCziEBT69I6Ifvo87auD8FobPzs8YldE3OiSswYUX4h+FAJku/VhXyqBh+6xK43C6EMq9
wIRprEIQbtU1yynLGslwDSsY3elBAphYC38YN9AXNlGG5N0b7vH7E6HOoF2Z1FLW/AQYpk9RoBgw
9QKbAI0HsixCDhts8K9qrl8+3bK+hwquP7uyLvjFfIkODfYYHAEmDBj+eqZGHtqb5uCPHdWUQBxu
fBqAa2FjVnooFyhgBDyxu6BzQkX/YMuFHYF2yNkesDKGA9PNrFUIbn4lWM9pFJ4c20lmGH3MvCz0
9HOmN4JmpRP5aSl9nJioy3mpD7UsocAoTZcYiy8piVP8GzzvT6IOUDfECXSldqEAflKwSThfnoez
FtanXWi8npcvp73z+xve6ZhGx5wtZqUwx/3tY+OR0KdQTLzLi28BKly7hoNSDD5aKe9Mym4Q9WBe
LPC/ENA9+WPs0C/g3UxMn8Z2xChyvqo/SFSgK4zWOIexEYIWfYAtBsnflmFFGAnMqxUzDy2M5sED
3g/8fPeWDdzrGRYnyWi2V+SWue+8RrambWiutlA1CpK0FsM0p8wVcTAQpcS2Azp1VfU9nSSAuqxY
2Kb6omIMQGbKJYgLhttBdaQ4YoxikyjEGfw81pNOIZ4AXymfUYUUV9M0QY66AUKfKfnRmePtg+mr
STOiwtHAxJVXyDCSvkcBEb9IfD9hF4hqIsAE8Yp17hZtKs9lWszgNp0G8L6Q/qxvDqGVERp6FT/w
Q1HytFqsWC6M2OFO7F8KBcIe3gTK+7ObjyCGH8syPJXUOlBDl+uvgtaC1z0qYqa0VJdKyrhbBkJC
GYPGghHPP65f1cEuO18Orl6D+TRSmMwK94DXU5oSLMmjR2IaPRDwCKJlAb9QKhCmnrMrzlTlTLHz
unk+zFgzzOOLwOc+pWQ/hw3Zouue9lGRAF4RMRLXJhBXkPWfF82OExfn0KsVmpwT4oCxnAZGGuhb
P/VXaSNTRcK1yI8O4UOcamzS5sbBH7Bmz43cD8+qFcyJWZN0rvKHhEMC6Zk+KYZBFeQ99uiOCq93
3+ukP4xKDXQZdXK85NW0CkI59h7VLI9QFyOMbnI2Ze9MW7JNXYNlq/5l7HAa157DzCtLWCu/L7La
oxhFzXRclUQ0OrmgfaDL4rORmEk9zFksNay4/T2puJPa/KPSkERHuwF8J191/+pa0OFMPCaKRnmI
G/ea5/hMMpyli6FYDbol+8ZnYVV7APojb9oTmGsCCOFzVYV4bTy+hLpgdj0ZKQ1DlfSZbqzd+q5u
76YY8uqwP8mSoARj1VbUDOrkVvEjO5YR1w+RLu8gqfehnRtIDg+1359GHNwNtHLt/JJCNmIFlCi6
hOuyiq3VIlJl5TQ9M6Z4Sp/UAvJu6W03u8vfpymoXzZDCa6+i1enye66ybbRpFrbdneArK+DiqjU
fSNPbPe6GTxYm1cQJ8AgkklzAAoIpDUt5NkCnYBfyR6u1cWLXyB5b4r+MODUL7tsuO8K5UzwOrBE
8wfczavSXsI8wGcuYgvB50ZJ9M8ptRWo8ESOesUCduef+C25ZrfJhg9kJxB4hvbU13JelPX6yEmW
krcRdqcVvsl0bAwdrNDnHRu1NN4HlcJ5IqXwJmsEQEC1FffrEnQ0hKLdJgzzYRwTYrHEmZg7EM7t
kTq6oD1ZYIhGRHLMsuKYgJW40QiV4Ne+5hqBVArUljNcxXqgkP3Q0VMBZV2zGyIzlfZ4j3j3FYGg
UYgwYIUPDpLNA9sbc3CDrvSBa7bcVeU5Jii7Vie37yrhhYbOrLpTH8s0GepIEOeDqmOF7tUfuzyX
+WT+phbjuXQItihTNhxVQcxY3JtvJq9Hdpk9NNhb2lPMm1nUnfIciJummBpYftN2EeCnDUm/EbqQ
/6aDTpN4pTzSlFSBz7r4A8/s2zHJq3Yz1AV1CdmCQ8pamD7um65k0hnzF8wj2XSV4Xh+Kp3fzHyD
0O4TPHnrI5DzSpIRyCbh+wJXAzmHrzoDthbOY9Q3+a1nY0xb0tmXBgakE1LXBVhZm9YQOidzOuFn
EY3Wao5aySI9+TmUawK33XmG47HGL2v7kgn/990qCvadlBeMJ+A4tWnLLlj0vaBZ2aWRCn/Fm5g1
nlm15wXEFkmDHnZGcZM2bZVO/40iGr4mxh+Jst0NX0l1Eb0WbX1bUQjLLQuzJlOZhwBU9tuNBi+7
UTim60INRCc0tmFMdWuvHPMUZ47ROSF2Xywg9PMfrX9tc26wHyUP6cTUWrFe3C17CGH0TNrIxnLH
4mFEbHJgU1AvEDv+C2GUHOb3OZpI9qTY54QXvuOS3WdARB8Pgr/CNBMMCeF6/GJ9U2z8JtvTIOn5
7pRoGawZs2C8+desmdqkX3b0DAu8pmWIjNnYckSDTpylBdIdi2dUducNx+0hqMk/BLgGgtOuVpk+
JYhBNAf2OMXlpXuGj+iQkl0UN7nGOka8qOVoeT1b2Pl4xVaFrQEaaE+bQhx83T/kUn6omS4WZPOe
wPYG2ESSgCczHQNhcmcyDkQ3Z2eFIhhb6VdYbKDcVMWE2R8glRsCN7gQ23J0iJvR9Pa8z72cS6k0
rh0iAQyrCulopYhb+jpUZUPW8yKQxzgGI3H8JEKrvy4RieDOYIopVySQusiybmTYABXWSR2mt6Nv
RD8ahTm9KsvUy4iLHy7KD1pz3sDq6mhoFsFw+43kTDfpoLy0elwvTeQljtx2skhUafvF8VAfgDYU
5RhZnRKaBGGl5C6bQh5Hc4dd5PCehyUJW0QuPhiZBYzdSo0f6B/gDxMUMYUt5c8ZO4X4KBbiLbCN
+FYUeVCIiGa0rs9vmBo/fFXyE8PznRgfJpP9vooUUqebG9cJiylIm8rpayp17U+3mzqhzpwyBq6T
sVa5GUWK+4DmpgvZzO0Tj5meSW15aeeQltnJkePV9zMZXWBiifjhEQFPR69YtQsnXMoKHeOCdWo5
IdHjSFTJtxBS+PHDhLvPcWbi1eDBz8u4a/79vom5ONAQmMomzZQNUVS+QRoMaDIg7rwwBUi3ibv0
2VOm/xxuHYfA4KHLVfh5rGIKnuqDmW2GK+eJGUgtQCaD7tE7CgYsfUR7D84bPHH/dhXovoIn4b0F
Pm4HSTH0UBbou/wBwcm4AroUaxGvUOX8x3Hz0h484ApUsNrt583L6PaTur5Zd4p3jcU3Pi993Y1x
ZtAYZAQZUYe2dC8rkLXTn+nXRdokZ0rTPIQAXS+65i37dmZ6oBlxDSMZterFWHCr0YNS1ZmkywNh
Cty2DNJqvfde9oZHxQuDn/Nv0yuptM/qIQ4/pbwuQZGsvrB+tzKDHOEwthWDj29rDeLf+zoInFD5
v9I4KuKD7voTOLbBMnvLHzyujqSttrllqqncA+wEE7VOIEXscSNstwVThv4/1lUzcejQKDB4rtIF
45eAMzZF454m0V+ondeVqNSwUoKOJZmf5uynnPWrDC7jA3Naeh7EwhFxOlOLSHjEc5hGm7wojDVe
ZXQvS+cbNSH1M9rH4B7JoSHnSxTP5weGnHMUUYT8C3oVjhRla3rHuZPh0Gc9iUj5Vg/N/sIz/dV6
/LvmiGEezdNjR3gcRqF3IcpUhdkd/zEgQHP92/5e9Qm8Ik3zqGfqMKuEVxg4brVLAC88LWwoVIPp
23U/k3QWO3aDTCZeaxZqpg52tMV4zgwa5O5j73mv/ruFka+9YfIM+bDj98spm+8eSvKGe1YVPG2e
3U7+xEaKv47Wgv81JO54K3efVcQAN01O9Wx2fLwFnD7xwb2EabBJ4LpdzZ7Vo4oKoXEQYnjXR6XU
ZPMchmhKYZI4/n/TiAyr/Ovzt/QXcYEwbILdkeNoYjwWeuu389k41PMj496XG3rkz+Wx9jcp96w/
xViWppnhldM76ZXKr2t7CBN2moo9FqdASThQLip0az1HvC3Qs8yrMsuTk+D7QJb2rMbEhi8SdaVt
AZv+xcT+O+oO300WRbcTjjJm5M5KVL3NbenYegBRF2lE50ORCDSZNzSAAUOR8BkpE4EPprX/9ykh
XAi0u3vuy7wQ4RPjgUH6ZdwfEEDV5WBIoffdAJr0tvxcojUwg6MyIEKY+a7/uWihswvacs+Mq14S
kN+jYydjngvNMfOoF4UFNCtyScNxTq+EBPiOZpHd5lbofMaUATtTn8HIehkur6e91ZnJjs83O3B8
4tTgESsyuIJK64LRBcPCypZx3iKT7sJFbbp42u8SyCZUtQ5cjuwNL9L5o8Vhymg+lzXJFz9WOtme
9Y2A6CBqR0CS/zjzr9xhHqjDkYFNcvbUh593StWYkf18wz8rPWJlzRgjWkL3hOPI94nl8SHdJUcm
hax3axE71D8sp11UuMRB5DgjvL5KsA1OQkoL5XUQeZHFjVQYzs7Qmr8H86uuVlbHvho3YI3FURvt
vPKhASjOSAfN++LaY8yAcSRoJSY3R5xmQwMwJEJRnES7uDzQlEYbMaKAsup4GVAFa2IL7Qbkv3An
rlBfS2N7Mo86gRYWwGfsesUoDJ/jStkhrwMC4QphRBqOHWhuqMiUZaY9Lz2vzjjPz0NTAmbbwRTo
f0n56G9Wge47YlO3yT8umGMF8U4LFgLFtvAVPCzprdnAg5uvRX/RuPDOUuO5oBd5vyE1+BproRe4
XLx5gQD+oJifSerNF7dOf2GpBOOBWommIVOnNLjOHjzFphaYBdygFIrTFib4Qu5c7CEShBhCivEu
FJ3ADOAjCKh9QR85dTJ6Jm7yoLwxmMJLl8Q+50IAAz0gsKbCPmG4u6kdJzfE5PXDi3b31+i8O1rN
nLBqN6qxr4NLVtoeHcKb/Vz8LMaMWiRnMi8PvYmH/nNdwr7Ne+gFYj48jws72HqSYGLMhHdsITXo
GyisGPKY62qJYX7MSxsHjMlZ1iMsSFaKz/H/p3WzR0zYuHeZcj4C2/tZxhZ/k7Jw49TsQ/lQY6gY
F4xVrYWRMX05lOQhd3fvnvQ1s6ugo0WnhvzYywQWgOQXHCXfxTucvCHuRQ7uSTCHId9TmP5Z0plF
V0PkYchDKZ9UY4Ye+kj2EmTS04pqPFJAcsyv1qkdfBcOjrB0Yq0Mrz2aXuH7Wln2DNhHQzVenz+r
hnjfO20bdHBw51SrM9y1zEmbikvNH1GQP9nHJUJW8mw6Mg+cI7Dk/QJN/zMuhOM3Xc59qTXa6h0w
AhTBRC8JdaUm/17chx56YKjsoX/wqJFN/kGA1d1+/OvAUxMFQ3zhtX3aBm008bFpDM3A+SZ+22+c
LZPKhuTH/PQKbncXiE9oRALyc5CyOuuWJCYPp9HVHmscuJzX7PCPsrLQH/+pKIrGx2NsJGGeltfj
T3SxvQnvt52itMQmS1dkOMd/f9WALV0ZfmGtU5a/N/A9j3+vJ21OdcJd7g7kculvihn9YBRlh06j
QcrfJcko1gWaPc0SKqEpBWYRr4vIjF9aiANfdDSI70biHP8gPnGLLLfA/7O+JoBJMvNCNo5w7xUH
ctjzuD4slyJjXZQ2cXxPqEymPvpyMTq+6QjeFKS/K+arZRz85bmpLV+DGRLAc5vTKjxgmOzK1tN+
wpACdmH1U4f/lbOAtphrPGb0eW2anYewKS5KHd+Dj6Z8zxXd0ymGXzRxPSpX7fAzFd7Hd2AtI8r1
afXWsJvTWMiqs2q/JLWucNvFdrOFyIz3XwSDBejYXwZlMNWLFWt9JLncumoVtHj52DkqySXoaXY7
IehTuKyiRxKRAJujOXrgrPn7F/n47wCLRysw1FXM+fRYF1e+bK+6ZgZHhw/h5qHGpDqcDn0hFoCF
FG4pHQVYUkTi+YfD24+dwJCi10LloOXUF6IBCzCaW2u9CtrXUpmhub3PH7d2+FTDc2YhlxZ2sC21
m/50hvKQkirHOc3C7GFCCV90B+i+X6KxrotLrLRP9e+o7Kj/koWDiIuwnx8me3pI9IAruNefkUNi
D14gRgZ6FLeveQnvgx1wVCt0hCkY79J0EFi6txTf9gQs+YYT4UFbSY932gCzCUKGr1RyaO04Ka8c
DTjoYPeZ3VHDaknUVNeTGxSR2fGEWBlWL7QT2k+wZDnN+2c+GScg5+/8UDBgLq9EFWfi3LBQL3JM
oUOFzU43IHtNx5EQjq4nyInN+tqcsp95kcYCDsKxIJ7rrmWWjKsNxkIcTDjLiL047wreJs0oDsfp
DJ0DT+StlHXo4k5SstDMsPi7X6RRVJ1gg7S38+WnPfwCD4zBWFFzk76mtz1JeZNdL7lKFGLuOEnb
a0T337Vz8RM47XM8XDwvr5f7txHYgnD0BI/UDADSeew55+fQl14zLgMHn+KM6r4tZzn3BWUzqNBX
FVr7bvhdhpa+HkgGGQO2V2+B12vbjp3wxq83MtWv4uq2nMIOZNBGZepCL7s9B4f989iNgM3atwEO
QPDEU2e9c2zi0Wfaz5ttdm5I2URziBIaRYNXg1Q4sGpf9iW+0ouku2kiZStCf7HjRPmmhlogF0dP
6ESDtLFPND0Nwup7/XGP0DeGFgCtGy9QeZ7wVd6a9CUTLWvNsi6rivhmTrqzcv7sNJ2SYlPAQ+Tq
dqg1DE0PeET57l7pSHWP6Jcxq7tjw4w+NS5gxvODA6QQ3HqAwIZwyeiIhUSDtQudNSQfNQUyIzEX
Gu2OYMbTgppgKG+SmSPLAjbksoynQLhFqfbGK9MgjNAipvDWQWKt7/P44FTnRLL99a2TVxY8vFV6
7r/cDyKS2tAOwBRzffjxJXbXS/pHRXr0kuRsyFoBbJAKoHZmb8B7i9Ob746cYoO7F/EreBwLsGmY
67NpqtNBMdp6pr/DNCffYOOx/xFbMhXkOtTugr8L93MyEtTsoM4xwfquj2YuSYp6ocWQYqLsBm03
kv+PoiwbH65NNTLxp0Vv63Mo5IHfJbWXzIOINRQnHuTDZVFrToumHoyU51vpPXWPBOEKPbUuIgKZ
oemkUiC142EhR7vtIuKlWbbcE0/yPTRv+i8qubzDh8WAUjO824SCNvhRu1dWKJ76wHo30sjOMChi
FDJJBi7hKSkUbuvg4FCevrzO6TL6JZJVTMafU8+dHwlBf7zEN7Y0hRrURGMeAu21UBH6WNhSgyOI
tUnYgUlnXxt1BIt4gESkwsxsudauAHx1TEo46RjZcG7R56ZcFHo5Y3OL/LAo+2jQw4K1qkOvacDZ
GLmEb/HDAeGB1tQ1eE/BKvjiEdfCG6DVzOJobCNvQ2z5zRjdX10plF8LOk1S36y0/cvbirQPqM5O
kGRzbF3zyEVtJ1Dpg+REzFS4q3YDQ9mv+M941nrn4fcg0GiScn+GMuatWVZC28U19ROqUKmrhnGF
MPlx24qrfuVq4NNUEFXYapSqObzt6hkiv6mAYSN6wAIaXkHPwYaGQ7/OID7+wNzVkKGMy94vVVEs
2BEweH5pizpaWPvxqkhHh+HWKIT4cD311EE9pcjcSc1LlXk3k2r0QwNwaLjDlxCfQ2cUeGJpKP+H
TnInACye8YlmdzAJjsEyTU6ANlUKUaIwuV58tjc9koDMnv7DwdiJDX/utF3Dq3YFrhchqP3SC4LY
OVuxSaG12d5uDxSZfWRyIQZwA1rRm+1446eEVIggWIHH8iQyPc0lZzS2NzP6PV8OENF4F0C9t8pe
GgBKMKZriYb00DK8pB4EgtaNs4klbQYgrE8S3uX6+8by6wSMhA7k2ihOf+bK1AtU6xTuEdGP5DqK
lGVGKjY3PWtcjePfxyukv3Gp2WNfQewWcv1pZfNYkHiB6GzP1pxtJqISeDq6rLxqA7XnwiAST5W8
eIML+Ae15Ev9vYmIfOYygWqUt98+cN1U5VasUg3BBwX3rnbGfJ/HelkmBP3Q9hTolLAsPPex7WuC
wrf5TplQyaXuhF39Ay31sYINQ3q4vsxOdia7Ac4qE9Ycwhd1stVll20adQn9wulEs9llhDxsG3j2
V85kSq1HjRENIlPLa2870yDVQA0LqQOtyQqrDkSuGNg1IjIv2XEwUsJc5Jd0We/sBV+GSxHg1iQn
ufpG7kvgfgb88Waq9jRSlB+fG8xXTKe2nfTQmC1HAztURmwmA6V1Yiw0Y8NHWxYPHUvsgJSLr13R
WsbAbUzhWdMifiZv+Sq8ltkKYtWS/RbTiQ+egVigKfw+R6FoEq7dh9FgeVmdoJxSAHq/7mGVSBsV
PD+/dn8+v75A+4hdDWd0oxodYWyx8bNIjFd6U3ur8YkQgQnbAGOsKCTFJAETHgXY+KZBavqo7AQU
7pn6b6NHnEm4Uq2eiRO4S1hKGmVFCrZs+0rpRMTE8ZCuIdZlrcpBFP6KQpgf6MvUDHcOAqXd91f4
HaKYt7SPxMTWWG19wrutZv+F4c2XRRk7VNDjMScv0PWpH8dtwn7BaAcnnoy7ZJv6BdVUM4rTQh8h
NWa2h/ADD20R7e1zKvCE2fY7+dASLF5BsGQ6YH4LgteZgu9PLs36RSXIQrOsLDLdeR7dFUnebaAm
7LWqSwd7tVWeFAhB4ZHCvI4OXicVrxCo/yAkmds4KMH/WTPKmd93tk2aCBI26jZOils2m9ilZAZh
19S+WACzLRhU7RezkAKd8P57w8TZVXhZwTiS+6jyYtMdhY3PooRo3Ith+t/YIiukGhlmJffAiMWT
oRGwk8PFwTUGICsiKNq1Yseiw6Xblu6I6sq+xHDJ42AlsXiSJZ1jA5slMAVXhZv4ozcqY7iMmE9u
BUXLvcd9w2fMeqe80mvz8NweQl/pkSmdHHSQrmfKX7A6f1X7dYb/BKWJEXdSUEm4H0K5tkj7rZZg
Q9/XJNEN02gFtG88EimIk+f33Mp2KAqI1hlUZ2QluZgSjv61rL7/8JHBTHt/6JG36WOyp6WzkIIA
IlcFjLHPhvw6iUIzBMMqFZ+BLJrdE1uh5aK1GQVwywtR70GSOrXpKN/qkC/+7MpQTfp0dsAu2iw6
q7+nE8oGdn5PtlnS3SGy3kUixPjQUwkKYGY7c7q9Fkk383LRDEBw0ns8sjbarkLRmvVA3IIseic8
oSBdEALavAun+YRiSE6Vn4XuZUgM0buO8plLrHp5WrNFKcSin0HOnltpRTsJaVyfmRkGPmqwHaK6
XLHchzWVfLjbnE1diWLF6NdbV6jRMyR2Cwzc9XpZXbG6EgGmRs7wSZQ1Q+ZS2cNc9tjjSLYCl0FD
OKfU6ODrXK4vCq90c4RnoOLgpOtfk5xYnu7v0VwpQjzQxxslbnjH1DgM/rlahEwtt7SGbImGsq9C
+CwQNd3I011SZ+X3cdw2Cv4AkpS6RN6BT9rp50zmMwhWCUsfj7w9s7bfnufBJTO8WHycGOnJdtjg
9enMx+vF7V7M84/Otbsdb7zOkW1WQmv/mwHykfrhtD/sBd7HfF806jNGRpc6npv2h5hPHsT+nV5P
n5pUUU29L9/vEYWTnY4zQGNgUSsWvqBIpYJ3KGipfzErmAtQVGDUsW6yJzoaq2tsDNui6otx99XU
7GckbSLM3sXACn63q1o+WNk5zwI1IRfl67Ff+I0PQTR+jidjzRtxZISJgzq8XmBsCx5Y7klklGri
Y3vZtMobbd4K/+qE5WnXRiVhv6ZBKeGDXDt9GFWBJ0KxIGKR1X7sxkPvl5SUkX8pLF6Thu7q/OKh
KU6MgZMGKosy8u1rfuSspgxUCQG3q8fKOhn433gVvsFQCsJGKN/u53tIwdB+Nyr3veQqeRA4tkjh
VbEIyturk6Xey7ooLOUEnQ8m7qzISxZkRn/pQbJNF8xRFR7Jtv6WIFPWGdzlhgnGg22MeCZrjXgx
hDZ3qoZoeWFMqEiLuQixnbwLQrW3olmqI+LOMkSxW+F53iOK5rb/TvdBvzF4JvXvtT6fbIQAAcV3
0OmLwWEe60DrBlOKAhqQo2wXRQbpaAgqkLF7hEB6eITjDBbg/OrLXRmFIVz6Kd9saihSRux1GTlc
aMgg07PzRFuj1DllZuwyRwwrW/NcG2C2VXUd6I0t220NX7r3TySdxya6VmmvJNl1I1sdDOK/KgBb
NNvFGncGzVzeteWde24MxJ9jujYARe7Bs+RTBE1JvxicV30mq0HmgvRIzdkwgsQ4BulrdmALRH/V
IIldbio2MQwAfdJ8tzgbTHUvEvPBk/f/8nf8KghVa5xRSpywHzD6BccCgajn8da2iY4yUDV7ilcr
Vsiw8SQYmr9DX+4tXYek616igrfGZvRvzt8ua7mtv3+lhHfCtjUffQwE4pLCyuvyJi5cD3mIAoXU
wh7Qw7qEh1NuhzYkogUEIAtq650+X/gha8rRq9pR1gt2O4KFJ8jS9RO8qWQUN2bgUO47Xa+uVntt
UIdPJKjgDZOk+K2L3IZuVgEYVg9PxdMT30x2opjbpL8iowNENISfZLUQB5X2ohplqvUphJG6ckU2
czt198skElv8g2YHQT3MxpDrO3xGabC/z6W158uR+1M7HPDJJsAN6m2Gt/zcLgCA33WEgIDR9LuE
LkbrgUpoDAFvd169lBnNsspQTPp+49PMMfxQ8Knhx44XO9Gidcmmb/drLhDV1J0dAU7CDTIoXNSN
6tTLJSiQ2V9Z0utD5T1RcAjECEWjqMdswY2csej6QcxSxwhhNO2DnFq6IKqT+yeRqM3zOwg/zKai
94/H31lf3YBbU5CHapqyPM6LwVUcsZxO9hYmQ0OSfzAcossb1+s1TOoN5QNoPoZWecrfC/eJ9hGD
9cWH6azDv727/7O+HEoKEblVC5nDC6+GeFCZf7pNcg1aBRaq+W/JTcyaCSy+zySkb46wFZeHlCRS
nsaT71bsHyN3kghDcQYGLKaJJtji1TqqFIjhsghn0vxMfouqsW4vSfOUENoI6mc7D8PSHnYo3NCi
z9+ggjeucLvqEP1yLRyg5V43+ImW0BADdpcvjPnMp1kSvNHukeJKV/deCUAetyK0AX8YFIRDyLxb
NHlRJTqasYF0HynZLrmWCgNwFCnee3zU+UFF2a0OIwB/B6BaHKfuIARDaUqRO4Iknw9MVBXIrHUh
6QMQh3tX9fbP7/ToasYjZ8H7jO5MNNEKWs7qJk0LLMLleZn9TjcMwT4q1PPGX7KmS8HgWyt6gZTj
RMrnvbTA6mWG57paYtfYdIFU98v5KKJxY2RjnlqOqe83Sn5jCLTMKiqINhGoVKJFr9i+Ob31mTMU
pGFG1IDHlEHsthYniqLGvmYQSt3KJcsOsqZQSNT2n8nXCpBPcj7/pdzT3baq1HF1yAhMZzhmzkml
lZ13P3Wb12Jy66gmQWKxPT3AqgV4wA6VQzb49k0CtiLUvniPebcvteTdsCSycKxUQbQFxxkFkB+4
BxVWlZNjlQla8MeQULdKphW/KA7W4anCLv6J+dGtvfJtenOrqVeALcCpJQIIC985ixh5WLcjVEE5
BWLiO3WKxVjJ2rxE4Ae9vkaJ65gdcUwv9yvk40AxfUDITxYcHdCdXHQ4RaLl81OACC8A23YYRfIi
aCrBrLDzSAOZvWczHKPnaxVimWTYv9DIQFb5FHBtsxrF3O6oknilJmzv084qugrXpjCawxz5ejAC
yjecv3TfDzs+Yp45TL15Q46bJE4DgnjA3lGG/nOmrf0qG0kU655AbVr5f/35B4nK/qd70BPC4Dbb
cIv9Ew0DK4a+iUwQ/pN+10oXkkZZXoH1PlWDmkh7Adff9gXCy31CQl1TnkRJLGUnHwDC11w5cedA
u6EA0X6uemkcJZLx8C8hFwzmB30UjUOR7ALUQ0KzuBVYsAbZTDQNObFlzed1aKkg5J44ZEwWSmm4
BXuz76Pwn3q0FM2EhqHvKz/ww84OlCEA8b7d5g+tmGOeOodHIXGWIZ/jG/a40Ryc9TQi3dr+P4Ky
P6vZdpZ8UQlVLuVMBjsX3YBSzeBqalsCcuI2ShHM21YX7H2Mk9wf2CtLTmCah2pr1e6ZFJH053aQ
+nTUmCxDrfnL4domqk+tfeV4V7GdDd7bzq6MyIQbYY20e2fMG8ExizCPS09AwVsVZpBQjVsmZoEE
XdGhka9y7IQoqNITnUrwIHYqoEOzjMk1ctH3UtqwdkhxT+2BUtgJfUCZK9XR0IQUb0qA09AFAYin
SMvc1CKhpWg9j2LYdk/u3rUpUkUEzR0Yuh22Yvh5i6VYc13oo83wnpcxKaXJCgKor0JDIc8LfdXX
sE7F2e1LRE1YnndaRQUS/o3vJfJZPvbAAa6e7sAr6c3ZPFjW+oZTJwh4n5A97WbWdGVmuhCvvjQX
cNMxJTJqPSYAQvrJJiRUE5R7c8wGjCAg4neFJysXD9HiqSv5UMc8ap+1mWNK8GG/NxppVLgnDoG+
idt8NmuPGYi3hmomu4Y7hR+U26MEQmtM11e9oEbtH5/embHbq37ZoK2YrmVWiESQESq4Cnv01fsb
s0HFcYmr1Gu/u7Na+NFgowNIsB/XAcKd4HTVvkJsjFP1Hyi3RVx7uIwCeUWBfKvIa+XMeYBt9jLE
8hLZcyTyE3MHYygmV4Fe9jnvEJJ6bJbG6m61WKsoTkrIost614mYPZQPknmh8gF9t0FG11zTZOwi
IWyZAzIzpzW5HnbBd3MrviaA6v6UzH5t83gRVRHmrJtGrAb+lab2kbO2K+pkHnQyha1UaEuIbPUQ
CLPvbvlj126KpAAexqbrGhiZmuu3NYoQjA2jSCN4cl/YwF0603tc78HME5fB7+FJa00V9pzo0fyw
pB1kIdrzQ/0GDKSZrPPj2foEN8fucF3z5+oCl+PEc//fzx/Z/N6PY4wfkZGW1fWk88nKsl4x15VQ
ns3qxxC/YA98yBLFgWY+PE2aMtTxSEKIeTCQUEtGgBbKsAzg+fnx6dITc/543DTSL11neMAYk1Ej
YfSKv2Gm/b/9kp57InXb1Bai67Xngfdy5ZM6YVphmxKn0QRbvF4Z9egBeGL7U2S02JQRoZ0tCWii
aWU8pTErjRVObn2MRG8wKZVlpP1qYe4GiwzZ4nhJPxZx/sSphPejb6Uh6ThSCPtQah6wbeQZLvzD
+9nOfac5YLdY+5IjoUl3Uxiqd0gRPUcPAyqCpkxhlJg0qeSs/S9c1BEvrECLMNGqu5BfJPXRDu3n
RgGOpqd09WgH3vM4stgd1/deMJPqLDwVbkm0/vT7UakQyU8V6AZIbnT0gUkWEZvyEAz7PaveU/RH
2I8ZgJNYsGi/pcpkl1YszX088GOpa3EsNGkASPJuCeBNrOY4Ykbr49xjzRvmk3jxn/JBFTIpkxox
TGwBeTKzS5JRy31QU0oCpbF9aFDZtsj5mfZdBlCpFuOP+jNjRDwQAiHBChif65hmgurCNmbUd+ME
kN1MnFK8YbS/0xWgJ5mcrRHJDJvJ3zJHDANqdQKD7YGcDH8OZnHP4TtPMzMlFUdXjABf0HfXqLA/
ec787PdGvJSR8RaVJbVDU0BCjGwlmSHcgni7zyKVR1v1zneYRl+rLAjmGlcTuPTIaM2Vbe9tuLQy
48QVmXSnjlAxC0dSxU7R+YFJBbGmB8F7gm36ubsec2srcgqSmw78aCSOn99G+7DVtgxX4ltz7Gt5
UGyKzmLNvMTLhAFFuxAodb/XqGDp53ri2+wVzJRs3PjbjeLtTqWdRgXEkPoY+m/wZOnKMAavFY8w
a2mC2el0L7/HEBwnydKlUA4ZocozZO+8g16JMDB4phOA5bzeXxpSMeOTehWIiKeoQ+6DQwtgztvW
tB0o/W1n8yXrhGR1dPj2xVV7I+dwdXv3/MboFx81NBHw+RHghjqWJKb90sHMyeZezdm+jz8CVx3T
bh0v14EuTbwm68NdYt1sZjLwAdWDuwFqa3xk/3IDAGNmmNn12lEXBRG4ISjCc+3jcB60rosWA0hI
6UPr62G5JGS5Tk004AVxEPBf57UWlZcEBTvT3tgUlDFQ8hYbCSS43zSmrfViAJoK8jtVImDpWs2E
dAVUPCK2qB1vUGAze4J/43nQK/qQ5UosNVENYc+eo4YU+rTvSfB1r0d6JuxvomghE8mQii8ra1iJ
dda1U/fNJuLkjKCUkF1YEZW55fc8iEvRq9uRczBLlZMkoxYVO29dTvP97LDt7f5pIvNOHY8ta6Jx
y3cEtytrKXo5802Ndxgxz7oSbR8wysc/v9+vgZent4JZrbd2uovslziKN7rSW97Gmq6r711Lg9HV
/p2ShPmc69IvvjhujVQka/PWewsM8AwzZzWYMw4mfkrX8UaIZWwHiMZCrS/qiBGDf6bE3AsjXybX
6GmuMJ7T3GWmdJaxBWiyWVrLAgIqPzsgPF4zC9biyb54WqQazXkig9NLiQnoY4Xep7AjUpBo7zkE
YpjNkD027dM4thHdqvDvvCFiTZf3wwlzcTPGA0JMd8NFgoFkO7rOnhcVELr0eg/m+Mn2aEf0KaSB
uqXNwpllPpk5X4/l2q6aZGtxp5742vgWKHJcwiKZwZPor0BQJpOAySZPVpd8kNAvN/W0Ag2oyFVU
05P33nqQyPpSZ0g8T30vdyMA97ybEO4eJYoL0QI4E33B6KyhApvgaKTVb3sk/a8ZCd/5SAOZlzgs
mZ+kc128smSK+b1Rr1erFJ4UX/5lnTfvZRI3dyeBEc1EXFq/WFCrywMGioSC6fm8C9W1OFuUGnsp
kqMZ60UkS0Nvw2XNs5Qo1TrWoWQPHSz0bPmKkZPbX5DbES6WAZbHwAmuYsFt74wJD1CA5s3oxtf2
P9YowqPFnqFUmWnMUZ5RXx5mNmMGiS7gS7tziF7rDc1+9sHIRvogOTN94717hPeXlHT8JudAY723
srLyUmfDwD7oUkJMZu+cY6fB/+d9GnHLqkBXZZjAGzGACnE6lGhkOXH7bLznr+RnV61sncAjvTU+
1nGQZ+fMUPhNkz4j+BriNYwll4mUkEEBMq9Za1dxFegx5v3JKL1coLHqI7rbypRmvvl8gIZ32Yf+
aBs6ap//M6VEft0OF6lAcowX4NwMyN8CVjBWzHQDLHVK/Xnm79nfLVUIKrheJf6lvesUPrUQke3q
P/LeH1HR+o5JaAqXeuk8rAy3n9tXSfZ+2MtQbthiDEu9MrhtbAMC2XrDBT2hObgHoMLi6d1cZSfg
f2ivW3TZCYN9pNMH3bsgQjLvFwEwCkoLGYzn0B+ksw+j/MR6fTHvcBqiDgun44YxpiSOpekDOc46
mtDvkwvIuLuu4vRWOpGm+SAs5+3IhsxZhfo65fdu/R+S7TadfyiBRM5SObXqWqM7/BdtUCa0xAxh
mzPihK36KUaQ8FGk/kMn03bh0R2F1dvkcDc0WMUfNlHn5cz/KP+1sw2es3WcleOvS16/2Yp2xUkk
4VLUIrujge+DOXnLi8tmJDIMXDwtHpcyNoFr3aQwJB7zwvtwLBzJDH/thIgFXLv8/1o4ZXbZ+aBe
ojEQ12G/1CiXpk0gw4wsO6OE7vKmGJ1r0YtBNhxkahDeORxvMESN/bRdJAQbnEyF6fdbi2iM91hy
fxojAGJtGZ5OPAxo13vAtxbJeAZuBy1Ns4l6tat5aJucs8l3H4YdHe43ANgRcoRGe3A5PtkDD049
zzzBCsctAtPuiRrT4rAPRNoeA1bRWfcYFXlhha1Cmj4g2NkdIL2vSPDRiMw1xfEsBM2iwzLqQHpv
r8HHWNFmj0oOP6RRhZVf9kBCKBK7TV+3ngXhYiKkCdXyrd5PKuCTdDwr4p6h6qefynWKvUd1Fttc
GqZnWSu+eR5k2JTlY34eJilvVWnWGdkIItLpe/5+i/XqCkukeZnx50OmCwElCc+gZqVCznvv8NOr
Ta3ssKkUot5gSmDDreg343CL/Id/CZ4gIoJkmL/K0UaB5taHR1B/MTTIGdwIu6124xsy+YaoPWUE
A5Ievu3PYQ/Ef79YCUVBNbf13TazNTJWu5s4KzvoaTnV1Hrl+hDpmsDJ2mI3ITYyfVLS7kuiGZJy
EjkYCjKJtFhxOkY3H7aPNxEvpgvkmN0n+E/44950zl77fGLHtYHsbxRdA0CIHpsxPJ9qBkhFSuef
5hMjg8z8aJNknv/3E89EB6IdZ+S0EWV3gev4sOtFj05in6E0tw+K5+pEXuFkd8GIKUURePwSqvg6
ioToJT7iiYIA0CAM6KB1Td4jAtv42UPOBGGfuX+Cr1/k1ln3JAKtpfydQFX5/Q2M3KLqISMgyMsE
8Pyr24I9Nhes0OLTywh3qJwgY9SyE2Iojo41s/PikwGfrbRgPIrxLiLTrMw3+VbqeauziZMF8iXs
qAbOAYm9o0EbTQQIpX1Edk0ppzlMT9zF6a08TQ/JhaoQCMCvKzKhH7cu/W/0wAL4Vr0icKdul2MM
jkITGVFlaMYA4NTJCwIGUPWiFAFKpZ8XaidU85tZ+CvIMrUWa8qIS8MP9D0KitN09OwXbVYrjY9/
MLE42Z5XEAsf0YPlFL1ApoDfPtAlgmCaMyFNwdsRyP7slYCuq8VLahlEVDQH34uCbpm+4yRYIqHM
f1wWJB2w0xwYXfCnrspwK1KKhtd3y8oBlwrGLMXXwpXsCfagdkP6IL8NGKuzFwpe1IalT8QDcpeu
JpkyNr+fdYjl/P7cnMs89j5fLNMIqZX5njEgi4+0mYku58+JoKRIC/NqAkvakvj6H8kICa94OqjL
5FoFkicLfLdRaZbJJUoB8BIyg6hqgt3ZJQv13Y72Z5Qs4hO1aGfsE7rZTGMWCaPnbIljHVejG6qA
MFfBjR2tDdmYhjfhgFxehjUvQwj3wq1xS169vwWDZGM4kwu+8crYW2x2tSzyIDqaajX2GuXFAIg9
2vjSo5sFkQbb1nhH/HKzWkNv4XK2T8YfVYz9zdu1C1MfMHQZUnUEVP9FFuemLHbOKax/YQkizhvc
A0jcGQ8VgpgPpynONGsbyBm/AVtiCMwpo8Ii2d+8kZuGVW4wmgYxMEXS0F+apUt8NdLyRRTe1+yp
nNxWnZDOk3AgyCoPSTGlBZLjPfBYE/hIrwOZ5qpJBzCayXIyNtpJsd/XbryjQk7qCrzUKwNaFn6/
IyqgQF80wBJcfANgyXMItoou645zKw1AchFeoh4V4eusgBfCgdMBM1mZ4AGT+puz5y8Y9gSV9IHr
Cuu30toBbjUvKhjhGzF0oXYHsWyEkLtR4lyKsFs+ndKG8q/x9ILmyNHTenQxCI6N2kcNk5HqCOFM
4YvpXbu1fLs8+zUxYftiPEj5EXvwha4Z24yaJgk3oXH0B34RrJF9WMclVkkOiU0ln5SKNHZPZxFq
gJr29hDgwinyYZSNpD4O/umdgzwMsHF+YILuJR3/kvFCsSTwAxliiJXbPlmDE3CHqEhg9BDcTN2U
quQbgJs72rjKo25se6vQRGH6FkiDa1mB1YrzB8bQGrwDoAxMxwo1nzPd8L1m9veK0ob2DBwQFyJq
Vg2FUgM9kuLxnZL/kWshor6pUey5LbKw0zxRd9df2SfKmgo9oCFm1p+hqFhJb1eAbunCwjeAASpX
0viJKHqIB5qbfw90fo7AFYxvbvJBIpRdacneesN5uBDvxPefsi8XsoU+JCt/U3Wi75dsdtAD6iro
hZrNRRkLJQm98LDeWrBKSuRoyNOumsbK3OWJ0ozyf05Qah5CI3PDhwarHmt0qX8RAHZxZiW52nYm
JpqVRocqZn1d9bpMkD0NzQiYCQig2MSEM0tFddsrvYgLxlph3wLbH5pJ5Dbci7q95jeqgiGdjPuD
hfEkOJJevZAR0I5hu+xPteoInwNt27QgHfC4KgFzQr484zcUDy9NwLMC1LTQxhRTR9wPXAEU/gO3
5UQa3O9wQUZ3ULekBZj+oBl2zOJOatGIRUjkmRPMb8vf+ihJzHwAhCa6KPiR3RDCP08eRlihoiB0
6z+FcBmanGOOsufAdXPMdVQzL/n8c+2DyDMdNluuA5Z2Q3Rq17UI+dC2JNklqHgeS084C3Av84Uk
klsKP0lrVIzK9YnXUG5RfjsLISW0m4LBSZTkr0fHMgdCLWmGa/s1VntlAsgvIJlvunMzgEQs3ujX
fuzt/ZmhL54IdNUH8gtT7u3sAzb2lsnmH7zju/RqUNHM7zywLwKIxgBqjB5G6eHCo6iB8EAyWQDO
51OHpzwD+GMPxiz45KA72UNMEdiLaTgUBzDXVBXij7FZ1PGwKkFXclDaFHqiMb7IqoN5SuzfIoyp
C5L8rPHu0nH55ILVwzjgGksVlU0YhYCXMIHDuTuNkN+TX0S9HD4Q05xGYmQvFJtDWJkVA131gBPR
gwy2S+DK/uKM/G7vUCLgnKsXOC0a7sp+xnYwIPoL7sx3H/zMeZ3Nnq8CqIo4kkCUAFO8OrIwDWLG
Z3WAiS+mG1kdg0Yd8b5rSK5ZrzOO6+VSljYmR9qjusz67WEy2ilCr6CQgpbjEn0DPr2w4wv0Cw2S
6vNuC7YckeF2U921UX8PPyry2pLfxFXsonw3MIOeDjG2mQ9UQsEhyl+qTxpnMPmmuPGZ1etBkmea
kviR1039G6w/A3Pf/P4HAL3yDltu6daB2iVdK+Y8xhx4HYFdaUdGz+nnjPFIcqKN4iOdQHMxvRFx
cxx0Lm/xEqqS5m5B0NLfGFmTzy/TXfUhFwgFANDOh0q0rA3cBKDU16jVB6z/cCRUZaiDi2wy+AcI
U3jT7iaOVgN1xKqjIzWvo6N4pvHkbdk3kGEQ2E3kOKG1iPnmHOBp+Z0qjr4RXNGf5L2XZjq/JzZM
5egLBXEtL+3i/7UiXzkKTpT4bNUNXO7HiWC9JsdQvDEh9tFTbM89AQAB09j/1skQ290brEtqEgvs
1lJk07nlTK6JZ2tQ7LzehPGUU2Am85n7cUXGYOUVQRkzjvo3oo8h1uD4+sA9WcjLVYS6HK9b2Nrn
FuqktIOnIVMvjeufskD67dARSp9iRtFfojcWShjBWL6v2nY5MTCajVHIqVYQbihlfYaYpa08Gqkp
eXh76DFKXSau9kTSG8ed+IXpdbcpIvfzY5o+0l0J4X0xogzCIzwx9HyYpCb3CkjOdEE93jgGYNSj
MxYIcxV0/Okwqt2cIijm/1pbmhauJJfqmGMVPc1dHu5lO3osZT0tfsy8y+waqns6m3rPY9Z3fGd6
a0j5mVJnjEORnc9m7m28ec5Fkq+M9Ym+LWjKqxbMpx+Icb8cr1pBF8qbDSSOMHMqrZ4eMMjKkGDH
P2bYNmr+rmUm42RJfGov0Xpx3AHSx+yOFp533PBEj4g/34orBC7r5AxEvhxzN4yu3wxnnTRMofAP
jCTVKca46cbOAX1voRhH/ZEJYIFMkiwJ4GAyXLedNcxXcaoCMKfn0rAml+7ylIy/KYi+wh8sdSvO
ZSy5NmZ9xZFkx2+gy3IjBcDyPmENV/XgZCEO04BCwqAscV1cjrPy1X0N4bgBLkIRtAgWJQcVxH5k
T9gf0fQoaOrLB1Z+WU/mAAl0gAsaP7ryRF3qtXne2+WJM0YJFXQj0hmVkAFYEYmsGhEbfQpC6NyX
EH5zPOPOJDKOuE0zMIAyPCGNoD0sX1XHOh8FuungfIuXyvcdJpCaAR+bNJvKrfBzn6UFOh/0rU26
olEr01GD4cAstQXDF7/jNugRQZPwzpNeudClko8wrV5fVbpFVtP/JwXe41RhJ7UcLUb22dJeGJHR
nMxolx5Z9HD2T19GVKdNxfYcpY+zqDtAxgRCFkHf6SayHlTAeKEOZi790KMX55FhlxUUK1WEH8te
rF8v6m+Yhps+mDLGJmu32zuzxs5DsNfYv96T76gZcGzM1vHfiGR+lv+1dRhCDHnR6MDKRkQ8KRyN
Bfta5q5aZlgcEHDYUeCPy+UI9xdF++vTeS+EZVcWQ+MZLWv2ldV88U3ZWRAAy4It9yrpc3nLsotL
Yv91Mr2zizubW0gOyrnMl/tlhfvKvTM8M0lBTVRkQTPDBAC700grXnAIwqH/f9N+a+l6LM4PTKRI
+r2St/TJr+h31q9XxZLzZqqZnRkhP7k2r+g/Cg5A/2/LctaLrkKPQtsd7lLn6jsdfeVhFCp2UaDv
S2xV1xglsgiF/h40giohzNpF5RIrhISGrlWQmBuc8U+86acjuGHrm2jsRmjpZutpwyZ8if8CmmIh
nAZRwzoBgDp6jncIWTnLHQ53BPuZkZA8z4hdjxMprR8iyH0zQUIM3sA1CVhofVksqylWTVZOF5Lz
V24P2CRuCkhWgEz5JH5H5VdagrEnfoN5GwZkzGa/QmiyKwwH3U+wHUx/6LUaS4yaxDxtj2YhFGBb
3Eo37OdDt/vfH4ekeCCsM1rLrBD57vPq8OLWoYemhhAZkhOQ5t6qMwH/HIgtv2AMb3TrahS4pJpT
Ch0dA1RFrFHpxk2q1aAFv7OTRSjATpoQKmfWetVPoCcKiCqh3EFQ8LbnLrA8capgd5i+S6uRha4S
+T2BL+oGPFiL6vk2PKC65Fjatue6VajJm0Ri9u4Gffxa8CTSo3nY42PVdCuTrKyDQKe67kT2Xv8R
W0aC+MoaW35Yt7NWxQXAfAe10peXiixRpKWlNph9PN77x9Ci67tnQjI0dvQZSYRfu2p6KXF8BICJ
xYF+BzOr2k6kLD5PWszJBeB4k0D1E/eDgfEh/84LWOIZBQ6RJnrJBbIWc8eIt64ugT/U1ejzqwwS
BuF+jNKrhy6ws22pZFkJ2yBJEiBwGT62xmp5cgShUbOaqM55Pxbwv0XENtXlumvhU152hr0Sqa7P
pggDT5s3leVi53KrooZkJOWwc/L/KLfkp+XwRAj/Nbs3/o6NZA8w5NHYANbubwSOurC7ADbMAETR
HZjlLKTrReO/0O05yUbGIXezomKRxKGlDyudxp/QMNMyiW3O38XZ68TYGTvkiNla2WnLqBG4Ahfj
cj0hPq3JMDZViJt8FiffxoUztEZz595GveUV4s10Ys/qto5If6pTACYFpW4RbLb5S0zSJPidbehG
jAZ+C5hcU5Y6FoCyqtCy4aJEHSohPTaw/UpgG8/NmhMnefoVlxP2iUt2sw7SRbP7Og/fC2bNfFxI
JFHZnaMVt13VvQZiYHPuM7vA/yMF7XLB3XT6zUjnOVhyq+pYSdu7D7Z8y/ptXZ2HsriWDxBFEHTr
ipdsfXFQnafZrMu16FlmGbQqbg+BEKcYIFTcfVb7vVi2Z3wjjXBlnXYiFAuZ/fxYqtbMWaqi8xVV
cOJMhd6XAFcOln839ywq5l4N/ztVqHAGryUjev148Gf54B6kyrkez1hX1l23qCu1moUGuUYei4Lu
XnMl0GhjWk49+huOrqS/uf49Lbi1QGtdAwmWwp71+NhQpNH8FDF5TSkcv9MWleK4KiNqJTCcc15s
3w4ZCT7tmhgGwAK2mrjKbEaxZ0En6FC1Rq4kzzWCOGv8rRd2fPXFeWNcl50VdYsIG2oTHgxAtMQ0
6yTB5QDsgbDjYR8wbNaZFLetqJ4BqFFdU+kJsXO79m0BvjOUHf58H5Ctbg5Uta7N5oAorAwVjkdu
iYFzQI018acKvCFXujVeD/nZu5QbT7fCjmTqc3FQV4oFtF9RDxEjflRs6D8U8XiX00+2nK4Xtr2K
coLLHeWTr5n5dq+myTM1yUaQ1IUoml3/3LIvhBG9kmb49H7zQMWbpYAllr74mxZ+M7EYfstMvZq2
unE+VBFtZCANPMmDM+JYvyUM6PvJn1CS52uLttmO7bihlm8otR5h/Pwtmegxf5mJyA7ujNKFrQZR
gLqz2zuD8YQhcFSc2lM+KHhuygowX/5Pbp9Mesba6XosQjjMn8cbQFdeXGgtR975/1Ve8RtdN3Up
D0+oSiWh97yj++7DMsQ/Xa4/5eOHb7IXW6H9YqduM9EBxlAxaA578evmfs5X3aIMmk9yqz7shEj8
dcGq7j3uK89MRxqK1SwkU3ibYjSo/e5uwoY9F2ZQlHTqF/a2ZjbuVb1h5u3EZZ9b49ajBJnR9Qa8
BgBDcbmgeRIjySvcjYjfF6ldgOBIAYs0yPNkamM52o3epZWukIp7uMV73xeyhiOrpwnHqpjJYkLM
GLVSojBksXolxjrCc9SIMDDpEkHpjJQmzkMMUbrKQeS9ac6S4XeH/uxvszLj2Eg/PYe97YvzpdJj
U77WXewApwyPJZKYABhMUJjhljf+aXuoX4s40krxiMogqPfEm/fS1GQ50/EzZhDfhr+WQAtew9KY
6axOL1KcZYLOeE8qcnye/kiuGgd7R0kNidqfPnBn8/X7gXk4Lg3jmUIJRKMINY5IUWXJji6bZ+gI
yc72huYTdETGn533OvXPhxdRDi0KySvVbFnOn71bQRsIEV6FtVzpHPH8xQEQKXnxds4SBvEcwFNU
3SPNaYykqz0PqGj1fC9DFoCg8W1abJ7tip/I2E3Ky7l1wdzWbiEsOuDgvArX551Yw3Id+nqORi4l
3VVbv83SHz9XkrL97pAzbJPOqXkFZY3ZVzSQlBGaGOGscjg89btC73v3luezroFoh/1lJ3NGLKBl
W7NqtzeersHZYtW6ba6JNNTiLnTamzD6X1x7waf/xF6cLO25VUNe/rWHVIlD7O0ixdmUqBA+oXlY
+lzYwPP380rW1vJlkRGZOwiBr0uwDHhqEGAQAtL1gaGJHCxP5F3FFgnsVGVd/9qYInRXaSYHtiaz
NEourJFRSevzdPvRfzT2TVBmDtsV6fPk05qo3f3Hj4P1QwEGLUmv4syK0a7a9zOmNzDqdLsw6Rdo
w2HE6S3Usk57frk0Tt05KCBeP34VTDPTUzTw9VthysKMjazCEnR+kNpdKSMxELFW+fTSfeXcWhv9
mkecvdo3cOEsH33axcJjbqQSi/NOi+otOzBOeMfMSVcSwsnC6OusU2kyoWXgf7OTHKBW4UYrr/Ln
TYVjVCfygfhoXPlQZCOancl0puxOLHAMjEZdqYP3ZtXOy6ee29UYbUnLwL6gxmm/8+x64ZAddyHR
vsw+KxFcpPtMjGfMfBfDe10SVGVFMFWAsBXM7FEhwfeOe74QHyh7ZklESpE9OQysYNutpB3wZQTi
Rf4hXEpm27bKP7Y5y8TCjbkzYhH4b9F2G/l7jXfc1EoCP4u4pJ1UASmNo2m+6hydlG1P22UQyrdf
cnlVpFN7yONV9JGQtaWGTZGAtoKRFXEspPQg7pasTwzeMJabrW2D7hLdct99PQVsvsFGbb74ymM2
6XcvaPh93CN5JvFweNgugrjc0qjPEoG4VtOVpC+skfujyxriJde/ibqpYaM012zjWftuVJc6MZ30
MCOYcFHRS6S/oId/sAJnK/XhlHmOwyzD4ZEL6OPgOik+Yx0CvHkAywehWWpreFQut2Rv+bgekFga
VkCIROWQA69PYtbwmuzx1uWwLnwlnNnS+exls6Q+Zk7bD7kgUurSV2WJp9n7QuxIuqBG/jj7Pguy
kNpPckxvIocKkduwn6q2cn7DmBGrveOl+xDkq+/XvvKFoJ8LlekePrxDbfpOULwOVchWbQF4dooI
+bLGXRIy1rZXEnN+6NNh/AXOfLiiwi1rCjASa5vSowbh8tyMrhkyQKz96372dRbAB0trg4J7SH8b
U2MHa17UNvRajnJiWR3REdUpK0nuUnPxvzAhuKtlwEtzfXsyKP3S5x5TmVQLjWMOx+/v3HvyZTQj
2bplRdGU2XmidQZ9+vgbm3OcIOoAht2WMBABln/aTD3xzpJB2Z6LERPEkmekeBeqg80uZJzSvkIJ
BmUTrm2rdWjCEq6E17r/z3hivEXASX4NfQgRcVQmyBdjr07bYiOl8xkH3WKsNFJvUEVU0LJKv6KC
fkBEPnv+1V8ul6tP549CUUKuV11WoBKPEqSRWRhNuNovTXcJP8qMVCdquo8zC4jhvAwGuT9BnCKP
GMSkZHvjwU2dXKoX+upNyV1gCmLCRTn3m1xoAQzcBc/JV36CrQ7/lV4n+AUT9x6BBr09Dt69HFo1
bOETVHJXitjlR3pNlTYgS6mB/i/Fr51s7uG4Ij9CAGCrYLBOVUqthZmV3ib6JGDXfQJocULD+GOC
QPwjCOXMNnNFwEEkHoPL/cTowxSeqzyK0juL/6Sjo0EDOTMCUhIXabRuETJk9cQLbZVNovGe8us3
K2H6+XZBiXavPA8hPTnMtb+gfl0CpCb/W0ZT2FrVcoFXla8mP2BaEhkh1cqeS4sdckeS+BbRTzge
b3k+eFiUU5ZQmjN1Zqj2mvVjdCbRgwdxAsB/qtDOaYunhMZP4XVpeRcJ366Mr6DAlaARhfKQouMV
EzJBiDao60ySdgLIBoQeswYtZSAylaEHKXqBAf9Ftob9SiFsuAEoWaUfYhvh1dQK5JpEtKSox6SV
Tfu+s7+71hD65WC4wd/H2HOpg6PRSQco0J/jbULbbecw1DecmXDLwDLp6fYk37CyLnuTKD7Z4Lwu
PCkdPSCFvMBD98vSLTAeIpZ6umD8rBDxRs4N0vL9kueu4nqakWyBeh8zGO9Qqitct6p5UPTi6xIo
dE/Hn4e+Q2X7hcobFmyu6gviwag2g6C5vZMNnZde5tUjvhKtWURjKUM85YLqvwD4ZD+56xue3A+Q
caSdi1qyKKY0rHbOVwUt7yqQhHBYp2iZkn2ZkfuFW19iSddpDCX5l8yd1VBTM67ixWEkBR1SJIZu
TCgPcB5z4u2LRfANVmwQgxDPvK8CNrgfvYs2L/7HioAdo85VKrQCVpXwo/YPii+0jKcTa6Epw7RT
qwcCR/+yHhxzF0SmEPsulWwUcX6FWfH3wLetzOP5vYBsgZHVNRbmXoKWSBV3aa6mr4DEygRSiUGQ
TXl1S9Vo+mp52psnEmUnu34NyaI6gePx8UTW/gHKUuDp5peq0y+4tiElIp5/sy3NZxqvJBrpOOvv
5eYBTY81btloNvNlkiFbtt0uNITZkVFDlMxMhJELoklHPveMwMXawN4fgY7vju1RphJOLOORJM8z
dTc2c/8T3bX+PFdQK4DbpohmDMp23mttzMGa7o6QniwGawE4VIeryl8VlXaVfZ0XHN4YaqFswpFF
9VCj7qF4E7ZmDnVh5zJok8QTqmIEdwgYXygCbTj0Jsyy0PmDAlprrsiJ01IQjMfamM87PFZdc+DU
vxxqmYTnXzJLLgxIXgohK3qWAIAgC+h5FnwCJ5llwXkGYwzmck2kSLy3cJqbnE62YxpYCTI/sIMi
v7dLVGW+CmZu89KHnPR84m3vTT5cqMXlToorrIB//Mly6h0hv0FZ7EaJQQcAAsBC4kEyWcC8+k5i
yXApTnmAEnNSfRCVCwuRr4zznxkl1TFdF2fO7KmI7+2xIa2ZVA6PQfpfKSzT5LZNSzsR5YLi7lI4
EkYHK9UvCfw5ahfI7GX7Vkw5Ri3awYTDYjfQd8HoeAeKR8BgCZxLKEDwC8FBgu2SikZts5nZEcZ4
heCtiui5DiYZ2Fq12+Qmhhalbywns4Axj3utMg58IKnOVntLUjDNi9zljj23TGyNa/YcGr1mIqjI
1thdOFryMVdNh/4Uc0B2sY+6DermBtnsvutf4l6DVMBB0ZP4rFpY6ykxbMi5ig5XIFlA9muapNKy
hHG838SwlF/V4tUQm5y/wxpRJkakNhpdW0uGOE3YrouMIcdHVrK7fPl7E66qO7buFiHJyFnljgmL
GEoAUGhvLxhnvFtKkSFvVrs/wx4TX0Zr/xXT9cNYbV5C9FGmOj/NzHEnEXmlILxiKUAJdPQLOz8j
JXzx5bhslQO9vySIjIFE3ZnlhK2XvrsIWkg0CECP48ckTd5vRxVg/mob1LsYmjor96x3T0vhhUUR
wjbQ8yXe7trHRIGr4BvotSoszMmqzeFx1USXp8qEiL1ER9laCHVe0nAU7tNej292VcZSqrkEzsoe
Ni/4y7p415zUX2bSlvv0gDOUncpgoI81lm0lP6aU7dVMM+8vMsLLC6ITsmakLA0x10eOSjbAiAOa
J9SRFUrJDou0sX4Ue8SzMreJqVeW2Ho8FC1gHBtdne7rYA/z/Irvc8TR4laQVBgAJkImX8ssgZ+N
QIrK6SHCY+ff7v4yOAxp/qfoPCKmQScgvfkFEZjFaHR389AoUyzJZVio58O8HlLKMdr5skMmFIDy
qLs1nOyovC9tG5skVnivIpnFOMUE4GhGgJO11tDihICIdhxeROr0uFL/VILtmOv5hcRkxz6dqFeN
uITvf4iq61g50bXER2+P63Vb5BsRx6adKIm1zip8hiRxtHgeo2Nmp8kW8CEVnwG3Bf5OA1SoVUvc
odoVDA6qemaKH2FMjEul+6qunTfuUVIpp1X1smyfz0ArxLwRZr0btjEBnW0KvaTHRixrIZlv8Dq2
DlJA4FaRNoJSp33g8lSmylvd1n8lwz1JBT4ki/rjolAUA0lo93GEeO6OFan1grd5//WsUPfzOLBI
Qj5fxNjo+s5/BCMfhDPj9Q+AK0Pz2rXX3bZ/yv//NQ5onpt86yPGqeV67FAsasJqnumCz2VDfmhN
gvFl/qai7KvLTl1qliLrnOx2dCoVaKmxiWp6l+efYNF5Y9Ys+HvOVY6iw9oI8dllzlm5Xj8cAIih
P7+iEUHg021Z6HGX8qFR5j16DIW77Sg3a5X4jGXIoyP5+4PpWlxTUbOsnAXsMG17OlCHhaNUwAYU
e2laNwXxJGqj67+0/qfoMLiOmIt/7pxWgNfnuYzvDdgVgz9LH9tzg/FP5e1XMc1B37R5lOotxpT0
m+CFNhKg80lkO2f5j2uoQktFiroTUnGKXIILLs8L5MO1hbGyl6hed9orHL42bkfVM9qBlgI562ey
jr8sn0CQguQaROeAB47NXovXM50uVcAgNAbMLwNhNlvUc/PyEnkxeoB84HBoVK6AT9eX7alaPtq5
P4iCmc4ggfztCQVXl25YbevUk7EoOSiy9j4DvvVS3+qJkSPc4bIN/Ru7CJ4aIe3hK9ot4wZ36gFl
u2tkfk+fxzTtfSEQ3z7Hlldq8N08XikgzkhPEj9S6F9bxQXR4gGOp6fqOh6BVE5Bwd0OkOT/Qtgc
LIRa+JnfhZhFKYgssuTDdrbLbDGybr+54dK2/WvqK0m0fo65w+t0iSI1rcQJE0IyOqAUksmRhsbq
GZito2GbTlhJFe4OLM96cTlEzMjrvnCXXaOs9nm0uylPTHy7ZBRdeoe0iRlunIGTA9oHOfPDu1c9
AECuji57P0TVgPNQyHaj9PZ/GNfT8jxSYJT3IfJ3ku//17tLA4gAirfPGrluT10BlvZPRiG+6MuE
YJ6lvFOe1jd+XHXDo2J6tJatUr6P4zfOo6gHPV9z7EmFf0hZqbKCDxa8YqyoFJgSmBfbtp8So/lM
52dTty9ri1n76WFi18kJA0PeR7U/LjYDIETlhSVVh+9HYOVp6Ir44Fv3jG9Xz84VzTf1vc6rEqle
snsVqtt6PKf1wAvqN9/7EkkmBsMWqmgp54dpTkdtHq2MCC6dQl0hBlq/3DBSe9vGcxBOUYUhABjJ
l9jPg4n4ubEr45flz5DyxJSMrbfxujRURJcn9yfWwypc8YDbyK2d6/u1btyiYVJ6n+F7tXD7U1eN
BhMHLn2ahbWVGfswPlxdj5cKWJ/FXc9QfYZpGy+WR/MnK7t8dYzzbOdA1ivm84yjX1PKyWmGHv0I
AZqdPGECfxm2iNQC/RcWFflVjsCulVpfgTlvemUPjlyI9Y8c7sCZkfn0MzRk+tcquam1FDjLb9Fh
yoEzTJ/D15f/2DqFKPMd9+zcCj7jwH3mBjabtLqjIyfOGsM0ZqCbSEcp1e/QWSL7/MucDE+JhFD2
GzR2ZwXFsd8rUA+p8Xlkc1lzgYHGGLLKI9bL6ywR1ewJawAbfKOaQd8L/8X6U7oKtHdm5D0wRIfz
PSHZStVJl0w4VHrmfmahq80twQHakh9zK6iVrgSYc7MV1cadlRk+c1AkRMRr7Q79L2rNNH93ATyr
Uo8ofSaebpreJlvdjPKbTfWWK/BEUzwpLrATwyLwQDjaHFNKTFvxAdV06ICjpIUzNLA7lk3326QW
giR619+hU8trbfWqwOHXgUc0rEkD1x73Fo02ldhKbDsis+uoTTXPQdkuqUCA4q9itUqy74ifv/se
74CL1LzBaw2BjA0iDRNmyMdPije5RMCaWi0CuT3XHo/cCAsA91lK9tiTRjebYj9NsDBVy9HdBTZh
DD9KoCaOtPUnIOW3ZCqjZzgDu9OJDvKcJ39irwHGbwd/rOi2ZlUKhzTX5DPeURXpBdmtTMfNRjUM
cHNrnJIwowej5+IrQBEZ3zOXxpQ/Js/ExxoUtzn5A+CE/oMDoyzWDvtq7TbEdI6Th4ttMZXjwhCh
WPrCUQKHk8+n87KsIa++n6k20ipkBnlVPgvECQ2Cc0pSRqbssXK6bzzyX3WIIJehdp81oBeLeAoG
htuOZt5AS/fuyJ6/bmEMbvllWsa4Wkv9Ahyi/0C851M3hvdCbB04SK6nZHOAfZ5Oh+3Cn/QXBmhE
KXJ0QFntBe13PGVAi9BAyZRcVmLkkz+NALBSdQUn6d36Q+SRE3pKmdJ5nTw+Ms5Z5icp69alD1zm
KCAN3dW1NE2RVuKo3oB+D0U5A5zs8f84oSsxLVaTsNrwNWj/99thNhXpvuNlpRm3aXwyLDntr/ur
9BXDXz574UK+2kgGE/KT71ZAE6TRqCBUDqSMb6MtttKTa8b1iYcvZlGDIr7jUbdoMT/MQc0gYVPC
aL2rFgD9g/7U5PN2ig6rWu4+XYyjRXGLJpNE6dq0bmBu+Dm17OeeFKMUKi1MXFEV7bw5cfF6BB3o
PunGFASC7uSpj2ZhxP4WWIWQp6SgXtMIbcx7/r+VbqPePzkATUFW3uwTaRaz5hcYoSRbduDbTbMd
bfLxRJA3GwQyoLLIEaPsZWYbrA7BzlVMIlMt2LEnL6B94ZTdzZ2i1xHyr7VCCdf2I0rCX+Q1zaU5
uT0Gp8TdXjw57uYdjIxtGfdPWxWX0kS8gdQqamI6fJisTahNMfnpWXjN0mVipJX43RfpillTjY/f
gAFRraDOEE425HxUh7XfXHyBklhmy1wu6pKpAI0EqoVH+965gvLRjHf4h8fUZxGr+xoLKH7SAJPl
rya7/nK20w7p+LIl+G4znSHBMvg1nzg8LHhv4vD9e3Lw5LBfA3AeWrk4R/B45u5Hr/U1veFhNcbl
0tX/f0IILyRHbOoExewrdUfeklpVQGkpzrJieYdDiYRXXRttYQvqosStj4/qCx9psWyxjJfdVqTU
pTdVE24fau2c2w2ycCr0JYEuhrR02gyTVj2mpOmo7UuFn7X9uHDwuQaUONv+Nxhq3iCNyVO+jkOc
wQwEvPB/g2IiIx/CjZfTz5PBdw7kcr7KWHHhn844OKKI2xyviDlkRaUCXOBkB8gcg2vPLwXtYxbp
Sy5iXjVPVBCF9wEwd9qPRm25+utBVow3lRtF6QCKS8vb5cSl186JfgVKBX5ezyxWcXDOgKErZybs
1s+lV4nASUmroRlqXcMzcksEVrIXd7S5wyFJ0AMm/H7z1lMJIA7xSgtcM2HITypCzShNxyGj7Coo
Mxr8e2718uEc+t7LSZ8gyWMtMR/eGnyG99QEebo4Pm4nqbr0Z0yAhZRPHUT0FvfqTGAOzIaP305W
OhuyEDX2DeLJphl50vk+uRPJMHPv8OL5qQJjihJrrFfgkA/quXTLZLQh6Smlpe2GxcOM12tFCxzh
7YBiuKC3XjYj2l+fUDjpnC4UljiCQLnDsNoZ+dgFFrPhHEXanPGHOPcyGwyWULkVumstglkkZsKy
+PTi1gi5AqrFGkAcck4OUSC2HDSJnspV8VFM5Nfdx/WnnPMfeZ23ZPX0NXtQPPjDc3M7zL3kvGzu
7yPgx4uALVUyUrHZj4YoCU3sR3m5CVDcuTvX+Giuzw27LVQxvJeOy4su6QvWRE1k/BDAIHJPAV7W
8Mt4mfcl6FC59byq3iJalTn05aUjsZM/uvLNYm+D6L3S3Kp2p+1rud11SKfqfMat3hhRUqt5PbOP
u5vGJvUre8O5FpO8Nns5sU07fyftJxOLGNkxrSU7zXoDGQj97ulJgVg+GIkdLDsJZKjUCU8mCkUV
F/1WK4QLsntxldaPexeycBT5D0WMEkig6xH/FRDrDcSW0sT0ZUaHRmv2tilZE1M1dmIF16QlF6iA
MW2DQ+Yw8xukMLaaQQo1gcgoG1FWi9Wl0EBpRuYp/bhVQtor6NJR0EgaTZdEOerFxOiMOD7tKsI1
5knqDfNubNCq9lkBxp+QdSui2Qv13tLto6K4+Fx7V17v+9hpfQ5OnfpfF/ClCoe7anxkT3zOrCsC
54xTYoRp7yWGWdHalKxY5LoDWhbTB/Nbnsb6CfmzU4oay6u36r/YnkyQ9SJyn2cM3L8xZvatoAdk
y4apPJIMSw7Imko0CM4ns1nx8EteVYEg2VDd368yL+6zUrXm2r7eOh9poYBV8jSgOlY+3piQiBj0
4pCzLd5CtxNdwzSwVsbYibYlqZcL3z5cc1xFtNWENt+N2Uux2cQdyDlOaG2w5yfbWUa9l1QS/huV
5vM/uxWLgr4KSHA7mS65FFXAkukSTwXclBqmh4lpH53l3ZqG3kQhE4wkTMZNl78xLHWGfMzG+yCs
kDRFPZt9wh8WfeeVg1SQuNgKV5GUnMFZYRxcKKfqjunwcR3g2jx8XSgJt7c3UAP/tPZOUjWYyQNc
LtGPvGtkgJnRiaaMdks7mbdCvI/XhofMMFEfUArFZwW2Tk2NI9HDNMYOZIdR9EhwGQe+8BZ88n0I
JIS22DH3ZjesxpUHqk5mC6KNpd4Q/P99+NbAmNOeDDz14NFvd+4cxpHi+m6OSltUcyNJmWiu/5Ya
Om4ATu4+EywR/wSMU1U6LuIw/qgmzfj7NTMzlK1d1Jmfj3TE2bZwYZRaF25sKP7jYXEc/NnEqpnP
mGTDTgSnk+B2+F4ZOhErA6RgVbx/uhoUP7x0FX4Np7kjKx1tenhdIJRziUjWspK52DkVNlJVodu9
xHPm5sy8R3YAEJJl0VeYTuOad7qzgF2ljQfbWz28ZD7bzuNHmMGTD+D+/hoXDlqdmZi2Q1wnCnJs
qVAjcAG8b2nJ3Zlk0DWCDpA9E3DP3VuMxqC2FHwEReXqAfO5IPriHprlotB0zLMKJoGPHpKJGjHN
ioEprCGaWP1rkZonIWJlcaINFIRWD2MBewHmH83HkFqSezlBmBWlxViwZsvJIiwwZqpsEaqiZt/i
TfmbGNvzAbdvht9wdMHsRRzDS8az0orfuYfiU1MiOc19b7ULSqKiXhE9lwmoqIUMwULPv0LzKuIz
masO5VdbO6YKWHM5yPMAlU1AIui8Vv784kRfSd5uXeqACQrIjl4XHBkeCZvwoDygoxA5cCzqw4Wo
ap11IgXrYdj+YFTCKsm/CgnWJAlTHa7+KDEFjHqzGaEWI3fTAQJlyLnKkYrhenCzOju7N8A/9S4q
y1hor1B4XZKKVrd1SD5gK3jgnXkiH4ZYLPz0x3PIrsKbsRUfPVgIriV/uylCV6c+arrBniUz0wGl
oFC4ot/XKLKpzltoMfud6q9bh5b6Qx/SvPi66YWR+G2L8Pi6thXUq6BE/hr2qkoLezAjsLRPjJn1
/PofwBkpgoXXBB29McdffuxxLw7gqskn0A3ihRmHe7VyHiAcCP47/Z96mMa5chdik9f0cYhrO69p
xfaDC0439v4YMulCiZJgRXRVyo1UopVTiQWB0ndUP0heNGH4768BW5mDewl2D47MLyjCjRDJOvBI
y62n1mZFyVhwubZlkell31Kr1QhDK09nA3mxPdP0wDKiCkmkE3xI+6mMWaPTZ3SfWzyOTZQaQmnX
tWd1iiE6ALoXhzENdmmBNyRzXykleJZ8f5qdNURcwBoKEiRIS91IR1Sbhwt0/Y8shNlMjsZ82X/g
xCbsjH3Vs4whzf3zPH4iARO0xl0CHfyxvecqMfDRcP1orqvtWHIdhyODj16vS2uAaP8JdFKH+ee4
MTPIqCPFDlC5aCnAW1Gjs9gc1ReNoIzyJVtMN5Wo2wZ9PT5mxEg6E9uGt/94+kNM8muDPVHoesVG
1YMsjOwJWh1dFTRbAo/c37h52cb5T2HFFO30ZaXkaLKduH0NYi3JPM5P7okHfefkYj3DhW6muVGy
Zs6R1wciObhv9BCoNUdxOfYlN0bKLG2hNZPxJAg7il6dbx5lYxKDlTXuzENrDF+Aa6vB5elzM2wl
rP6AleGAsnTTU/FuYPDPBaURM++FbEMaOoqcebrdichcZ6QdRmrpB4GVo/hqJa56o98mkVtgr78K
gkwJUAUBI7JGY9PQijr9fIHL8ER5gX1C8K+YW8TYOLyR+D/CqEYozL3mCoxyOLVEBF8iqFpOvbT8
nCIVRWUVuwv0bp1kGyVPZCKuS2isJ7RMlMohHevm/S9vbDqyTDJ6c2W+T6V1WzvbvH2aUCA98kMp
cAZ4OifEXYUWKKeFjwsLDUeYQLCWi8uHZcuuyqQajuWOf6tdzU8Jjp4GaUAKemYWdm9RLDiPGd9k
1Yuiajhfrc6nk/y+5yal0DAvep6GmpML8S4/J3LZBRK6Bkme03H40Sz1n91bre2ANTnzb9tGeyK0
QYPuooRJMEBIMkHX4/B707F/UfhNfQp/1ac4YYNvgWHRbFh1I9cBsnkMI4npDudREJ14aHQCqauz
V5LonLse+zufGZmH2K7zi45aERWl4es5nkCDTSYpysMJll7G7ziWqET3ld5FMUxRfFbtcYosmbBY
gi3pi5V9yxzhs8xMQPxhbmxJGYemP+mnMMk6XWfgPRcltf6PPMCDP4XEUtJTclFJZNcSJ+Oq8PcR
7YsA3TttHPNPqZfiPn+VdAu0yQfeMBN17886LdtISXvOMVUpyDhM4jHyoZJCb8yp62WbfpFo7ffI
UEw25VnSKbvg+lBVL3f9GLOZj/2/qzfQ8i/DGIlKI/PqHHITAtMIKJM3e59td5TTl5d4xNPVYL2V
YpRMteh6t1MaNERJbXRdN4hwpqtOb+nhDpt6TnGjWz/trkhW0IRYeDgXsG/6gHXSMyjhJZsdzfhS
+cFojfB2P5ToeWzq9I6mR6M6pO5f3NR2GeCDO1pjtR+C8GYn8Fs25XUNt0L9Yc+56W4tOranPhxC
cYNOAJ5lQhGiIg+Ka1Hapgu5mKTKGbBp6c3aY/HmsZb1TBHYBTonPIzyeDjSNAJvD09JmEO5IrjV
yLlOOrMXUd32e0xq+ihv+VAtqm5+pf9yFWtnfF573MvXNcQ2dsESDR1ncCaEQ3qBUG90VNiY7JYU
MYrC9iTr8SLEBEizoTAFmRqLxttZxYiyG1Ly/INPgUO6Vkdps98sf6lwSC8pFZHJtHfCUh8pme13
2SJxCdTs5+9QVpT1cHHrnrXkEk+SAOjTN1ZDiJCTYY+sdxrv1irli/24r2h1EkJUVhnxvnwyXrtJ
FMYJhGNyP7jX+MPQZZlryd9D/ujTDKWsjBG6lDUcX0oLRjeV6nwvnfdurStsy9lVSs2OuPyvy1Ss
6xRgji5FKrWLqAS7EKWrhQG5KwBdOFevbaxbn8gGw3QMxPosmxvM7ldLmJ+o9fIMc9TiDh5fy9OB
KVar4jtSKVwHfrzmRkSgNsjc73mkCA7gfghjOhrLnEBOkYdeU2Lfoio6YYUhQ7dfJENfxk8+zNuB
cvi0ADDF4FBUXeoYil//xExJJRqPjnUjIhiJzMsySfGu4e0WZAouPakOgcGxx+qsNHhpCbDRam8p
EtIz0fBFeoC0lO/8m95fadRaxkMLdwsPdGZZDM4U+4BbtKfPAPgUS2WsxYOk2d4oSqVhxnsiydLL
oi7ce5q7lpEb3wUqjF8NQwA5YZc4U+4S/qiiN4LiK7U5ZqfCGjsbZgYju8FDFrjfACcEaklwD/Sb
jyrG2T/kfqxVHm9RmdTf4niM2T38fMVj9W3/SBAhfy1BeyWUtxWlonDUmCZHyDeYPHdfQ2n+UBAe
c7CZi06J+sIFIkdPfxboMgE9Hf0aaQRL32UN3Uu23JtMltLgtImpBeCBFEHwvJ2DaCGmOl5jkn7J
ozq6x2xHn41T7Q1qD9PVwSpAVe4A5vNWog6iRmfRRJR7/w28ZXMYTsTL1ieh9I9XB3d/maOESdqN
HwDEpZZI8BZCAOIh3fwt6FnU9/4dTRqUKMKBeBeTSJMZNQFkGmCz7t0ssrSPTGw6R29sd0B7LnRs
wi5BdE7vhDNvYEI7KgecX/quYRLewWChlvQsHto6Rp2a7svrTSuo1zp+m08HptVDvE0cyLrnjAB+
iPS6FF79KhiVsX4eKQWuNykTCoyk8RUl6nsUUbWctqs53s2iR38JWQzdi/Ko5HCZr3Q6oGE0nkqH
ySRkmP5vaD9ui7+tKuPh0ZNDf/bIwitwhH8YjBvvtwxZnUVepmos9fzZG2VRwgXgPO4NvL8agpCl
oDR2E7iKkgmpsCYQG/XdR3og8K0sbrRV78VadB+mUUz+0qPLIToM+OTH1rzddV053lNjIL9mwrZ4
PI6LAxsElyveyrTHXiRYuiuT6IbG4pPFgV7c/NvzBFSZZ9i8gfAYhngqllJBfxH/ev7kZQmD6VGd
u/qpvUtPJ/l5GICYGAilb9OffH38JTb9dSVfIYmuaCacZUhmthAq6KcS0MWkqZo7SGg7XUaN08pI
ER7igjA+wL6BAKO6l9qEc8u3QT0BcsxX82424VsO6mGS12eer4D94hn7BvE+VXbVH/9U59fZiBDB
KFPazgPwtNg6Gf54skJm/O+GUGVGkPRn9ObNShtSJeXWVST7kKtu9Ha481Ug9+fDQHhsgHOYY1cc
765id2z81JvwN/pLGDuqLXqNfmnTkxEx4QcTb8yce2n/LoEnFBcBmEOYMa2tG8OEzMFJtIri2xAr
yDHFxb6OvumlqS68xU63m2WaIQM8wz19PatGCf8a+U9MsaugQ7NCJPXYrFt73FWAkqhzUjTo2KDe
rJaI5+6gSybO9kGTUJIarD9+n1C9oTrzXcSqQ4ygMvy6QTacYA9XTIQ74QAWdJOOa6/q78bAwzGq
RMoKiBYY19U41d62uaBPoOMdciaRBZGjA54hMZ0HkP9DnstsI/1Ly5cFaIdu3zWrCtfpe4qZk19I
WLAahEpuoP2vTcRXXi0usVqUIQWcslQmMvksegmLATk19tu+uAfe+9TmGcl6/jU0UkX+XXRw+kaN
oInjDBLeSJDqJ7EJNmxk8UT0cxvi2AXRAwaNEy0C407thu94gK1TkKzcOT52FWFgU0LXpyF4JMq+
x1QdBb1mt4E3WrxIS+pv6QsKqvoJE4u+Tag9WggaEcARasflHnPff3rjm9j+YzRYgnt7q6UFyibz
PwbPWAziy+sLsksHlFpTizVclCJlLPTVn8vTlrtifWex4XalJ9+5lMCyi+Falc22REyCSRmgDJJp
oZXsEGthfCVOx7c+qcvod5lRIw+qHuag6SHlHuPsMV0q1wcxvj//YibpmLbRinTuMnclPLXnbkqx
PnvKR+0iD7Em0G1tgKthfC1d84BFybLJRC4CvUNQYA38MeAnXrKpTrKjq5c1c1lsq9vdCOvUNjjp
XsccC6IBvblaOCIGZI9huLOyHnkzc5u26Fn0uBiCiVs+xV+s7DXXxEuJK9tQSzXWKR5dyK45kUQm
hN+GaFVCFhTl7hKhDCNhnKX39Lb9A3vzVpjwhcxm8f/8SOh1If3LWhsx8ya9vxodR9tilGGBz2R6
mBU3pWIlZzBB00doBXSugk2srsBZgY0bVuCHybLRy8Jyb2AEpVN8UyDGc7ot7ZnX9AcsJlST0dqR
b/Enr7SlRSpRT1d5vCyBl6vsoWCJSGvuTFL/ii3FrDYPW0Zz+vSCmz/uGsxWln6FvFAjQuTjmv21
D5svolUv3MOW3GzgzmInRlEmannTspGGzAJZbOu96b5bI8AdbRA+92jvsTRfsqhG9+QunWbpDLOy
Cd5ZQczStKMBaQbxXTLNYSMk1HBGKhl4qOJpL2KSwAfljbg41QF4ig6wUuEMvhAGKFZSY/lzpe7/
F0Vp92lLsZ9D8E6x/AfiDMy5FyyU7KpBhdrbnbDt7XDTd7kDvm6mUnyiWbnvJGY3iz0kJA4rPETt
7QINPY8J8nDPh9ColkuGqW0QXwVc2iaWz+WlKahChCJ1dPHHDl7lVMZO1z1s4lTw38Dts5IdfGVf
IaqFijQIZJ8iS9g5WagPv+5uqgyj2EubawOIAQ++aVyFZ0ppRjzKkuGl9aB1HsIgiNRqLqAzj2US
iyeTr8/6847MSr7la7k58tvodp1k+ch9IoO0/i1vucDUqkBQDxNxLMmzB3WW4lZ3EO8OpNOH8jN4
DnJ5IEN9fUoWyA7OPFAtHtxMzCT74d50jE2XkNTcjNGHI5y9gkwCRgiDPCnEIVua5NfAR/X4xMyM
0UkM7PY/Mvej1l25PyijyXB5iC1oOph1DrHye7os5cqnMUlQiZCVkk570r/SLjE5iQjKBRHkQ52N
u5mm6xPpOht7GCpVQv4KfyjE88IkUjnUk1oqf8snzF1ujq3kTIwFKRA1XWLgR1qtuh7x58K1wfNW
dhfqPkkJurHAwdQaZvV0OMMZw3K94UTP/W/TauZXGntojcv0z3ExzQZyJOHLmCAnRif4VhTuitv6
kNTVFLKm5f497qxLo2vo6Lgxwl3fjkAll4NlzGeRxMM97s2GokyIJ40xNs9xCt9/chwv5vmYp/LO
z58bCuZhlRgHAUCDuUx0Cs23rJNLwUEpmM687b9mevdnZk7rGINA4pHnab9JvSm162MdxO8Rs5x6
9fynq5UD3d0xnYoESE08ewov41P0uuHuwFEqSDz+BhwE8esQeLar0wvhLIuNSrcCKPMooS6mzIUE
QKsP+fbdgIgC0JFFMfnam+yjTTJDWH5yRmEfQLCiQ57NI8A7xIfflgo1tQDbhmJNZHWpeksld3ED
w1TbRtKMfJR/16GVhpvaRCTTWS95GRsp06I5ZAGNdqpvlyAY194ytHkKPyDLgenr2Sg9PG/RQej1
hiaARoCywmd45mxQm1/JyBxgAeKXZLrQQPaixGxOUUJz7bc6wWLoSz6ImWk1m9+sJDCFNxqxdCsN
I1Dhk4L7CMqFbM11lSTDZQeS4bOllNseO0ROGdFGZpMoSbtiOCiSSz4pOemK5bl0k3D7zBtswV2d
ZMMYMj+QPR7+RX7sK/bDKAcRug/DwAh2vcOMjxKndCF8J2KC8tIaGP1y334oW+wvYS6R5SiEUCNA
WMRreUXK4ZnlT7lj1/GpVfD25p4ySbP+xEjLxqjzsb+rNCfxmBwZECRogObravLeQD1ZMnbB5ILw
7rX4PKI3wBrXLC+pFZnVsWfCt6vlam4+iq3CZun65BouDziIpdlmC/ikjJLq1P6XyD8JnCvnSLCO
6Lmu2T/YpRC+YBz6TVGydSHXU1jYy33aNt8kS9v0ZOeYpeuJZLp5Y8XvsenOLJTOwOIDfacn7sWS
wX9l9kkKL419o0/IGQQOYsUQnzioIYoB8eKcOHoGvJXCo/P9DKyYQ2On6b1j+K9vkVU4b4pHenPm
GT3XmY4AfYgNH438TdRrYGaG4vuUWcZT+x59y2kykIeemgbIpRk34/pL8+G23h7OlyuCF+WX+4dQ
LKmeQon+SFJwf+d0Cc8DrYf6nbWoEWAuZs0sv0At4mI2vMh4nQkQ23xQGDv7wPTITcd6CEtyfA1/
W/+PJby/0LXo1upaMU7fecJ4vPm2zaIyyQxewJCaB6+9DH1xqf9F5ji9OlyO4jgsdtXe0MOsVzad
u+/O7eH50y6NnkOrEhDEzzILoa6zjRNeKjzIw/U/TTm8RfJ/LC59LfoiIkHnyYePKljakCEzLulf
ug8uf86gtlSmbn4mZwkUn9haKnOE1pPIfGMArfr2Mgt7bBbleYGKqG+IuLWkZJS+uf+BEUGXVOMr
aQkCNFnduknOF9mInbeSevE10QKt9FLNsfDJkYWac+tCCysHA4nSCAAgd1peF8lOlvO8CLKprZ9j
/U06etKTWyiVlIud+sdc9/8NgLH1PdU78iFruKLQ4aeblCO16swxQwqhNQfuAE+moonC7rUmY6Wi
7+WtWrpKEG9xkZOsg4IbMwFw/6hUqn57jgPr7NF/6QajNvg/lYZ0zl/uEoulDS3tfWOpN6T8ZowC
c0I0Qit7TKtcs94+schcIS/1c3Aaf1/MvDkH4+MdqGzMa6YJVMbGFRYI5KKrnmI90/o42YPBtVdU
1VecOzjoaNKaOvTPqSVYDP4eZaPVYATOIjZRduZ9VE5EqB9StsrNwsYnwbfSw6DVXFpRJNqdaqNe
ZObkXkG6L63D5GiqHh2+s04OB6us0wXnmEMbAhj+G/w/XDWVTJ3KsuAZsAiI72r6nBtvLiDo/QE4
nIPYzjI+hy9WSStAlpY0iZpa7ZyvzPR+Ru2ci+loHR7RjSTIpOHaWTp9B4rV+2qw/LddPlDQiSfA
Hrm1IaDWnq7u9J5EfoKoLOZIj5aWLPkAQx7U/MQNx+h/KBD7UyBMa1TUkFNESgwpbjYCeRLn1zfa
kCnHzrU+l/Wi/BNYazOmzB+hqLxzyhcJTNsLpap4MxJnnTqI6itxsoNJLTSA5pLrkYP2f2GTIUBM
aFDhufuO9p6afZPR8kvEFBF2eJszvGPSVxN5vfxbXiYr6T9P3Bdy1eaRQlhQSeeLaHKnXDnEIzm0
JUyt5uvuuSQSebkU/+3eHW6T0RCs3tF5TcVft7n3VqwthCWmjjsOjbtGjgXW8W3+Ojm+QE7ZFB9L
SjZfzGM01jB23JewmhRIAXU5cJqul5J5CCanh7A/04Vehke2BgB1AwDIsJ338OhCw21qIsKhVt0W
soNjQgIMWocNhaji8ULoMM7c0d/m8bpm4UdqSY7rVhuENlSh2CyiI5CVILnpdx8wo5vh0omFHmnS
Z8C0v2vraxQa/VpYm9Rd/mtv9YWb30da4m5nSrfBLxR2jTmzuVZU+j9RIlhjgt6AkJ1g5r02urdy
q3crNTydGlW8x2Itzdp44l6zbSM0SV77EovSwIRhL1cRtcbor+M3V+ijLGG5kKi21fdWZvwEJDx/
tAngsgM8G7G7OztDBj8ChBpUphftn8mxJCCiHBu/yzF0Il0PZJzNHTY5YouSTVYSgqAmIOqf/d6d
Q425tdRxZmvilEo5xXmczRqmeUOxN8rVIeuXMkeWfulZII1n0UGc6TgiIIMjSAkATHU6SD82xYve
L+tXIbwlAYZ/uOQAd2R8QvYEZmikTEc20vRaF03tgYaVIZ20+JNFAx9iBYoCPj98Zlt0WCYEZXbp
TRrECrm7j1HUMvGWIMLBLJAs+bsv1TaK+uK3f3gOOtA3aiVbTb1lF87eSQBMa8c/99fuEzMFdlX9
k4VK4VscckopnkQzwIAwQStNtFD5pQrxJDHaJHpdYwKG+Uy2HtuiMiJ6c8anAJFR6aKd1GeYAbHD
0Q3+yFq0mt9MSFk5lOrVYedZKwKtzmh2fGQCH2pkT4HAElzB8qVjg5q3sZ0ALJW83NMDOBR59hfG
VdNasQid+W7n4fUad8uw9tuikaVyDcIyzxnODx1V6a1tr+k3BT36j33QnwRjpYGPi/3iDbxGmfXW
LsqV5aBN3mH40hr/Q4EJjLaJDGhg+jzvc+E1sPKNqn2dm9MlyFdA55d/d2Aeklr60sqqYpfHBJti
X4U9noCh1quiVCMAsFfmys1kwrcIgb/sZYrBbbVFiXX/q3hMMa5KOfLp9XEArv4fMbc3T0cjRbKY
M014DOy1syL+yf7JqRwk+8Csmnl62S7NiEBQrtKuyu7jtrINuiGXY4StWh7lQ/1y9NPbmF8oWa4w
0ce5tGQiiQzBQlDURB53PtY9imtKKeaccjFz0f016CMEa8ceH2TzPCIBNIyp+IdSxwiuAD1+nmki
Htwp0cbKxooiL4e/4wc0CuBTtghurokAdsVGI1BEhojwKtQnpDdfI4vxcA4DO36jWkYXPX50+PwK
6fnsB+FwyP1Jns96yLDdgWy1Y8R5bKQVc277GMeatKx8mC9F4l9fsDsXyZE8XWLqfWprDnFz0qRT
WLncnMBTcPYFDi0v6So3QW/DeQj5LMP4gRvIqYvI+ehaKvWmd31/Pb5btt2Pl/LqPoXBz4UikJ9Q
anQqb1dN1pdH+lT66+KNyF3j5EoN+rZ5hhkjcjnkNzUkgAsHyzuirOBKl2Ou8bL0sU4N3XQA0a2y
QmRAVPxYytEpoIdrl8Wo0gyzaNrdIc6utBzCHozJRGGuZX6vu5/yuiyW56B0ffIWBd6enMjjFTSi
PLSMQuaRcNvOu6Xc8yUinnJ3JiFYgwCBfgHyp+vEPf7A0015Fw3OXFN7yWsjiBIJnoUyX7AiC/DQ
kP+JDPpO0Iuzs+cHaYVn0CuYOepI/XG+jE6ehJ9lZJLsv/5s6uBOP1Xws+0284j2KGZ51aeoOWfm
GO25dQWL9tYXLFSDptfswI7dR5Eqq1/RV7MJNg48WKJImZHNTHvMlh78vtDox2HH5u1oJbvHqNre
6nQJ135+X1zCPVFGe7oXlRtxTvjksItK2AIlUCCZd5rmJQnC87vvoXeni6tkS0nxR8C4RVOhNV+Y
tZk5tygdBDdVIb/eFuZAcxfRXZXRl6JBUB01zH6yGKMuM0KAE9AKZmzbGp8v802qns7QSImsA2Hg
/ASAPFD0Ssbb+7p8ipV6RBPu9pnKK5XcX8CqjC1Ilczb5JoGISI/LE23b9eQiFerJCpzkPgGwiuv
AbORWzLS6S7t4X4B+CR3tZQ12g5SY4ZbYH+HfGKWv3YFSRrC+6VNPgfbEaZZqBq53nL8hbRS2U8u
sz1J0yk1e8nA/PvQ7DvNTMfH1X7ocm/win25V7YUoWvuXcIXEaqPQF+YB7YbyjVrrK/jCKsqxKfC
cLzo8l6M+JAxUzlb6GLQiU29zG6i69fzZQgmISEPE83so2zfVfNv8GdKw8Gdee3O/XWzhMNlwBEo
mhBZarznf2PoEByeafowFJ5129W8TNogpQIooU6xpn9v29/M4vVRZ1nbtInumc0FTJ6ItzX5Bytt
RamF5ojLBA7MQru88P/H/pnrJtVsbXSwF5Oh8G3v66YF3PJinCw7N7WwY/UmlFeyXI1sj+6VGCMQ
nCcDAie7+QFdGlksev3ZasaSm4uOr/AlXiuuHmwn/rdwKIODLREPG050cmj8LDQeNPzC0zEhTWxG
Nd+By5hnQ9fFmzr8Mu1vodhxG2LVcAZDfGCVFUOS6ceqKh5c9MCNHQSJ9gFXSxcEOUIOcT3h6k1D
0kxPf45IcEi1SrrQvj21cvQeRpgeeUj4rjGmrn6dWfJhWoaJFK8Eg4hWnYRf3MivvaNqbdf3VsFr
ho+UuMkP+CZn1I6wMvslRL92gTedFxW+o3+/j88zrIC7a6kWxwxJJuMfXS/7/lpPSGQrZ/TxcnyF
2WpYjxnERIxTG0TSufHYw0wV3fJxqDiR/Nw4t1egkTKulSas2x1W1ViZvV2vK4NP7oimlmrQiqUY
X7qzG/QQxmxCW4P0dxOjrsl2TYjJrj6wAgKH5daVZJY0Dpze0CUSvY9kuqMrODIpyg5J5Wd6xdKo
FHR9S+AfDR64fyCDCEC5C1ObzcvH6xN59bvI8ilyxjf57dlJEvrBdzjnJ5stcS1dQh2hig9wTm0z
aQK8lAwQ0WlaEgLGA9OPQ/YXeLo+14kHFtXPHxkM6pDV5ySQ+eMQSaCssdSOqdJzqpbuXBMtdmzx
Qtt1vrBj1DfejSxtHhZpSsVSCDaIed67M3j5aKds034tBPd/8FaY+ln6IahDhSO4VqkBiPiU3p/K
P68AJMRGtVKFw+BGUBN8YgO2iGlfYQyTJdWHjJZmGD5ROujCxKyg0hWHNHuLG5J+XL8kvVvOipu1
7FVES0QLFyV5mD5IlHyCM07jHgzhlquU27HG7833OKKLeOg8no4ZQIM98cFCzHO7bcztFblCCYuw
0u264Esem2qO011COW6L0fdj58oEs2HczmQiDZiSFollNrRZGBmVmqJqeAX+xZaHV/SCN8gfh6Pg
77KBr1OlPYDpyid+vnWzNR3OWqyRUrtkJvmLDiq0zBo/hJoDZJKgJGjmdgyBt+3+Ce0qjBTe8YgZ
9G5HPlnQ1K0D+MB6lpQqdYLiwhnJ34qXP12sz4NQS8EG1eW5jMnQ+Ixtr5DbDel3Ah5t94IjBQ9L
un+qLG4Feb98MNcJUvOv3FArQMxULVt1kyEmRE83Sy8Bh79yoBNO/jdXBiGtEtt3nMPK9D4TZjBG
Tuksv8Cucn6Awvpk0iU166OEwoEwDTwloCYA5irMKlW9U73Qr91z728RI+ycUy0YNNJP1OPVg9rP
r9hoAwq50TuckxOie56Q+I5J5KhPEvaVZxIGr6k/IjpUU+jf+V55VDHvBc32yU6PcFfxTxsW7wsb
JzCKy72TUqLIZrM7V+iEOMGqTY7qLy8Brvl5kHMqAf0WdvFv9nCucmxVWMW+bvE45hZakYuHr5+z
dP4KqysRQU8HJhggiEbhRdlDy+v0brIdS+39/kFfaGQvfW9rg50P1ZiXNtb5PM34DCe743inC/SY
M2h8+MI6LEDe/B80mEgJ1PmHY9Zm7k6KvTG66nYiD1R6x/6CE+IqeOf22uLVBmaZ/06BAKqSb42X
NcEna4ozMPWcUK/WFO2EJKhtkfqJ6GfUk8kv3OspTM7OB+xm2FE4XylICq6+GOLm2sVwVQdJkwZ6
2v1x5BaQZpdHzKQnzvXhISdnw9lFhxL3EVKqOXnlAQmHrQw/Q3uIAMVxmx22f6KtSGJ9CnRRtrNx
5XRDi6p/HOpKIFNpf2gPjZdyTpW4v3Wt81D4C1lmkf7pOSNVHQQixWlOdKg1Jyh2mooOKaF7qPlO
PE2tuzqLzQqLqwrX3f20drpRGL+ni8gZ3QPGiC7FUIjcyWUoms0GWErSCy/3fIq356SnD7ykb/+y
dnPjeFidrxeYt7BGKbcp7WhcozetO1q14n8lM5NhVRakauVj/wpFNHjn12lul3m4sBAPgsRamuAn
DI8GzpZqxCQ1Jl4E3MLauBprjCFMxaADcQQRqkNAQN9m8Kfdl7v9RoFUxRkuaI+C8fN9qMj8hyMv
GNbeKm9Fkooee9E99lN7NwCWQuinEc1UwoQnM92ncLIw5+y83DMxqRbHf16HkV3aTbc4rAY7BruT
9N4Hs1oJnrpfTkxv5aRfI1bJar+E5NMM5qREtgE5qao++YrQFHoajq4WKTNvLr3F1740BU2b/E6z
i+6RCHYnHIBrIN7nLEPQ0dwESSy2hauEyjnPypYz1XZkXAl3t3ldVg9x3kCVpwotsfKEuYrjRM6I
9OsF8naCNl2qeKPub9Xj5pX1kGJXsjeHYX5oL9CEoguGkFOeTFTe/bNm/IEKcHF4tSyujYfCsIR8
5I74aSK1PBCfVCjNsIL2q03KfpsFdM8neBKUy++P5vUNuKOUYAbirh0ucdtD8nxLJcEc8sQDaVFe
6iaKeaer/jpz7mNa/WcJ8DNN8uyCfS9LqSqkfqUn09ck87cvGa/JwAtOcsapKwGUcz/p70hrQweA
S094KTBfMgaLLarriM17j+hodxU1k9GizJIPgfEQ7R8oQ4X77SILW9+4Gnv854/7ooNHSNuDX3CD
YcI1WIZpyaOqOYcr4FpNQTTupph4wZouN8cY2EtlnReX92nAFIRAMzXMmqvtBWoqCQOsTfOCGu+h
aUaKfPQigiJsG4I3KXYyN7B0bg2fA1gWNgodaEKbOriTjwON6zdiLuNUKFBUR3NUeBx43Y2bflBV
PttmphH1U66PO3E4ActoShfNlKuwM+mKNHsS1Jqxex6at9FAj4K005VGM/jbU4ObMHB4SYYsdsqN
AGTs0qDKSlzNwnz+oE2gYtnnZMQPu85RFrKSXd4sqPMg595Tvz6HgqYS/+Ek+j1z64qga8rb1ZE4
zgk486tFIcerFTeMkeBtkSKZ8Rn1zE3edKyeqbQgnjN7eER0IljrVLUh5UMGJfvsXGc/BYhCktqc
OJreRksZ625b7LzAa6a0aMXMMiJY/FcJ0MMYh1Vf3e9bpnORyxReMQNvdTNnO48DpdFE2hEX3L6A
cBS6q6ZVRqGQSGOmXW19EZA3L9qf3LxwxsJDNWmhCyIbI1+nDsy8b3rWZHhX/Xiw4/iAsnNcckbD
+ytt0kz1OdD72IKOyXhNa0RjPthaf6Gppk/cr0gT/xasNAXhq9W7t6hK2kxrH6DGXt2tgnv5VWxJ
XygIYqCdnx8AgMzPvSsAEW+ibAM+auunMA+QSvLaFjhvglf/7QJaAOCiplq+JMDUszbHV/mlevSs
bQ//zV9M1Nwfzvgv8uJlS3Yb7/Ig2mYHiX3L18V5fiMYPAoR6mLhL/CO1D+6jHmQkpJOSrs3LEQD
R3wKRNbj2raohH1eKc2iKtunj8bowIwdCComF4gllBNLEoz5Aga+mvA6nZLNZeYCbeBR0geyJeFn
nTpDLd4pd/axeAqmEXcbd6D7Mt3PanBBmVA4rD6uY1ruaOmv3yDPfyi157MLhjVleu05yh+t7+fy
PmwpwIqbDhiJ+jpDz60Q8A5EjN7JuO1F6f+aLm5I46IH2YD7VzlU0XMpv1vD+nNfNHr7Iq0Du93S
NnBIKSC+bycf18Kbkm0QPFNAWfGwNC5P5KZwDujNqIDekYYFnH1HBcETmJCCh5W5K1EfS3noCsfN
se8cL48YLKHho+1XrQk6EbtoHPAm7W3DOghVwvMEmc1ctgseWvmvgwwUPcR+zHaVRFGv8v6hXckW
ko4u2JMyVp5jAaP6nyQxH1AGGLx24BPdkYBaEjPAw0FhK9iTtfv4XpSwouSd4Qs1a/aB+Ynyvchm
QpkvesiM3EbJXam6dfG+X3v9M1FwomBcK2AifTPAtm7blRGTxiDhuLnrP/2m7tYsAtHB10YI5Bjq
bVRs6pQjgZ/mqp5VwshzDM1JS0h3iIrXo/A3OhFFE7UuJ5/vMnAOmh9PFS5LI1Knz+fdo+qj67Lz
zvepHW5VhCQJrLbj3OEPEcagCZ8wiJv3QCtAxL91xgLzRKevQrMOSRz4dN+uxMm7kpSBRoU4QYMo
QrKY5mmZoOCATBhtjks5f5AZ9sa9Xpo6Hh2TydB++K7JTT87d5ij2L+DyPN3N0FgRITrQsJAvNsX
YjLL8j2tp47TFEMse4mBk9ag5fIJ0eaO86MltjLqStl2gNPofAEAaDE/KiTHiHOCpLaDrpwxgiz2
iL37IKsaAzpMI9l4plxB1WcJpw3vxzzGfnHJ0d9EGeAwmTWLpFSHr4f+0KCczROQdGNIqygrpg5m
qN05yJX6qhnX3eXkcMIoL9VMTW7FEKWiWhMSRDCN1ze6MeRubcx64xYqWnrIphJ6JwkKI4WETvAG
kXgse1zpTamHdZ2r1YqjmCpbZnJ3n/uF6c/EhmpRZCfFdtwVFQmsRVyZ1VGwa0DRwno/bkggmPqD
+7KHo2bb/Z+YbNPMuYQltIeKz12Aqa7D9mKjOzqIG6b1zoudMOfAH+/8OqyqTL34vCwnI1WBoZUt
veHUp+zrmx0r9wibaInXYX6T6JUUjZOz1ydZ1ktqgd+NkkXjA0chXBNpXaoqTKLyKI12CZqcHbFN
jrDwivQT4ALmWurgJ7C9b9Z5mzqNbsfpTzZirm5E77FFZGn882r+5RWFEo1rZUDRgK0RaJdxUYTj
mAlX6Sn6WTA9y+GVGuxTadpBTRgV+ejgz5hEUHF0uu9ecr85Fx2oi1EH2Ijwe0cM8BPUymt7JMxy
C3A4ARggoeOqUNEde66KU/dn5BMHUIdTLQBkPHOzmtFmib/jyoJVy2NM9T6VyMSZQmQ5dFlKscvr
0NEvSAEPa3Dy6NR+lcRmT35rYpzOUx82uG6Rdpkmt280uXjwp1MI8nog+kMmChT9lRNeFKJeCafd
tIaY73QP2dZOAor8rkzDlk7UPA1dv4WUI75HiJqLvCdPFaUosDAn4KWpiwCHxBH0CsGffT6czE0e
mNucSJNEb/gwJQXBCYlYV+bUw3HFr+EmANNscRix6YQwPfjXPwLM5ChyrhIeBMDHCEZyHjPLzTmU
5G+BVyPQVPYaAX3SCrlnZXzxdUajRfLQiBFWOA6PwiPf8zcLXzjEww8FM/1ODjzIutW8TnMLXtQG
JaDWLF5/OErGlyCDM8U+fJKN4mijKKfzIpPHHCo6lCI7KegzUJblO22KJncImsVFZNNhnwPN5/qo
bMxnFfxMXbBHtJ0icQX2I464MCEoQwcicnG/TrCP/kgTTLkuQ2Xii6v1kVfJLZHaEEne8HHCJO9K
KZTSp//O8Rg6+QWR9GpyC3RiYZt5+KHTPGly0VzZZanuQvG4Vi3cWE8gotpDPfxZ5x4pkVkRQC0a
k2b2yrAEa5Wk35ZoJaAlphVAJtjalmpW/zO488HZrzFcLPjRuz3pNLqdDHtFo2yBJK02S473FDPt
ThJtcgp1paZ1/ZR0PpvkSiN1konlCJBMaNVKM8kMAXDowAWjkV+lFxe7V6WBxr50HkOgVje3XkJP
XGPP6wqfUfQpXOnGL0vrAvfWL9WdN59MTxQxcOHZsuG/0xONbfPkS7qqCWj0TLcUDwhSKsyV1NyW
nHD/QneBoE85PvtKE6zjYhqucqk/3AYsGYPXvoqgpwJ7Qb8D2S5bAgwDSzfklcfuFrhRC24bSae2
RVYvhwsoiJlNKl81OPcLGJTOGawWZKUX1UNPsdmfXNNH6+n0PQtHUV6bw1DoswVjqmfRJZl4wWRe
yuXGZBYqGmMzsa3vgaAG9nWdD6Skad5im2PVrUUlOSPcw5IYA63Z2X+S5YGKnMEl+fK3ZTVaG8Y2
daSKu8TUBb4fEn4Djo4L2OJsDLB9FV/RBR1EH/JO04vv4cdXtOJ9qXZva8dhOFuDJLrwEQdRLQlx
wWXepiviXrwxQ5ck27okKJRcU/+KTK55S1RnFgBXFXhQAu0HnA/Wq8+ZjAP9asrcuVW3caneSaEM
tMu24qj1T7TyL+DHaUQtXg8p8p3aChoV0X/axA3iq8Bq2zYgnsutGCqFRI4LUBes7iqOgCcr2nO9
RKa+0uAIqWkPq4TIwq5ggaqgybXsLg+OZyrpG+6TTWYrGYXalOjpXXBUta7sTOv78ZWtMB7TgAP5
KMM+6Kxe7EWL1o1HcCfhOkSD+zq9dQc7EcjbvS306G1ovPcWikGofl0JSSi4i3CgxcxwPz8fCYPx
tdnMT0hfQ9ijQVCum2kFOMy2/wYFzhcBJYdt30QSdHpUO0GO8U9Rx35IIM9wy297F+YmBBmNGr+A
gtWbNPrQM5VO3tFRIz2HlBNKGozwdJtipj4ts02/QAS7dJ6v8vFS3B1fXH5PLvZryOOhGCDdCQvi
QvEocl/JFMBXeb65vHFCvi2jRWaGJXJ4hyGYQzvBEhu58VlBVYahF9x4yGRNr7aboqqxE4RHFHyO
f7tiHj9GANlQ2JrHOMV+052lHhhPhwqdyM5+1GwPLB0vWvXC5HAnxMJLzCkaH4dK8PVbc7cQ+CPh
D+Z3caTuqnVORfCcff2NkUAq2GFwUAc9SXPPIknXGTyVCIIWlBnVzLyEnL/zUZv/9aJB7zb9VZbs
0aawmiksRkViunJfA5AUHqDJRKOFj2nVgqUjj6bdlVuFF7OqCff1QEt8Y17q4oyQ0vFTfp5rbBua
gZYGTQQBLlQzm+c8eIpOpj+pgvAzTymVqzXjwf6vsf1hrTDg77CWM8basTr98t01uu6RGsmrd7M6
jgUdwJ44aTYtUGhaw6BTPl4qGwoFOrw8KQlxhTEPCjkv0p+juBzxwSe8oNL0ahXPZ9NK2d2aYDkd
1Rj/Iw9bv77yWrP9upGClPQR7ynLojg38ZJKgjFzdARXhs5gFDQEuC/CiHBsv/4IA9Di8za7ZP6N
JeowhFhdas25EW0rkc1ih6fhcVc83r7GaNRHTQD/3iLJ+K5xloNi1ccRkYbNvh4rRoJ658TkNmww
mrumjkvu8KiNe1bHcli+OG1BzqzP1WfBSMUtH/kZi/jjZ/us3n6pPe5gonr+20j+d0lVLimWuHer
S0yOIF0PGcReDlJSR1w8aOdm+VOovHq8LWOAAc8DFhypGDx1vOPXyw5YXi3eUKTKfODPzcddnhf1
y/e8ckkiMOvm4Pf8P7DD4CgKMXyxpkcMQBKn98Q7nKN3TT1vgq+QqZFaH33+mqAW/s/YasmH7+GX
eB4rvCurY+p5i2UKfu0YJFybDrWE44UsIqnGBLjg/JHWnuXH9rwQiHaks2XDIw/CIKTv9E3ZvND0
g2Rmi+epmg5yfJ4TOOm8QI67iyOo0qJGiPLnYZSn8j1h/vwFhsDHQoEKzCMzP8SV4IIT4K0Ax7OU
BBoZpb4QP0y7RLB9uxgszkvb1L1QwPftM4mS+TAoq+VkU8z+VHA27FnUGuw2s1wwPTnIL3oivhlv
G0/yk1LG4zxqIGF4gdDNL/Moo+q1luHwVQzrxOvq5FvsN4tEdhi6oM9QbjOxOwL/4JZL5qUrfEKc
/AJBWM/Yeqzgw+Sfji/PHEX/k8A2YuU/C4FYe4OSaRzyxojl1lgfn/cdjJUlw7lK7//gcabKUSgG
jE2aymuC4yihXl9BZofgMzSk4308zkPP3GmHksenzq5l/QSSp6xPmYYBWCkSPuJTDCRwXWzhX3tE
CW95v+Bk9/mKmhl5tnYPkpaFC6tzoLq1omzcfazJHcVRIsSK3V2wdrBJYMwsa0d9tBsT//T2CtQo
InbftENSDSqHTR4sZUdVQiSO4C/xe/1d3Q8/dp0h1ygJUasF9ozkhniUWdgZ4P9H/fTNg3pfpFv7
M2ZqCpb9uiKsmBbYUowMuStYZ3LMlNhzktjtGG66Lpdjp05qjTbJ1OaLlnUVm2MBoQB56AJxJ3qb
u6aXKvVx37/nHhWHu8Cz2pX+Tugqe571XEx9gyKxoXJdjEoaEYZv/cXzplUlFWVI0ZeZPJEsM32P
NX05rdSJuGcAzKqjz7wPPOMcSlXv8AasWAvB0Z8cRi8hwOM3oL31Yp5oTyloLeWajrz9i5CIiNBk
pcqFEITTONvsIreyb5qMGFj1Nz/5FWAvf9HRNNGG9qXVUi3dSVuDawcSkT/W3UlzLYZr1LdKf2dA
ZBCqScdupoyx6wibKSzxkH1odDJPPaUUrL7uJvtXJft9n3jY5NvIaxYcRu8d0qvytqtEK6y6pQJK
FCKrdbjLjXaRjrU3XanBKVSFTo9DKyrU4yBlyLso/2VnL/WGLWzhMJbXRRhgEph6hHoaclYZ/qjT
ZxWDiHWVLrkJ7Ifs1wc/ooFGY3sN/7geKi4VVwGZjG/WYVOF06YIQOrTakI5qrHbklLyc42zP1wu
uwV/dh9zMGB/apWljqJGNvxkxYA1JbpEfM1p3BgjAtrP71oOUWcQYXKADj20iNumWFcNwfjjsBTM
aOcJ8wJno+kff2XqWSguliN1WWSfbrzjoQa+I6lRQ8ysCKKTBjbQ1h4TWlwcxN3GPyRzWAPAHuA2
1ZVqwoN3E2G8rJfVJVLCy0nYFmiH0x3hTd1Zi0NnIaAs1PW1oBKoGlTeUNlT9n7UXbQV8jehvUco
fU1mtPNVIJWSDXR/R2s7btO77v+DUWA2NpyNNvcaD6vjDHcfHtTmj+rKGALZkjgort3iitXK+js+
pFGAMzZsCBaSsdmPFB3QYEcrbYGtXm0LLPAgFGo15VW6cn3k2odt3TkdPdq/MKZ0sAWon8SnUA1P
8jMLf/kpGb5PdV0Ieq68eu8lYxFNlMGciQ0cgdsaFjY3JFv7MmArgWuvJ65LXUZzAajH1Exq2kUa
QhL9dpN5OwU8b4FS1atuouH3h6RWa4o17q5ZIMgrSH2JMrc6qFX5uJaxVRL7Xcdh6E6ZyFb0ip/7
nC0esuWkUIuOUQTG7c6d4UwdObcyAmjttTA8t7kIyX/InsE7Sot81r2qNiHmOOSbfhOwXRDOmgxI
1lXVDH15h32tgIj4Xg8p6ti3u+Zjg9Qy5UCx/zETwz0d9Tdf3B14tPwi7UedpYGeQpy2qz2eGWuJ
n24l7OR8I/IS3bBIkFRzY3hL40j9/VhQTYReO8Gf/yxbPEbU7pOwEXMLxOOGulZR6fZiVkMaJ4GY
j9VuAsH0yUFiOZ1roFux1CfxodEGdvv1WbdAkcYXWAkzFmxz5v770wc7pUwJPc9S048UqlCtASqM
is3SySRR1DE/4A8IMtAg8OulAn3JTPYQOqQgbhq0pdr3+xpiICpdE1SA6vWbhWbDbp3fRG16260i
LF0vwW8dJ3xK81vZ7QbcQgs91ukqYs+rOgV/Uboj3KWst0uA48p7Uef08GL77lWjNpdmF6fCC038
1GiWN4ZYKFnWZ1HRRt5zaa75PEuIZXzEKWP+fYk8Y41Z6twPBwJ2sfWQEgAqfSyIjYsLpes02jXq
NMi9bKD51x3CdrkDsUioVbSKTNUxbIkRey9pdaNBGoAeaxB5qxSqamJ36ljU2V94IyJ8R5tWHRuN
mbSRqLl97Cvi7ElweCswx5XF1WUqlrt/MmlEI/KtzC5O2mqOUI9OzPcRSfkf1avAqLq5qzZbIodo
qILqboaX86DGwAPtkprZpKoRoAgI8VJE/aELiodky5FQXk0MHRD29zvIy5NX2ByK6wMkOPP17Yi0
fQuFGosM+rMsmtGvtSSCg0gAO/h8H8Pjbc15qNTMzadWq13Ctxox2A+XdU11N98OEqAM0HmokmSD
Tced8E/4ayX0Qpl38YLgf9udFIwDmH/ATIPnxWwll97jN/dUhak9FaGyptoEQhPRbr0v9SNrtkQw
ytVJJYxxYqtlQ2TgZ6BBPqjyp+nBxcgW9DKlgUcNxEO4nBW9RumuN41fPN70ZDKcn88WNLAC4DcI
C1aocmgh98r7QunwvinYXL9a4605sTVRoYkvFUD+sVGMzCzwTbsp3mTHX/6WO7iW544x8Xa/OzS3
nViY/ODd/K7YaVspHyXYJmCnSwVcPEzfOkz5AY2gUbRY7X0BmMeDXEXmqy3FanlXVnmJPcOTS82I
WFsLF1/uoopGs8Sj+7UBb+4ggM60HMAbR3a7S0QijgtmnAFDPVpV2SfMI0GQY9cKj2/kSMRbhNNw
C2+9AakWG2TFHjcqvF2B1HvczH36qeJjUJZEgoTirznz5kHmUHfOWZ8QBL3Z7MBQkB+LPWDVSiEj
ZQNaQFaBdz6tPy1X1V+zh6eG4UqyLh7qizyiAmFsD1tno6Ln5YEG9f3nKXHlRcRX0HIPbpwJ20ld
LTOQ+7z2DIxuCW4V1Ttpbos7heT/v/QlZieD0T2LV6+r2eQtn5LCCPj3kkJJomXp4gcmyNT+UjfV
FCDlyEFR1kpoElkJbLM/JdHUjSY9TKhucIINDubrD21nTtgiiRTDpFm55aEsiEskVSvSYXANx/Ui
VJBwGy3hBQWik/Yft7oRQI1J1ppAQzPam9+yGqslHEGh7IWVGy+1DtEJaQgzbvb7G+bTqclauO0G
5j3EiioHZv0mFBHL0KtYmHbLKCVl74ADiSIgmFrwe2EeaxUnoATqryOQNdQGNDDPUuAeIE4rVlcy
iv7Hr82Fkct8SEdwy08Bsb4HTLONronVJOLkGvXZGmWNsoZpWl0a50Tp0n1sEJOBriDj4rbsAGOQ
pZybbFX1S2RmSarK1IOdiFEV9iyvwv/+g6i0m3TRF8t3HyEY3lMnBQtt4gRAWOe3XeFCKvMQp0gu
ErPfnLFSAxYkBHyKfFZaaZ4yfbputUCnO36BUt5A6DoNG43CUl7wgkXoNXoaTr2orLc4prLTdR3d
ksNE85uAWbBV14jmtkgYxXtYQ9WjiAMNBtG9UvAqtyJ+tg/MSDgNvq2ldMNygQfJSmiIg3wsKIAJ
YlMQ0jZ6zZtUAaJHP/J6ET1IKNcdKpHCt2kx8kWwunWCsbsanKy46dJmeU9L2KWOELHBah/VzX8I
G6TGO8yTVNWZCyzZtXg+oFjNih3aTaqlbvaX49UHdVAoXilqM5s0cZ90C77SRson/T5wAw9MYSIL
Aj4jIq3QqaP9Wf9JVy8S3dUNd5ZDcPRJ+qMPgH5fdJ8b2W2R3mn5FxZeiS43SHq7bo/YG/AFf1MN
ZgBtOCIm10KILF9n0zLQQ8dCH3EbrLluR3u4ZHQjbSZ7P7Yk4D6ZMR4YSN5ytKaudShD+ILNOAdK
OLaJ/GjLSXmHSlss326ArrYgMjBN+ZbTEgyXYYhprn2C6D9tEzyOr2DpajNUP6d5BFnmWX1Ynjr6
s4A9NdAO8CZZ70Oed0LwtXbOPUWTsaVWXpAZurMnpKS3cRE1nhIsXY1yKmmU6pxSr02g5J4mpzD/
7goBKPOK0YU19aReVJtP+w2lvp6q7xGV6gQcNv0tmarZZMq4NOEan4zvSvJ3Ut72rfOkIlsGOh+P
TnEccXYeDuptf40tk3e9JfD53V7JUpihaMnUzca3VQb6Bb42VIqOy45pZzd3XI3lSE1tu6IFyBwf
lTd0axWIzR2Xy9amSujHTCgKcl8rHaMAgjNstFclbGlg+WbbHIeSJT4mtl7DjNVe2coSzktU9GZT
P7VcW+lboW+BaCdKSrGMYt3LEmSlmrwTr7Ez9ohk3S8dhSWd18IGyqNCzsR8+AiiL+XonT1+tr8Q
+py0b3wo7Yt6isLG9Jdu1fTa5KwO5N3utXYST3BgWjsD0u8B0QajKs4Rqqd3WfULGwGD6AgmXPqy
2bjr0p/yau+His+aXjS0ezVBbAZt+72+NW7eSSSA9zG3x5j+rLGi5FcSgHg96SWeuvbFOkjtI42r
Cpy/EHYsImXTA17L3CThKwllVdPzgJrFdbUXULeQ5Ne0U2NjbjRvFrk/orXZUm6OZPKnaF/evsJW
Vng4esPCdbhUoZ1opNBLlyPZkVjMtzpIgHZ/L7RvFHDmTZOAn49dWBTuIjQvBk5SMyLzFeLF2Tva
5klXxKI/tYyXMQpk8bi3ywRztuof72upFXN4Gw+rZ/XK/uAvYCh58JfexTGCR2lYRYD7FpogKr2O
pcFx1wXZEr47R8HUlshxAUNou+jRMZpk5sQgxFB2q9+mnB8EjPvBDOEBkQvHfDFlFGL9kmM4fRmc
Wq2OJNR4npEoJPIcWsRIL0lE7lA+0aqINWOeJRGEMpKW65S92DqGgAM9iCj0NGD0WM56jDHpMAkz
K47eu0ewGkhuvBaaOHfPK2DGnjnGC4uiIYBJcY0CT4+UzP2vNFJ+JTPJ+Uv1Dw63vFWJmDTRNDHS
fMAyaxbqLdYAsGRv1RgrvHa1N6O505ZvFmp5F8yxIxejoDQySaxJC1NOumfBKb9y54fmUj07XM/H
0kEzIFPDGC+H/MgC74ItoRt0MBT+xVbNzwsZ5muGMUnqY762Sdx1/WUC91jtQsNbP5YEflIH/uOh
DgI6aamD34rRejUtHe73dD4/9NRuNxp4bdqfA1bCfN9wmNqaw1RaIu/DNOZCA6Z0AigIkJCajSU9
MoRxYZbSFEIh0AZc889HGE2F3AGv7stXAmLchIV4u13qz3ZhOfKdg6FLxmxrACfhu4hx3OVulv24
ui5fVwjvj2YKk00ZEfeIFepqZd6tbUK7rTfTIgh26gclIRIgtOPrTdKKTWlDDHZhTuwrvKNxhZ7b
VCLh4j8gRrNShgKEDI2bj9s819sazTQ6Nrh2xp0If4tymAotqjkZL8ZTj/v9tHoIR9XSXo8tLtCl
CinFmOT8nuyjo75U/ANEkMmTi2dmOdGQoHQqlh1fr8BcPCLOC4h6EoAfHFDIb4M4bgK35RskQB8C
8N7fmAVliPnQkd6uziXz12XIaH4DkZ+WcWqqNNrymB0ctdjPlgnNbp/vQCn7oY+Pg79tE/9MkEM7
fdpXhYJimxhH7LrY9i5xXHMe3kXtytl7MBGC5rfJBO8bq3UYKrq9xgA4wCIxqmMlcsWqUtb8AOpJ
WJ9yGf9SB1ENNUwHygPdlbfIkvdqcf5X9ebcoyy2Nk54DZfUOMZm/9iXO2z/4TiOmwYdnAnLpytt
VOb8tZRfr0Cj+htK/fwiOmu1AskPgm1NRAsg21aYJZdzhf1Af7XTh9xW95jO5jd+E8XbGlEKMkZr
XBCUfdf1HGKivpiOAUOASi9EWVLzI3nWcE8qltFrRKDD7my0UzGIVEokrmcWxUuj54R8MEzPRqbH
IVKfeXuXacauUBu8zsbEku5X9Z8K73UeN+oxS3Ao9pX7HSvGjZA/Z8liEs59FmqCodQiHmq2C9aQ
Uc9bdRPzzbzWzY5zPdsKgXXHLWHVydkegeKDRQ3IgPLBohY4/I1SDRL+60K/GKkfA8vPZO1e8y5/
d+YDYdw7dAcSuot0uttBdTvV0zLuvnaim0B0LkEN4K5o1JB+BJcm+s5B6GQSJCQ/HNZ3pbK65sjW
F5RaGDvLvo7SOdeREOIi+S0I3yzv5+0SKtf6e7tE0okcY2N/pKfsuTqo0Ljk2SA+hehZsp7CC/sG
qSboZTdJKfyFHY9wsHC/w3XeeGC6MlmWfmTGmJ6TN+FZ9uAOOG5AfnT2uJA9hSlRZZ7PQn0InlGz
8N356Y3EI2FNyEfASVrI4trI/vnju8FuelaEQlbQDzStTBG3lQAqe2gnXCLn+tk6N8+uF98V5smf
5VAyTFBgNXEuq8efz1G70p1RC6Q4CGXTqxZZUpNCepY1nAvjFojeY/7hVWrrSk6AaUXOFCJ0Cv4t
JFRBXXOPUNj5aQJaO4PbPmHELVbJ1amUGC7Dm1Q85OSKNvZyMm/2EjQyqwyZo/P4s+X+3U82rytB
45A3oLhYnXJkK+EjQJJjP553PYGUoiLrBstNADDctUYiNOkZH4C/IO0v0/AY7dwHvZqcY15ZNAe7
/rbiMa7FnNMtsquy3zcKH+FXLRHgCZRYzOWXFVG8hQAlSU+vqwLUJcMI9myDGWIw93eIBv0Jdx9y
xEC91YjoKSE5QrEIjwOMP7p90S2vlJI5MgLlyUWpmq5apI53Q+P130RpJpm7ocujcebaV4QONaZT
CuICRQlL0hTIyuzsVKQG+Nc+hqplwFjzDExG6TZZQYUh1aDWLhfTLaA8Nji3VMx88b42bz0tASgE
APgi3b40JFMEmgTiD9YlY3EK9C7xPpEaDv9BLAlf/BSG/sW4pVflV+YnVk+FyV9EI10uOCb+JpwQ
lFkkuA+8OKMjbpz9YM52ZQdpRt09imEno+3QEk2MnUj+qmkwKx6GY0lmuCuuAsHvmGu4RimYrtYq
WEeaT6AV90VRVS2w4FfsQMcPWPFWsAG6A7Mfi0oV63aVwkwYssQ5Hp7rVLl5an21vpY0sL5x44ai
xImBH/1BJKl2aLvbhb0FVqOXs+thu/oLtmPQJRKmpO2t6BRlQRV/qDbZBdck/mDl4+qA3eg2cpwd
BHSMFwhLVtY68309m9lzNI+kS3sIHTob9P7qETZcOxM+MMHQ3iTN+Hv0FdlIIDYDU1bmeDnIMRyp
pZrgBkdFpAZ6LdIHkRlfkCMPsjwngM3VZQTAeAnEoMCXBQUPbEfTKh0H9d3WjS1ZCRvyMOv7qgnf
zpZ02GNUAlClJO/OpjklhkM6D/PWdSai2V8mU6mh3Fpb67KHAy5+C/1Pju8qqF2NNk7+L4IDpzS9
R+Dw3N/fi7uNAO+cg3szvDZ1hZgOuosfzIc3YBJbTBM6BY6QndpGLn/SmQMT69hn6Cu6LOeYlsmv
5TQfsL60V4vOpedCux2mTPDIQu4AUucWigFa0Zl+CW9IUld8f4B9yUrH2xgCCWCeDDBbtMl2tWoF
cZK9hej2ZWjCkxh+84Nrs2Mg18uMRnACcuLHF0Qltr1wObZY5EqhqfY6z2J+QHHiwgFHpgjfE+ig
Qx9NPP5QU99nv3GNAyBYE7ohSvACRawNKG1uWO0M+sHXM0iX4oOxvZqdXCJLto9811YkDYRYIEvl
RhZsz3Xl96BPqyplndFmsoj3d0WgLvtJ7Rs0KJhMDG6hpFsv6bDY7NKON/4x+e2J0w4dy7mJFF2o
ka5hB8ukHDWDdL4y2Fk0wznLc4leCMeitm1m2aFDotjVRwymvM0ap/lrykICO7xRbzjMV+grwtwm
6ODEJqBaVK2gsOd+Ieq7YuWDdfLnm9V8xnTT8bbqi9mb4tP5Oqh2UFsRAtltOX+BfWLTVvVBFsH1
y1V17q5ZHhSBwHll+Qmg7TfcBw71NvvJ1AyaRX4+9SuDDqbKcdl/8cBkyDifC7+OlqGawm97C9Zs
jIG2YCB85ukyZtxWW6xSugk8Mfo5nrBLfWvbr+H2wdFIvSa36U1TxNQo2My9D71e12sArcLkh0A+
a9Q090UWIxPaSqCGXXQw3s3MCVmTRZRKXGqjPz0v4y5hr54rEr93+nV6u9uKhBlhOlwLFJr9Iye6
yv3dcKS5Eej7xO4QXE8fdeddlQ9atFbKTQ4T8cMm5JR8iNSyDEO4eJZYegH9upXLeAoRTpzwkM9g
nF5OJnwhL6EuSv+yckE3PCHRSnT43zplcRfNVjGAQjQ1lzDAp6I2pA0m+JQdiulpHAjgRvayg6MD
LplPjdIP+9O7BRwo6ay+8B+0utzKCvFMS/RHSXHL8oXGZeepS2YDAUgDI95Ou68JEc7LfNIp3hhE
SsNxoXEQLZYPVHbPlwL6Sz8qfkzFsm8hbcXTRZuwWYs9Qa1RhySbojhVsl1six/45EveugFXgrlR
3Q/kDItKj73GGBWsahDbJBweq33YJpK34LBh/NVJuG/x8kFnaDuI9w+PWghOp/xd1Ld6gkpkipP9
AQdf8683eBqC79GRsW3lwmZnIZfZ5n5G1Rkmnph8EFd0orVQHvFbo841mrOethMXFIJLBszJpTy+
fW7xUKuTg6xQ1PPD2dNSFtPC4EgHuv2NlCQ1eN3DyPgCL7izrfSIerVGT9a06sWs0FgZk/oGq042
p0FoN1FO0sRry3rEK2GXPwtK5OBwAKDDEP0PUn1UrDQGV+1oMSKAErtwH/1W9FG1qSe8QlSAFJot
kHPYSWeRY4QaOoF2hO2WcwSHOG5THkMNi1T56Np5CTZsmVigbb4E0UbEVqPYOFvpkVpyeFV4jhEc
lshlx9fBEOq4UBzH7FLLAkJlRVqsfT7xW9rF5hJNsDanA6b+zt8hHhb+jt2QXOJApsfFgcRvqOwc
LC4+XCoyQ4k3Cx1IVhyRKuh4UgXFJxxNkRP7j544PnDRKVq5jlc6UmseA0NNxAH0vH5oEtwce4ks
9CDC6du2SyZ+XBprPPngXYk4vPMBCqG5/Gz2ONfS1TTlWw8gjYfdNmIESQxHTA7bWx0yIH4pNQVJ
Rr8K8ZCpRamtOHUtCKHXSRG9cc4aO4NpMxxQNDvWu5Lakuf8fn4OmVo+upNEUqtr4l8VFOS8tMxm
oS0s5W/F849tuWpfAJy8mOa6D10uNlQu3DnvzgpNcXRSp4M2LEEdvrQawRV6WmA+1tgI3nnldr6K
yGcAAlKzdgkCcM1ZgBF1g0xdUDp76oJ8onFZDs+Z50IvxxtkyvheRf8VU5gkV5fsIHaIBZxvLZdu
BuGxWbdYtb3Il0gkCROAIuM5k+1r5kkWrk0B67f9OardLlawYm8VKt8PUeLeGKBiO9xKnt9VHaXN
EvNrrI75h3PxPejAE4ugBKd/dN6vhRFJIe0nKBgVaj4479Dftyz/Kzklrcr6bD5eYbeoS8WtsSDj
bP2pEnOA+yN3UD5CHT6Xy/aY13iQzQpZRSIf3DIcJJkDFB2tfknY/rRlFmg5OpMEkFzK8hlUn1Fs
wSy5JBpXrszY6R8HhWpKBynd3LAwHyw2hnF5sU3iseKaKjwLtN8P2EDqSOFVaotIjBWITxHtsLf2
UPQ0W9Dg+pa+bJ9ca3V4ldkj6CoA7AI+ulfySvon3Z2hXMI42mikeAhmKcRpcnXgS7GjQTtIvp3a
/ZYGTU2kQOtGDqbImS1lCMULjC03gVZbi6TlXrF7tHxsE1km6CfUGvU8TSLLXUlTfB90rq7m2P2S
XXvKH15B18Ef3JSaSHYM1EDsndj3JVhg2CYIyP5nunJ7akHhgPIGsQ30hC1gZuIPDvJZ+xYLjs+x
1QebFGiYr7u1ysQ+xpo8nnff8CZ6U5hDL/bj7618I/pZL+wNSHEBAzfPPDUTF/pP1z0jDGc8Muya
+VxRjlh7NtF2gKt7qFZBNbNq2E49WBhlAXkt3GptBzIO2jf3KqG+dDg54kfFDEEbr43FCYwfomem
Xg2H7b8dCUTNgm5lml+3BCwyEt8yRztTNBsrGyjyVKdUCDFt5l+pLeTLD6D8mpSfFVLM86u/UW7p
hOuUWLId3gtd74v244L79HCwd0v6dapnsGF2n53gA7VmjaxuFEczev0xSijp8uyP1Ze/cZ0TNNbq
ye7T/1asRsaUdicP7IY3FMCTcfjs5eoGam/ZyEtMbkWINeEX5k9WltGML5KVYCfFff+V4SMEIfJv
kEDLrwfErM+n8hEEyuuk51yUVIqJNh549P0N2vKMUgpIxgf2OpQLBQ+b1iPjM9VRwkLe9vuXN5QW
wciJgHhcVmCXhaLmxBJ2kxr4h4pb5LxJSZq2RWkvdQswjYTQggplUR8QdGSQVaf6mgt4bu8E7a2d
p+qYOZcBRjmUgyA4C7NObguXsx87ufO7tzRQbC4DJGkZxMRJZZWalKzjyp21YYpV6VIfhZovA0vh
BxoN7Rd1FLwKLnUwx0MMi+pDCzzMm29GL+OoXQmTBMa9MT1ByShfwyayOfr1oxh2PeawkCNZzMsO
bvIPN0obr1XAEyNdKbpoE1JZqINxWArHmkVk19thAjBxNx9C9vmdFoOtK/ZokO1wHfSXY+5j0Pjy
qlcyQX6dpdtboLqbeu79tkkPAF8m3XFjE+tVXxABnPE0S6/uYa8cY9wBlEv9zGNNhHK6TE4rEN9W
pbmRqkFPb0EumfN3SEfzYu4DzELyQF05RTv8+52CpZ5aSYT/aS5KauEO6mr0KcKds6swu8xhI8eh
ZFTc47MHi0819xdcHCsZ3Eyu8+/Ahvyap9aOPOP9cLf0NnM8ImenJYsiB0zxYVbOMKJsn19K6wPX
RKHNtA/F14vYuDDpnBod3bDmVMF00eQsRvSM7a1ddUy82pVzE/cf7LKWcnWGJOx9VqffZYQ/ogIH
GrWMU8a9Cb1IA9vJ2Oncn1W+9GWXlVzNXGIrJaiCn31vK9iQ7frnzDw23UHzGWuovIr/VtHe8aGK
XiPFWRrGY6Q/8bTZ2DhPTD5ouwRk2oqrhvjm8tZjTJS02vBG3jCFXBbjqJSLdbgPU5lEu/yHBHSQ
crkfge+8yDOQ8cQrOoxzCEw7olr8Unlzv5STlbkp/MdzFud+N2MADypHx+fTIRB0+GAfqgcSCSd0
TH7KCttcctLFMAIQ05gu1a/OwAHYaPWa2oVwx1oW2hgkFhq3NGyOgdraqD8u8JPAr8c0NzV0gvFM
Y/z2/2k0AHZKbDzY68p3aZTW8xuZ0U3ovhTyFwZsMfCQOVsaFh8UmhLP7GXGwXASGNduNyPIHxAx
j43mvjgL0/ppyIxxaVpo3MC4EkP6y1tkErWztfRwIlSI6BhJCsoBwJlQkvF2t/K4aeDKxSDG7kCP
4mTKQQM4R11rKT/7ilelXEj1/x9e/GP2rdj1KvOtn0BLVlxuPc6lDdI+p2w07U3xHrPvpOVu7XfS
wrxgDUKb4b9ayaQcmWNyVfnb2Q0JAqzAxit2Z0F20c00f/toy/+EJi0QhK4M9tL6jnwB5/OK310C
M357HyZwtmt2TEn38XWAYaNRByBfKdLHyW1mxScRiqKPoGFIB/IHLCazj43oys9VLtI+vheP071M
C2AHI5pXG+dURQDI3kzY3eMJHlTcCudjgR3aTqiMmwfxPHNMUOOqloE72pMuhluBUqGFxYcOh7t6
xMB9hiLYRHXGvdFjE93ffoxL4pIr3Ia7MZrjr6mGk/CqmNYwNu9+yX7Pzs+57uxaq8IwqYz3YMu4
cMbVaAEuRUKmfTdPUmgbtseZ0z/ehZ60Ks47ZCeVPCmpKI+JvZ99AsUGjwtHER2/Y7QJZqDmEvuw
2heSPSQpXEX2kWVVTts4pQMnAylG8bDJSbgKbMejf9Mu7fL32lhA/PJlhqpPWdmTcrScKEgx4f9T
eZ08D2Et7UFt0YhGQEQNfuhjrCsncRQkwrbxJFe3VDrik+uHGNNE7mQzgjCv6sOuSkqdjx4Kps0v
X1gk2bqDwlKePzep2T1rgotsTuY4tBkrxZ6My8Z8nNXGW6mgubFWfM+rTP2+a5CC565WwpYqXhg8
TXlSkq0p1vYOYmhKZPtoRlepMBw6xwAtR3ZVSscbj5REH3M4pAbuWApvg71arSU58rxa+cGO5SbW
noGHTdnd/k9RIGZoUJk1kqBatGMgahgoaI8sY3vU9uhIh3EnHKDKrPhyP8uuSWtIMwxRrJLTSJWB
GZw06klzbQATXatqecZK6Hjfn2iZRgekzOWnfcyh3Q1yPz4A3WUUgKwt458MCFP9h3aUkaO1W0g4
6siWtccBQ53WZTYaaCmGgmOwRI3PJ8qUrIR1ElWgMLSBiIP5oYzR5PY/U55YRgXhnMIX6TNQXcvv
feAv8ZcSnGuYoEUiE3gRtUGl9GeiFYFkrs4hz5slH3EvtEVQ0Od5PqdoyPH6zKWkuYL+4fHm3YsQ
oebJ2LFkCmiuE2E6ZJu62YWQKWhDPJDbNmMYTsuoCp/1UjJc+bpciWfO/V1Nx6zWkzE7hae36hRy
rXi1GiVsrYSug06BzkqkIPNwCQQNDc1NCaZLKG3fJLFLz4P6vi4hDbjSfWHFeDmi6cy1xj+nH2iN
fqqRbGpD2s2ezVUS4kv67cG/Tsl+KesStzUTpQUpgPPHU04XBHGC4ZADtmRw7uMDWai03t8l3bX+
C8ki3jGcfhbORzseCrTo0xVE9Z5lPxpncOs0/NBOeh6piMrsUVVu/XO2zbUE392S++EYCl/HCWiU
ar949O47rsJjP/K5NhxF5e01wxCM2E3bknlSuLyxfY4VUSY9/lo3H3YPp+tV9h2g6xdoJcgdLY2Q
lCFENbJFgvKFdRaj/jUqRNgAgEgGqp+w21AqXa+IFobJZIkQ9kfH5HIxRYzFCRQAJ1X2dIfyLQnt
2w0oZacUOWCGLBqFN3rdpadfghMVqOeUutJLd81o6vZKK37Wts9Q/5n+9xona6O5DMVaTS62fkQL
6C7ZefZl9Ls/90q7MIJArq+bte9SqVUtAa8i74syt45a+NbZetlDlhpriXjKYZqDntoVoCmMbbLM
jFcLucMdSaOiahM3f5D+13fkibK7df/xSNIobcQ6Q/Mur2D4nhwHox+oVLpmz23Rqyk2H/AICbie
oF05Rc/Tufz2FaxEucgDpRrbEhyVWcbPnZbNhTl71wbuYywjnDbDzD3j1aPWRNQL9j8I/AAxkzER
qEu9P0kpNeVN/KGbxsp1Wiv/em02jrcE7uzBx2YOUhB5pa6tsQX2OAsqbXnUDstoNaEJqK3wmsyj
kjObL7f8KzdDuGPyL4qzCWTia6r89LTg/wEYLNs+AUfK02TtFtcGPnAbKgyJFyOTs2JK9JBKYMfA
Cc3J/JKY3LM/8yRp8WFoBrHSgC1LH5kSM56diZco+umrjn4arOy093lqpcG5O88nv84JnPXUshoD
ZShCAzd0FBK96QyTjK+bf++GQ8rcSFP6xmv1FtfW1sBCPndSDAoPm1f7tLNSxUaUaD6Ah3/nVQPA
HoUTO2qKkRaa7jcSGVtmT/i7E/pU+gdnfn4SV89XFdVtQaVtY4uXDMQQx84XIcEtB0+uPc6p0beh
wQ+h/fMYGScF7QXQEb3tnGM802Fryrr2THpYLuEmyHCkz8qv8jNwBwQA97MO9cJFP66rZLbOc3Al
Eteb9YOBlLFhoo6IbciPyDVnN9StzB4yl7pkUit2V0OGpxYJtjLE/WIqZVdzuTmKLNoBrJouG3ml
fihEUvB3K16fBY3TRPWUwsPhyIUkgvNgXBQ6TW0VUIlzxrw7/mcmE2+Q9jo8dXxVQTy4+sFWOAPC
jpri9cr8zI3ikggUvP6xtd7jDTdoTFzO7OQcDbG72+Hq/JX2VxmTtcAfpZkAWvya85CF/O6Mj4ms
gaPyxqw1JLyBt8c4Nu6xpcjbJlFMyRii3FCz4R5sFEEm5M0VLQelSJSiQGz+28rg96dpaeDZ831G
qhWWIOvqoDVrMmb9Jc8HvwAZUduyg7Ab9rQ0LkThDb/VOrNb6hJV4/NAeJyWSZ/vGVM1dOv9TOCL
ABGDWgQIiUShrF2TOvq59KLXIpVTK67hHRrlhA/wn0xxiBCINT6IO1UbbCt4KmHU3P3yh7xFvvGN
dyGFzHL5Ks7GZtl3oCXq3c413/m3BId4E5sR/BTUAJRCOjNaM4Foh6w5XluZ/IDe/n+AHKZDlc1u
HESu5PsNxJKsqdQp0xibMbRIWH8uMkbyz6n+7I9/xIYzlMEbxq/Q0c0H+hcaxkSuWKjF/O7JheZK
GaYnZr8tkGpsPJbOrM8MvxxVG9sjUGcjBhcx97+OQ2ae0HEI6nq4M31vLaOBrj5qjsCdSRGOUpVa
YnffzYUYPo25GznqljGL0ReJ6F+nSXFBT0Xe8hWajJSSeBWWlniBeJnYScUeAH++bSPMilS7yE5E
ZiTtVT3x+4TePjKKAQXO5iW1pBBbQG1ZcBR3whCnx4QsffeAEQdzsmFxif90tfzmw5MCMfbMg6lf
S6dKbD8x3l24qN4v8OCOS9vhSJ2bc7pQI0HVMS4mIW0M9xgu/jSGl2ViiAp8aUfraobbyuZwCowq
JqwnxJqADtG2QUhuhqT1+8p/uuUhgNANTljOtY17gmxDVfF+p6XE0ByA58jLctq6Y2N46Fe4XPMB
gLo+E8/ZAfMkJ6y5a5TgrRGDVM+J/nf3uewjHn+e4IDNPqU6/Sl2I6UHNSTRBxOzMxLV68XC3yFk
La5jUNzNy+U/ISbPXcwKIXEgr0xVRDwkoVTGCP+1nOVp7bJXu0Ko7xpAUO515/nZV6QC1PpSL5X7
OtpzExpqDMAmoELX+zyqe8QiHfKEm+4dagEpcjhR3+ZYzIgqON3ZVkVnq+yjBg6Ll5OwHnUapn+r
jnPKeCo4D6Tb9Zk3clgi2os7R9QaArVROVthazIfwXyqvhSU+LsHNFChO3NC43imXewhE5vFtdkG
r76ycLs6zndBnNTtitg5C4XmVCb0BYScIXTCH4hI65ZNTgQoniOUFK0hgqgTYjzJmMYpaEz7FiQ0
DjIrYLDWitMghdy6zDFBgqeBDqWQIUjTMlh7KoBeU0K0EcJMRb5K8h+dnw7+Ay9jdR5VeKZSMJEK
MQugxoBLCk+t+VTCniOHfylXyYB/iWAyyqE2yC+N7MeHTbibL1IixM6JLhjKm2G1TsyLi/JVGTvI
uqO2VEjAivvELDkXQaAp5w5auFMgxodp8W/VWa/oN8H9R1H5DrpGFGO6qocRZs+2d76/m8nKkrNH
XCYwGxFK4Zt8nhK3MMeycFB9i9DveM/V27bS7W+khhs8//JlZuwVQpSbbUj/LD1jWmRUOS1USMbR
D7HH4MfDhNql/YvVHysic6eUcVTYlTbzeb9LH/Yw6vC4FTfCQawWTRXNfbDppVQiYOMA/kN/X8Nd
ifUMDUh3fI71IkCyL8280ipx3c8/ztUj5yv5QplNT8icvLYcHY+rWYp/u6K1Z1VGLMApAMiF0OLu
taAraFCO2czoHq6qIDi+QkdL/DgcAKp9RhAU7rPv5hTZTLlF4E3gPa6St8uFUthEiW6CzVqS5+/U
A9z8Mno3QBQ66Ubheyp9sBitTzNFt9BxEHbLiv6bsV7hmv00TiS4zBAgeswKeBPkNpfHnM/67mEK
rcFHbxgGNoLe5iCeXMGSND3Hcb1gDsX0V2Vvq6cyHKdJpgmCLr5zrBv5mFn0JqJUdkxH6IyuhBKd
6gKB3jFaOfIo8uRgWpC3BVB5FzV5vmC6dayGqe6us7/pL4JyrfwA9tZT/ac8Gg9noeuylYPlnM7w
4iF6tBq513QyiTlsGSNggAlyQgFO8m21mc4CwuNXFhbLPbXKEAJs7ouPsHPwMvNYlCAsoV0hwsmO
lI5/rcMTmF0sPtUsiVgE8MQgIXa+ch540rfGwwJ/xY0Z3zSGni3DQ2e98hZ/wwYQv9ptmPUBQyaG
nbk9aSLpVjAIgK7IA9kN0Cojqxt+idwKfsVJjydrk3QSjcn9jwPa1QfljgyETIzadPuDGS13ioCy
aBDunXAH1VU+D+gw7yquNweSm4VQ2SaHc54ReDkUGtjd4ocUkKHv1IgWAVvxyzHOLvfzd4E/P6x8
xp3vzMC4DW2j3QGU800I0hst9TxRQ7q5ZF55wgQ3du1Cjo7O28ahz+Nqsdj+up3dMFZgIrrUJ2Se
vU6gaH9Lbswicy0sH84xXo3EiGpG5XATgHwRWjZg18ryn9kT90smssh/KkacmpKMX7pVCs+lD0Vy
DyF/vjAwMx9lNDgY/S/a+JojiRG6ZA/oK7W00YWxAy+NTxbxcKIlaRKeodwewa1Av5fVqeoDMqjX
V4978Vo438FIbYJuP3Dv4AUrgVoq55S8eFhPXOFpEMLbUMNb1ZnfxrtkioiFw0G1nRX1wy/K9Blj
Bl/xZ9rOxPGLX9t61n17+V/RhzVIeaK0R264uEGdrvyQ9VM16BvDp98rQBJMNzjidD+ZhL+nTo/m
iZPoOReHurc1dktomdgBzuKnVKVN2FAC/VztCeoiwc7Y+DpgAaPIuY6Vl2I2PVVOp918jLoweBFK
DzWuH9k/W3HSC//jwzw2uQcB1G+d2zU1h3DWu1lsm1OcmRlWfI8KDwnVH74975iSicSIY3pSO0b+
7DmkIuRuy5oxQlSOpmkpUwEDFaP6SUq5FJJTRu0mXXQNDYHQ8U20ErhrzFp0JZSXaQmhTgS4FF/8
AH14Blh4U5JrYxsbKsOfRnBYQkAdp2v42r5XewgbV/PcOaevMcGaP/8Oo537lttnRlIHwEBdAGbQ
nouEw1g9mca/4Y6bk6mCmMer5PWpEzP8/Oh/t4EKrXVpWmpNjG4zGY5rs9NOmPD75ac57PoesciD
0JxgoWcF80+AkXq0ru/1NQ1mfyqcoVXY5Q3R5xx/3pmbqdebLtIaNgqzyCbkvvfcHd8tzGyJldOJ
yNm3dHG78E4xVNXNDRFuO40DwvWJJTmF6X4y8YxJpIPQfO0gGEmfBzYs/z3Uv9/Ec2XwYOHcUQPN
4/6D5BGsnsVC4/wPnnZrXGTGhxE97jE6KySvyeHKW7/mO3v/NRZNij8rqUqc47l/44HQGTJnc0tA
mavkbC0Af8TR7jG2zbYuEqBtsnJOPhoS3R4RcH/EcJhJVFOzN4W+3v5aBgDBFLpJTBfrHUjXpJFG
+jEjKcfYhb0we0T1nYVEgCorvrjEal8kBZXEvoRLEu+NAfbudl+QRfnE7TzOi3QE7OLQJA0C06gn
lYC2SbO/nbiDVwyIidxJ3H2/XJheCwOeal/E902TKJF1Pc639HIjE9KrTdDUR5SYgYk4o1s0sjiG
pTH1vqHWTvvebo2Kuf7O/gn2EKEcba249Iyu+cB3bU9Sai6ZCzGPMWNThr+J1TRGX9sesTjGmOe1
N3eLUZYBwuRkmndDjyqqhlYnWjm/FnhNah6Fbwh4Kw9AgH03ckr0nrDaXdU9zCozqmN8rbWCFhaN
SA70lr58yvTFggEyzLyaPov+5EVhMOXvRGMb/6OOZ7tII7D7riX0dtY+Ga5CPFKV3IsSCBIS5x/7
5/pBsAvfLT/wy55TRNg/yrW1GzosLEeolb5MRhyYeh0ly/C2rC3ZJZu5vv5zbAQfKz5YaEVLDEgJ
sFrPOrJV03tsVV2RxgtWw0PEsiJPkY8qQpJd5VY9XKAiaX4SBUxNuj8rJzgfOX3PFnnZIUNHIT5c
vHTsB0MKwtgRy58C7ztSZ7E0s9vXaBrEdvtjZXvZOnyiLYH5Z+1u4F8ZdV97Pq2WR4yz7N0snyvj
o0Fta43MGHA4AhsGamO0tVXebcRIllZb2QD7kIeDxa2r4NwGqxX7QrprHBxeNEZ/mPIGR475tX7S
osCg0oVGc4pGo2ixz/WiRMJOZXtAiPwiEC4tSNyJKzEoZI+9DP7YsW73ayHyNKvru2opgS0SZmB3
I9YQXdh4PT5D3m9Q1Ch/3Pgf27nNkJe2sV2bfRuJFP5ETaMB7FKfcw9Sr7zeC/U0YUR7TXw3jMwW
X3BathwLL/iJOVKnRZ8nHp0WOiZD6YtNizW9o84s2lutIm0cvYXZ1MqzedHL12ncksYl3VNaJXUO
xYEVSge+THAEdRoH//Vz5SEIzqpmQEj+HUNcYw85weMufnCvK05w8ZF3yjfqNlt+fG2pQ+bibVh3
BNZ4U06IVhn0HnijtstzXP16M+x0eXYzRcJFdLVRisXjWG8lHfU+GzkjYg/sI0YtQwHBGS4diEGF
8JSTWNdkBK5w0JceyvpaWQpbghTKS1rj5+85m04HUNKV8wZVq8C2F7p5oywslaUG1v6zylf5X3PZ
bvraIBujGqEvhvj3uTPYkr/2OTSwUg953isB7hYmncVmJ6e6yawe6VFoHVAGMIERjc+fFFelu487
iKAKGhuWtscYZDiimZhpsDiPm1wiiBdMhNXga0L06zNJEbKQBZyDg9dOsrKfsJjLCKyXFHR9AWRr
AN0b1wKyJN1z/ofBXM+VrWHJSuSCGRd31DTkJCycvhRLq7G4VjNy3gfgILFXEJSoKJcvP0UTJn2F
cwW/2VJy/N1uIPGXGbp9AtFzg+3gNrk3iqAmWX/qhqPHxEKPhX6SjnIWyXei/X3sBkmUCNzH7tAw
TvxvqG7mlV2CJaPczTkdbMzmw9wxv4hqYkxTNo8mo3BaDdv6g9HiCXBHm1ajA9LIdFzt5zrxm19M
pBXBHyVwc9ZzkGs46VxTW2XMMFxqdDLy4TuNxPmrXcH1vy2VasLcIMtcFNB5GV7DNtDUVcLbmzta
FWJO19pKaWZ110Ef56Xgq1Or5QAW5VRk3O2fxOkDo3AbeeV+R2DLjTNg9T1DotxeMWTfBcYc9/Cp
eDXuFnBxu7n0UBXHfOA99rswRHriUrHpHQO3ibhk7gxl0uMc8j4OOwr1cm4f2jsgzLHd5yLH3KAZ
A1uOD2K9YcvDQw1LYK+zZoP1EATFWbCfD12JVf49tYs4Nzzi+sPNMy8CXYNbcZz+i2P+1Iz1Zkyf
OY14tXur5EGe1cP/kuw1C+rRBb8lWauhv+KotImvEyxhC3kUQaYzLo/JjhhBD9ucDeDKwT+WH5eC
GgpLVxr3HRwaVNVGRR8hoxfl9fDXTL37RW3BEJ/Qy3rhOx23KZMI+mZmIm48tcVLPJai+yKHpN+N
vbea8ih8wvHWEXtJrJJqY+/dzpYWJAR6mYyiF6o9bA6SBT8tnKBrDvIp3cI7vDhRAkjN30NXDurh
ejUI8y88XOFLi3Fr8E7Al7Dy6lP5sFozDKV6gzhE2+T2DUZ7NvemQr72daq/ga9QfCIEEk6gLIOu
PO6X5DrW1jkwkmK9sAFtLkPDdZYqsHo/Qp55VX9kzHF6B1q278BH48Gzw5qv0qWVcVtLmk4YDcfo
WRblBZusenWu0GmkT8TsL2O3e8Ew9GMSDlEJxMLzJkT+9vPYHjvOxAOPhw/DGhGLu1LQFE+npUrk
yu/eRlp4yPbP2kqzFFJXpxl4dFiARe2Mcma9J12JgB+gXjZtEKdSs+7FiMC1U64TWgjOEpaaxLmp
hCHn2gXES28GwRCl1kYG6uYrkU34AhgTQxMbchnR24JX5afLIavLT/ssIOtmEL+znECV6IZZC8nX
GihkKpjmwpMAQl6i1u2LUq+UkMtFemT56O3MRdZi8Q5lOroqiui2VO+kt8rpp6NCJAw7u53C9Wxx
7KP/LR7F4MXEKdH1bMf+4W1WMp7doCNB35RJEplWzvWwxgeOcZbay9MA6sOCgEum/mgxiBMH5My5
TCumfOoZ6ASvzngnuHznjCW41NiHyr1QjjVT2T29LEPLSaNxSJoWo3F8jxOVQqw6afKN9E+cKn0I
i1qK308KBp6kpqGyhT+fdfCdhCzNM175M/pCsaK3E4k10ykQKk6uZbkV6rli1yY6KN10eed94S32
gTN2s2SfQgEdZIcOCKUInis+qRZj808Kt8gc5fEecRbcl4HUei937xe1c387Kd2eKnLi8DPmWCzw
qCVUhKHx+slcZ+aY1xknbFHhClDJxx1+gIccx3kgfGfJsQ8nquBXtxnfuD3+unQqZJtYkRlbzBHt
duH5BSQDBTCL3QVQnWbmokKD75aybqFXTFvEj2iQTM6+bODzzmJWZ4kzWGAqv88KSGnJk9/gPtHN
sbWXtOfsitve6//grXVYCHE3hwWmacokEAVmm5pqMKvvqunvGLx3nqlu+lx+q40jTLfHB9Jc43SM
gYj01ALpEvkBbC2PDrEhiuwiOm13UH7GHxYjFF50YJ0lCydGJ3fFVzQmIy/h+JCLWezguTLpZ3Vq
y1MKRYLpnrH/LeGbg7UdQ9rurIurm1bJ4g7ks+24ac59JAXHFwO2rCu+6RljORzAXbxLrh0OxMVi
NrT4FSpxn+vg7i+BVcWERDA0VgJmZG/4+/yCMMEyQ/duPVsXTtwBKmimmtGBxzQGbWK7xhnL7bBk
NJ3Hf1lq6OALydIqOd/lliBzyGWivtjUgz56Q/yK7d1BqoXuj72kDHexefV7h/W1FrPrKx89zBPh
Rtnxe1N72DJKJXb/6mRaoH7V1OlyRqB2QZOyihjqinTy+ZmThvX4N6vPa0+6AULt7ICYZiYMczqr
T+vKCMxCtpaRm9GU0i+BCG/4gigDzwL71ITOGyf40CGu+0XVulbOv1bq+8/9H1eN4Er54aS9QX3n
vlQO2yQJvzwgfjtaSZh7kQv1SW48O1Q82qxfbuI481b4DOfFvTsR7EkhHl0zRf5GBpfv2o4ASkB7
SX/D0a7MUw5/n+qxnsCGFTFGCvVXXJ9iFKb0rDA2gXlmzaH351f/tFZGgzPW5UlfSiEXj8Bjsvdy
UnlF1/brkKo4GVJPStxNAKwGHgBPMqcN/APr97ghFNY67Jo2BEZWydOUf1k0xEyBM6mZieLVPkQt
L8neZ4uLamtc+K9vHWf9W+qNfzyJA0C2/AQHzSOHt78hV5gvP6SExnf4//mk4PwPOXEXPP4Eoe1w
FgHdQcR0UnFfYIV4szPzIhV+YzMSATlz10SZKU8ml20+YqsJvDIscRS4wTutI4BBmqIymZaXeYNr
OprJFVMuYykf625UNG9LNQvVbpUUJsdJ3zdfJv7Eg9U4jIUQnZvriMJtzvYfr1U/TQBfCk1LQKZh
NFDcljqvdz0AgPnHtc86RpyjoyNmdSlD9zvaZtbiYg5p7xRUVnNF57yv7w1G2gMxHczQ7MHunvk8
SD8pjyph+A7Uqrt9Go64n3dqqh5KzhQsGzIYrqdqcxtt99D+jZtB/cIhL/QjkCy+VZmvMuWgg5MQ
5cWJJx04j3ns7NJNAk0ofBTKMOEmaNaDSUYmzATAgeSF2go2bikyqjFoLAQKjxpFy22A8g84jL4X
hHvHxpRPRijjYfBRBqfS2X2hOMnrVyJe4fw2anRpvyNfSrmKtmADGJI2U3PsW7rm+NIHRYeGKG21
ZxN5YXfRpjIulz9zb8YVzgP76GuutbWx3YNJeWDueu+D4JksobKf1rFR48D/6DAiqkLj53dT56Me
jok7kkpwGHsIPEhLd5J0yEqGHp4N9jiitzGeYG8MMw98lHP2hZH3xN4pN3aPVIx2osLsEOy2TNEy
ZNfS7aR1swBdhisUgcnAveqM1TY4vanfN+miPDxieDRNfmBigfdtDVJtzGsQc/0N+s5WwAOWCm1u
HDaCamseQGxNR/HkRXxIVmt8mbiqBwx4wW0yK2uhDGPQ4mV1Wo94/TZMtXHARre7B1KdetdA5VqN
o+obzZf1dvphh53/g97kk72X7t7ya2VzZjhgZjpotvOIpkJXqaUKajp83MCsNJyD6QwIMOi9xsFz
JwZdl7P4g0zwPDco6TPUPS/xMWGyYBVeIrpaimcyIAGnAvkSAe8/6+MP0xufTdB7MLi9B9RMHBPz
J7DQqWzjMfj5GZ3mzr2iUOlEXTpFEo0A98D1xZifLkysOI4F0hNnPTQ7+7Pr/gE5gFj496VzlOiP
tUP+1voM1tF/kIL+/qkKFdsA4DqyGvnUpHoalyfEPTFNA9vHaB1aDRmzNP234NNUedUw4roc9pGG
LZoee9lvWPv0iA1SDTgCuv+stgrri14VT77b/zhMuVD0R5DWE27PeACxFQ55Dce9zRbhKYwekOMx
uPgvzv/KZIyiGDtSjBXRNDzjppH2hTunav42+L8JF+9est6ZLBIfwzcoNWIRi+j/RxU2h3JyV5tI
fun1OH8MOAqAAQIQlh5C9kUNSYSOEAZpY713OLfbksWBIHvVgWyJYhb83y3crYxoj4lBIzV8F4Hk
AEE43K34YdYx5nfpyH8kogjjxI37IiDPkZnZb8G0+trYOQgvFSRQx+M5WOeFZvtZbMe9wkCmLGf4
ICD1ehy3EGtR6zjIwPZavIPPO+SW8FdpN/lnbEsWnHgAH2L6yaMXDGbo56iELPFUgNRSiRXcpqEg
cQjb5ZMOLJ6BQYi3x3Lerlyh1cDTicUAKoFqr1z3yQmp9KjO3Zeh2pvj9BdigUgzoMVf/4YbtmMQ
oYvZEBXn0u959isqt7ECfD9kMG4lVXOjzOGBqFjfW4Ji4UJ6JOollOkVCsXiKlgj7sOoeROCA7U5
IW/Vmb/ywQ1YphfT0FY6ST1XwBCeZeVKFZLfqsACMdpDt6eJbX2NZAhRKiJ4FSBkZ4F0SjIE67WK
p0LBBKQuRL9Z/95cAU+MeCJ0rWYNbjaCded2lC4D57aTo/2g27heTxRrDoBsWN6ClJuQoKiStWPX
7ihfdTmZ5Lp47NAA4L6rtIO6jO9sfn3DsJnzDV9oh6NT91/s7gWEfPkxcnOx9kK6/Eaz2+82/EnM
DNCHBbCcJjHi6Lgbzueo3KUOSiL3/WCzbdnOphkP1rvMEcw6rFPyX58YdLqRSz7WIku1NzOW7x39
/TUqZNF3SolSdDM/Uyk6rDoXVH0Ppxe8W4KTECDe/VdR8ruVLSvutPUYxgia2dsnrh9+5AjVlodj
ESQDh7bsYrfWgcRpfQEOtcvZEPjV/cXMo7np7J6Nbbh1PRsNTh+TNL4LPhIGL2kRj3OtIbCIq0zU
yFUFj/G3Cn6UXcvH/BOw4XZzx0Am97tPY4xrpmBPdEDNkQCMVIuDloIS7ZJjNA5urmVXoERG7U/d
LXiWEXoRYSBZJ3EPGsXH7e5KW9A2+JgSl5WGMrOFiPyyaIQ+jmUVWWeNDUyYuY7cVBSJ2pUYk1Ru
a2uG0+x+xDQcTvv8ShXytp50kTqqTpCxlD0idI+fGSTCpVee9DbJKv8WQz/8WVmCCNshfNm+U0E+
saOTHfgyxsEgG5ZAZnQqn8SD0zcukrggd0gcHiRcGATR8kW5Qgooc2A7xe0jde5J8IqKr7XlO1MU
sE2ECe44dkfS7gtbNtKvMsVbpf3CJj9UoDVEyWszNcRpvqQ3EZyXymMWP8JgzO5ycmycWuaRuKaR
wUFFSFScPR2YY7MiXGSxpETNal1QBpf4A4s/I6HRbFxfStJpmEb8Piupa0eI8cyuJmznYDeu9/BT
BFmIqGDifwpGobcfhMXOcqXAlJt33uG/zVQksctOU5TPZO/luYA43i9zIDEnUhY+a9EnzP9g7NT1
H6bwZcTeq8I/J88Kb3n77Z6DfNYA22uWM2X7ecVCotDgRKC4giVVcboY5Ajxwgt1Mbt9FxS/qpCv
GFD6WszL0SFJLTy/2yLbbDUckYNLiYYV/qmRzDW6L+rlCn8LcCQkdnGsc/v4nyNpOCyXmCGKlLau
B6khVIOhukWjA32Qy9/jnKFUJO+f/VgWYNaOvZo1gAoevnjqs7HlKlR+uSTLneHCsgc+aF3QLwjh
4aoiZIUePZHTW4rGifQlmBS4W61CwpVFBlfxlM1aoz8Qyy2EM7kcxrRxVDhngJHNzNlFF5r8gyTV
Zk7eVXZXYWk/LG+eVonsVbWLwLLPojUq9EfMAr2pc2GJapwMk2nNYNi2qz+1vRHAPhy0w3rS7Up7
4qbSX6ihnnKF5zsPnqhXplfcRWv78vDsDbIlF8fOFlD2UWieH/xQKnxmqaTFVllVbLCgIsGXA8gb
+9NQTtFV9dAeXWUPf44chj4F7+k29Mp5ujloZjGyT2yWZqf/ZRrZNpxzgrnD3RrlJX9i6HpUgQ8b
HFu/mj0iHDiHU6EQ5rsKP/6dABAa3m3g9MCxj9owsBaT6Mn6erXDxKbvG0Yf8QOX0e4OFtWrAJVM
OUvOH9gpeMgJOur2yImSRjqc/fgkGTnWpzTU9agB5uab6ZW3bDD7FY59rWMprHtWbAsBON+f2PHR
GJ2WaLrW8foiqSTr8sWPG762w9AUY/gDSC2YDOoeJ3M+2XgOr1OowG/eCW0uKp7hUrjieoaIu0jA
/BXYVaT95ovx2+SZ23r1AQfGfIwvXsH1+5PzWk2+Fxt+tmiCVkE540QoNj0MJNMzQs7dsVrqA7qm
on8dJjiKr/ZPVEjh+qXbk4m94i1068SK9Da5zpnqLOdAzs0ltbPrVs5d3Djs1h1vsr5OtlNxXah3
ol/1UXJSf5k74K79Iu6ZtAdYXKK75XBWHRsjZ0clzTZgriKoQKAMi3ldIlAc8vqy2/0pzitMu0jY
4moZhjDerQ12OT2TpoycUBbXOLUXSVldUkG+q1kpWo3CqRUT23OTzY+WSaJ+FfGL26hSzJkEMZ5o
m0CkzjD9jU6fNntZWvxJ/BMcKBbR5rzizFmeGqGXxsN1dorGTEK+64lbi3OvBeQGXUB3n1xsbXo3
BXT1GRVqpZzR5Uq/ZLYhJPufvrY+9Al9HHOuSZRH3L4mJippdcjkUO+doh9yUNxR/mCIZ7iQqpZ0
jHk1II3cYKlc1oR/ZNPd7iIQW9x74GnkJ9VH51l6m8Y/0bZlbxr6EfQFmBu8424v8vWmegmwTAoR
zu5RA3ltWXJ1/VgKUDYtZSUAAhGIUqwpAa6rX1yjZNSw3gZQkhabkDvZRGWLy3j/YQbd0BiefVLx
s42hy76aWIIL7Li6zv8qevPta8RSO+Cvw6DgRzdgzXClgGTgX6bzHTs/UE9nyDHOV34n39Qj0iwR
9ugeQyObVwGG7jGTcrCjvZPcYGaahhDSRqPcDEAzhTpzVkdcZfV1GkxZU29GhB56EUROra/G2ymo
WPQ6us5gSG2bfCrrVO9DbJxCqILsYxMvY9Q9Y2Nr2ITh6ypHPZwF4zW3dtDlm06lIfEe3msp/je2
sfYr+wuKAnY//gn/KXej0l5p1s8ORIfTL5B3PVBuHf58IoRDK4otUdY7BI1NRjjM+kXR+tTG9TcS
W27razdpZCF0LxwbmILpGdoaS3iSVwjVKgHNIkQN3eVolR+6vNRhwCzmk2tJj1f/dLPEBHAYnwkH
gyBpa4DfpsrSYHXy85n9SirkVzq74F8811m0/jB0BuXoDiUSbwKPrGGYh6gvir+Qpo8gO8pcwHqH
fc78zfKYfKPMYuWrL4hT7OmBZ/UuLoWDcWLDzk67oeRDt07HmNEum6f66EWj6y1MBZicUlScLJj0
P+X6gPaYKsuQn9ip9NTp2VmnodwILShgQRhDLPpOGnLja0e31sm+RX8s1Vhzk1XBDj1GEIxMwecn
OulMFSK3IGfem2ndJp1idpqArswntJZp41dlB7lXwUe7/2g/NUndNqK3UkDoG5e7jKz/Ppw07BK2
aPRizUdzOUozE2SDu2H7Kl8h7L2U9hztb/YiJLscy6fmJh72Yhy1U1YXK+ho76UJHEDhfJvsHVvN
Eb84HkcCf6ZyQ00v1Qif+Vo9BuFlZ980IlOi2W+yaLFgveUmbT6QxdhzcbqXW9xp4olDrnZuLi8X
ZhOiXg1Tsl6T/uPpmkZdKkh5Gpas8rKoavEB5aB3HnGAqbvIqg9u2wTWQQ1DW0a0TZk7YhHykrgr
n5iiFpWw0v3QvG/acpC6PLSyhZ5Va8k5+fzoQ3D7ZAKBFLz1pl9TkifEXthMAJbi1fUupjZew0Oe
envBBiiUH1HaV5cUZBG50goLxO42VffE9gJErY48Htm65ml6RjyEOdSy6+N/Q8sNxTfZh24Ne3xs
mfMe8hw7TK+tzC7WGYZ/bPVwJWet+2LJhjmgqjT2nIAGHQLYl/LFC+4R9oV4qZo3yoR4RmkxScFE
4ccjFZjMhtvxrCZFFskA19iR/3C0IW8ZIV9wvzl03r/2gd+O6bq1f9eBp+ig+LQwosdSPBlQuA7L
unTOQj6363HaQsuTnCd8UUe8vZLQRV/1yb2fi4CivHifqwcWcylOPE1Lbw4qrRuOJSJPSJX9xsJ1
/5OJMPYPf5kgYN6xSEMiGnD+pMIV94KgbS+99t/LZPDl/8XoC5oC7uXabCAoAj+PLy/2ksKJFB2y
Z5ULATXFtm1XJZdQJHDbV3/rwkO6Wvjuwn3SusjbbWcDLiZYLMvWBWka0HLOXN0tH3M1LBBOZJpQ
r5Cygtqs5cu8o+5K5lvYRqvbUl3B02YmVkqAMPS4iXKgEJqMCBywsMxSs3Ip8OUzihMFMXk3Qrbr
2ZKE2+5i6OS82XnrlvHvlNmTvVxTI9teZH+JDW3p/liCjuSzaQCss8i80tMI/GNYR8RThcDcIowA
bjhftQE7hMmlwCJ3mqAsFSZn3TjfPO18CwsruMNlAIX+7tcJUW8+113qta59xG8P3knFlwwFRcXB
h4fFG8yYR/9xDLFn5klnZR2lwDTi5svLgBa61unLAcjzu1zEuo06Cl5m5QYCV6br1ahzxouBpa9Q
clQFs8renMArUzm7sV8QfO8honZucETd4CeRiSntcJU2s9YzNP1IpnM+tWyBNlI4fXBtGMXcOYma
aINWey16T+dBTEFs5TWTinGc8hDTgvvkQjN3ZUlXeVZ6Le02zGBxCSZW5rqEtxR8hoyq8rATgSdD
1th9kSBZ8J5gbBC8CovjzKtgkC49i/VzLbhjRUiYYLs4m1ibHOis66satfr1vHGzBbiqsGcWvMqh
EP/KGruii2KcZT7byg5QNmVsVzn+crwnHOi6Cq7Rj11jDXCUeea42Qn9EIrzpRJ7T7g+R+ZjNKvI
s/w/skEFaMByZ7bSh/3AG9mfYPba8+ZccJDRoiRE2kxkBSx1ILrGzqH5mKXi1BMeleMPdumMSYBz
wP4B6CRi6pwewY1bgrNJCppyL+LnIAMBrF8VtWcBJk4XW3+W+k25gdH+sic9QlAyOy7IJ0OWL8kl
YMX3kCsLn6wWNhBXGkCkUOFfo/E6MV9uK2wUJMfra4r41BAB6X5tskN7oJ9eIDub4+MLfYkHhZNy
+7/1Ly5+1GJNlOKFr105rYskEQNbZTGqR78WLpiXE8WrTP8k8bZn9o4reV2m5u5xY2SsHYEm3Qy6
paKKSffkbz4JduwWZ1pEvZukUXwV4td/xp/hmeD9oQaIWRWrqVEAkFbTx7GCbBf8ZsOSzeFMIWHe
R/yFErbuN+R4EMuSjWP4nyclTxan+FEnyh4/tVn4TDC2jVCi3RWzOjEul6uk/lglwR7psPbNDjyt
vKQFNqRSNYhpEJ1x3MH12irLfHTZqCAdiSQCATGK4jFH0nhheX/qzuorh/NwPjZxERREhvKDPsHR
nQJKYnKQZdyWLE9zsWbKIw4NhkBW9xJM1XhxXe5WxV2sj/nZqFOirltpoU7eFNb4g6Cwj33zm6/9
4sdh5pYeFCEm8bq/ztR34PWim+yn4Uvpbo3p22PtAjvS6bZcdZEq95n7rNV2TnPu4pvDUI6Pp4Ea
SrOT9dPUyqgLZi8Cb/Uz7oDwwpO4ENMW4msWsEA3StqdXawZ+1pO9h1MCqN+jEfcx15rF/A+Y7Th
QinFGFpgI3eOXsk84UP8iZNCAi+a2oug8K/nO7QW48VbQ4r+rtPRLsgiH5IeJRHTTx/940ts+aiv
8kCUax5Q1vhGbhRTsj0LE+2fXeVx2yprLKRppZ/0VfU44jP1rAbFh3Q8Y0EsoPsplNSeRgoHmuQL
fw7FWdDtk0VXd4PNNZmhNRa1QQ+v7cA9rTjVQ7KQB2FBo1YYoq6GSrZPOz+TPBuBKDnLqTvu2b6c
qsdHMjv+6NLWbdILx7tDSfoZPd6V65PuN9ESDb0IzsTCOFNLhiYCNskcsKmgLOQomoIKE5gG4T4F
0pcPuHpQab5jZ0q/KTaLKIcZwJzOozj0moJLt+rB5QB/lcFoNi/N+lm7kZhMKqqBKnwZ2uwKk0km
xBh8kHaoivSdfO7gtPOTOlyoIcX8EbyUZBXwMrP0+EE6hwol8/yEytRxxjFDdmFs9N4xWGkiMPf/
/zxR5hZqpfu8yAKPRToK4HbrUhyUKt0FDCcR6tOOdmVjBMxuuYuGO5t2CMRGwJC2nSWMopNSSmt+
ZCNzkQDIzAdOqZ2ImbF1YHzhFXdtd3QyG/XVtbjj99TfCUNqy2pK48+IngpkZrCsFUj0/CyAsQQs
hWcDo3uGa03a0Rxct6q93V6o8LpmBRXdXQjCe+P9VyLeQllk7+9gB9Wg5q8sdb6GOq16j50d0VVC
yP4j57lX1KLRroGmQ9mEP9Fsq7DWFpRfrYvxSF/SrtVR5VZKuNzZFYR7j607PUUcxBNAavRlVmyW
WQxVJbW/WK3ruOsPJALjk6Gf8f9ut4wen2cxS1DVRYwAmnh/3aGXm9UwurwV/lOJXixzUoQWbIeg
JD5ZXJkGZL9wO1+G6iIQsicH+Xdq81wdjTGSXlFvaOsNx0eKqARy/7c6Ln5tENYSekOm+LnwKqbC
dr+JAjghgRnBl7LU5FrQjtszv6aSVk8bUKzj/uP9MMP9cN0KV7D8nWbWX1mxGffAminJskhx/4cH
/95GXVU9ziAyP2C7u3hgv/LwkxkQd3+j0UYnp/1YGV48oEsFrjBh7LUr/3hcNT86IwmCCsQDu9XC
VXf/eHF3DdBVaTVHuJM5tQxSepZPicHNmLlfnCSrJOJ40sU44QuK6E1DdktPVTYcBeo8/dmxkctH
nd9jQkosl3GLrTxL2che08bJqF9fDkALDQBiHwiPrHAZ9XJrv5MgKGnWjd1vn/XxTNNNYL6zPhv5
iwV5fXKj1nrN+uMEE1CvSENVI3Hq1P0LiEg1Dw/ztPjI/w7zy51n9l7By8Ya+eoRhmN5mtv0IwMy
UHXmYTp9MDcUT/+2QQSPLBgswDyscEw63AOBE5lSO7Q6zZSic/BbvUztr2r1j5YaVdB8Bbxusqi7
e/0MQFZuEmtGr3zIGDqJAZDSJ7A+1SdiE98R6Oe6pquJiYyQGH5KLjigjLMq/T+iaUnpZ/PjpYnQ
/ud3SSCusqITkBzBJ5d5gh668eZts6XJaqAiElM/5/WPnTkGDQwREbATGvrE6SqvmjQa+LBhLeO8
ejR8M95tj4UssGen7+zWrZD6fd9eWwBMHWEGdbRcehDSc7L7RedT5s7dJbuB/osQG3LoB4y/gLuY
jEq6YWtRkAmF+umgb8jFicGeWWFCX9buuHsujzDbJCQnT+zI2JDZi+GTkkozv5V7QuhF5Ewz0vlE
zO/NGNa+WqUU5ae5yjOPPZPH4JTBlk3dCfeqKtlknD4iXK5A4a7hOXPAmPA4zNphxNogrp+peaH4
1O8kws0y4G248rFpU2ZtSOeIHHA0DfceXHX0bcnWtKx4sk3biZFjQo2gbLji4pInRjYJX3LXM9dw
Zu495akgc6ONaP+PsApdoiaqcitQtzc7KUTWW3W5iq2oKT5cm4Gt6GA3wl1/PbSbxQgXPpukCHZ2
LJxZxJdlZ7R2/smFzHfoDaANkLTKdTdg4Ao5vyGUhiLrJg5tfmT4vNxzWb1r+tZ9B3AEpKrd7K+v
P/k2zx0MhRISiWEqqPNA5wPE0PMmpMOuUK4BH12//dRjagnVpYyl6pTDOsiEarRqbM0rAIyUow5P
V0mmm9B5ZHmdfbzKDW0xBoBD5ElmjpDx5NtkYQCBfpsn7rnBLi8fD1FYPy4YbugL+YNbH6vIjnRS
keR7f6YyyotFNjpaPW3dt/KKfDTpNBYFGjCnjMHXeSJ8Cp3TS+LEAgtftnU9M043+D9ovnmqhMUY
WY2GaadQpdebZorNEnLhdXsvOUrzdryMTi6GMFk9kpCw9dc/kut6etzNZ3S3/tEUNgRtui+2kE7U
hjnh+sDtxeC2WgnRCuo2WndiLYZdNw2jGgLRt7iO9rn5cyoK8iJw7QK1/T4Gt6dj8d2Q0LJS4j38
3HiEpZw+GojHd7Yjt+6AogmFUKBPzcyas4dCY62G6LD8r2D9NtpZMAdwH5gpFoJNMpdgepvjwCIu
j+hFfoJC8DyDnWBh15yPUOoauk+dkAcUP1bAuclxrRNim0k9FWGFYZc2GKMOt6lfpopbozB9xxem
BGOd3ZOyJFh+hkmRGVLA6xDLwWrHAfDe3/ctC595ck0h3KxKuljjHcJC2gXPwUyzxJnepAEptUQC
NFWgCP1IukRa5r6F4yeZCFMp0e+kzMRKqW5RAT7SXxvjR048rHM8RUj7RjEvtzSQFrzBPwwVfgsc
vx683mtOWMh4SEnxTj/IuHEW35aKvZu4mnZZ3WSiu1/cMLWCONjQuTmJr7xLzxMKcr9Kp4vT65ds
q4YSge2Hdu3as4iyjk9ExHfQwN95MFDJTI0euw0xizr23pPOgdEVKRSaHaBHevQ3Hvo8rT219z8q
939abNFBXJ4N1ff7isgK6CkjFC3mHJ7oGEgoqWrF8GQxpvskxfIzpd7pMICG2Dt2Wgv3NNwt3YiO
GbhfHFm0rvLuN6xyDIF7x6S1K9q7T/lSvun7P91EvSI1BYyfFVcV7wvQK4LGHwyRq1VEY2NphEZi
3tF9UEmt4gRGUTc1yPqXh0RUEa4z3xqw5lT23POEsTlfzF3btpaqRDQABUqKFdyNxJSS1ehP26BG
vHIXcdyOD8r+CkbTWC4qbxa+4sF84PHsy+gX/ezqwmeqrewN4wrGfLoY+z7VUvfc+24eQ4kAsivE
k3ZTwbeCtHCPkmG47svCLGF7co7BCjQcIE/vg3MYQOK1r2g+4I20iN+R1BiEXii5bw8U2U6gXrBJ
E5Af/iLosiQ1zVH7zU4G+VHIwkFHiIbGKoPrVFym20KGifvJ+nqCZkVcMCX8NvoGSyywAQHuyHGD
wEvqZ0KM2k8JvfG/xcRMug/aO/m1mmJohNcn1MJgJ2v8jdSGyr30zpKlLGdP1x5YBN18hYPANaBH
ZLfnXb5UyDesOFPbFFtA5L4Pez6F4f+KYzMftVD4nnmooSSBbjJfVHnaKMM+r3IO3q3+lceHynYo
2vc8xQ98HpJyowSAcmbVT8riA8Yh8UQF6EFQq2VMaqwD4b544oe5/vy6QMu6aVtV+e0S+h13pojT
jhfpqElyEI/VdTVBBqlhnVq81tcmwvGpAAix5IWeGuxqwHwiu1Ip6TaSAiYajbRQtENh7Du+kVUV
CLBmBF5I4VmJTZaIDq1fmi24Dqfea2JxIJdh+/umFvBoXQIwihi22mNa7idgKB8HoY7zQ21wR1yz
waO4ESuvEd3izg6VNwrbEKNv+OVZrPrUUxeenXIvkln5STvtcN2PED/qw7i6ce6MA+3pMcii29dR
24hs3kYF9fS8MHo4btDDjr9CGJTMRDFgEkU6xImyBst9wnIoFoK+kELV9qbTvUS4L7Kwl4j9twM+
oWA/lkvdGm+wggk/RrJ/DNgGoTzYccQL+n/JEuW7/rGezdaeQH+6FjtLti2jCF1Aw2Lodv2OEHCA
ui38IQyfqxZhNJKbbDYwMtmK/CDZyM9TAv5iKhfzmUlVH0k6N8PT5DevgRWGyh9GIrvE58JrY1h9
IzidEapajPavYMWY8B5rikxibw8zSFZ+vN60JI6iPUc0v9JXUrf5GPYQ3FGhXb5WSsDMffzLJMW/
qjBHiRg1i0cwYcjGZcj/bknCDMTmpylDPJGkMzqdm5kjP5TTRE3/3MIOp2KoUNdcLxUZJ9tsp1Xl
kQw+KYfY5eM7W6GMndFxsFlJLU8e1/8sQIdcebiLUaj51OcI+aYQJ1AgdVdZoYmARlT6MbK2XUuJ
0bvKyHefkKgJ9ophh3DGNV36gVAkJfQFbfGrGphHU5jat3ZGzC7y8bG6KT2kBTMqOoEpGeap16jb
dx0UXNhcs8L8mi2+dGEXFeBrz3qpsOHAIsPDaDKJk5t1U6110WeV+G0YLPFB8XOXArMqYL7yIFPV
8NpR+dlZ7EC//qW23sn22+lPhhoLdYe8nraJhK6YuKysw0slbcCV6AMpjTo6nE0nTfBlWiwFTGkh
SWvKIPyogp7otFRzy/WJBC12+zHbJmfo3VxVavNv7l2J+wlyoxi4X1tsYc+Q39iTOu+1s+MPYoph
bNy3L5qv34myvSeJ60EtNIAkBdFaprOF2HZz1fisvuc6VtbGywVcfaJdt3orhzsmOW2PsJpluoI1
Wu761Y+pORfzEHwaPL0WCax5HeWR+eVgx7Ch/8W/HAeiF+pAMydospYb7Gwrc+dB9WayXhwMi1gE
A+mapeJ87i490sPtuodNZAp8r9T+dPUNJXvhreh0tPOTuQl8/kmSIK8j9134Sql33E+xAabc00XB
4Af1B1lN/DBzB/pzLJjKnaaLQHnawwA8iZ9ISzwHvF/VYJWKFSYScYe17WhKeX9RSdgh/2pQjC9u
7SV4RZ6oxg2vz/5fVkGjlIhnPe0VgEFtsydvsYVj4gNjW8iXTBpY18vI4l3VIrVSf2Rr9P+Xadgj
XlCM1HXfh3fDeNmaoVmbUa8H54kL4qF3ACY3CTF1ZNqUU8+so/3iRuj3zTSKZ1iPwNdNFWd2KTvY
LcL0sYnqAhLwweaY/iHgrMPrL3fxTGxyJqGZmJQ1NgcEKkriaDD8vK7Sx8xrTHSQdaMLAHoP70d9
bWc+cJjixEWYHQFNdLawR7m1ztosgerdJl4TrULy4ecKEvR9e2bABxm+fJ2kIKeYdO5ojNmthCpQ
L6LFf+o6Y4sVM8Rb6TIs896PVrPwbTOj1pFjB9dVhv6zIayrdUvNsihD6sdgl+BflitwsPYJccn0
9yjSYK9a0ZcSyyIeSqGbhTU34pSgJoU4fbn45xxxPYl0NaVP64EBcCGr99sGBf46hK+aVqNR9dBF
2a66Hq6TBzp+3RmjJoJfZAUlv22ryeuD2dRsODuvE6eo7BcfDaQfnJEGmHLu+Hom9I646Bd9FuLg
ayXFLbYhiHStdpgeMwBtxYbnBuaHgR0Xd4cGNCFgnfeFkvFM64tTFSNP3q1CedOF2CCS0EMLjh3e
UpU5Gko44tTSeeROyXJeR6bK9d7BRaH0mdq/c3zdYt28b6jSav8uhtXfIHxigv8O0RSNWTJCCtdK
S0KUk1/TS9Lpl3qi+OzcfunTHFmtPGt2fyFSUtdwltzDYwucZ1zPmlOmLh+XMKIfrmAMEG8T7BP2
3/VWIf9pLhuqDlJkzE8wKoteVajeJCp/uS/zZjTnGWbSVzEHizp87yJKOoEr5ACYWj1BFUvsDDtz
nfUdw4mgcy/yGtM1VRaP2GoUUpkZjvJhZUrGDYooEFozIz1/MXF5qOQAaLKCYS0aInmYaPrQvJ7o
lrwr7SUVTh4y7CuEmLvcRqYZnKzVtryEwd6ccrs4PkTMBnj+JmfNObk2xegmGgF2hf29IID+Gw3M
8VppvdyLtIakhAbnYm7IPI7NwoPZv6v7c57UxvaF4MGWuK1Ij8AVenJC+6spE5EPEE/dHqn7opzi
U8M3Q2POXaBo3lg4BgWB9KoKQh0OGTOQ6kzKNl8WhxogeB52eiQ1Mgjtxk8g44W5Ehv1LXG/bDm2
ivLGD+JWtvZ8WFyLUQ0LLmMpgorurUvdAcS9Ph6fwZccSnE3pT0ahsLc4WiCyNdd3wVroyNz122p
WTzJtI9BqzoETkBOpYtr8QOgxIHahalDgwvaSGREjbpo96kfaEO4KwWmjCRaiBwFYuFHH9NPvTW2
tQJ2LPz69kzTJKFZveXx6Y65lpT4GEBOOI9YMwUYz4c1mqlCGeyK02ulyd+SVPcPCo9OczgqrtAT
XOYAoFcUfcr3ZdAWmZGTyK4DQsosU3/bOJbWiV8ZSxjcj1t92m3sGeXAuGNAO/fw89+hl9mJS5Op
te/XwMq5oeJ2g1ZIdC+r6cBgM7uaGpKRDGPQtS8sxo0PPxYu9wJko1v8zgYbcgGPW6XjbN0KBCtk
nqFuErK8s4vgtUvBnnf7JYr9U9vkUuKnAPy3g0KsbSJgqo/uiBKtC1RXmC5Bryl1mDgdDA2DGgSS
KFYR7rpjBCy85YmVcvd+aXj8gL4CXywNcW5kxbuJLRhQrFgKp/35CtwNiUr6gwdT3W/uN36bM36f
15McpZrImXl771PnfJHB/kfr8Ds3pM+9quYnKZ/PTbAJQwuk9Mkv/Yra3dWWHCV53gd0zdr0QLdk
nUE+hdpHHXo0zgDJg8SigLI7az1FcUi/jqv/gmpGldENsHrEkbSlh8E+uX7AepwRmfNUJ4L/8TOQ
vSblmxqKhgQ2b0XYh/EjHkkMErAcUvbmi8S38FslGJNTx4ytJSjozl0OBx+iUFcmgEY8FtcCirzp
TJTp5ZVUdB3JRwc6Ar904ay/pv9VBhJ0t+iAX2vxAKe1hkGvazr3uvct6YG3N/lmynV0FiMIPT/q
J50iAHgUz175V4PDottw+whoG/yItHJdTZ4i58AUtti5zZirEfSahku8qGuI1264BGtw/+MwSu9u
jdGiz0ww41kGvqqhq1PAYJQ+NtONaO/o9pc+JJhGATyxoAnowIpxFNmUG/fcVo+KDXMnnBFoa5DO
DCUM+BdJu8dEU8f/0ZyuVQvEYiZGRLCJuLNY9SoruY0saTviQdoLp3jd9CtwxM+y3Fc1JhqXQSfk
kgKg9cjg0lsju2VDTQ3OV5yTXO5cttEPH2+/Ji0u6RzPA/bStUK4S4FEchvXQXeL0vjOvsGbUfno
/+aeHt8dRcngbx2/OGf482rgf5ci6XwctYrgGGwjVpaBYtS67isHz3iWr/xNkERyOWWnIF7bpkaK
F3UtgH+DN1cSWbmi9cc4kcnrJMBzZgLq6LwwwvsjZ6s7/cr8SjkeTMYeWq88JJBKCXGmuGrTBmq/
KjOIY6lImNGL3FvKv4rSqY2SVwgHKuBofJYU/Cx64p3TKixJz+xWhBaCUFCKWg4FFjQaVSOckAaG
prD1ZHkmhI1Nmgr1/IRXulKHpLdRaYivfShJBKFD7ktzeDerFcFirtFbJMUPsgAYItWUFnBqKVUV
FS3pWPj7+432w/x+nt/tY+Ud3Y52y1S33Nf5VEbNmPAEZh4883B4/NAMk8G+1nZWsgMODr0gNHR4
td4cZR89QE7mJib1kMirDq+79ouneyW3yF32rOhLklrkLPt6TfMtiHTxwRAP4Tj+xels1EUqtS2p
P4Bp4y5GJ4Vv7fPU934l2Lb+5LJlzb9krgjb3QZi4fFMzMDFKQPafksjGnsDnQ424iSGtRg873kh
6g628vDIIUUpmDpQzj4m/hp3izqmrgpVVEctzh/SOs2ROc2vNR7il8X3e/bX+f5f5i9P3j4KpV0Z
TBipU8Y+pJNjSTg1Qz9j91xMwhA0P6EjH33Rya2uXg2fFAbkkZVKZkFNGRNy5KIlB+9R+M9XvsHd
tgHnTz/M9jfZQsxBrtSX8owUqqWZGhPhmXPJaWdHiBPyWWp2uHTTuE4Tn1rqRvI2f0kJB3aNsS4Q
oV6sjoCL6v0MMmUIOfE91GW81fwCwP2n0UPx2eJ23C9WSnx/B4LCSfsJkGG58aUtOdbk70fX2210
MUJ0VckV6LDHUSvgNXP1Isg+U23mHX+3tg4zwpmp0FMnAGW8JWbTDMl+LxFICzjHZ/X+xfz1obcg
xjfV3lM7dfcXNFfvWY6qLkqVC8fWbYzM5HszEdwtxoc1uaL0F+oKW2PqYJKLQCS+fmYrujWS6DSl
/jklHdfTLG3akJ9SRF5Cgwdm44CpbGR1ohEFSIW1KxdvSFGDZV38PtTzN28qUvCHRA5G51Ye4XJr
gTgHuoPAHU36QTfqe3V0uxM38dQ6HzIBC6hUjZL6NQUTUb0aWd6Uqt5Bhk8R2sjS/ruHPrTW6XK4
NquqBJfElLldbU6RFYQai6XSlIPWlGbPd7b6wC0bSvshBBbdybSaOmLr+GQqTL7DuvdjelrdAi8U
xfEp7FfIt4WIWyDgp2fLvyFwob2ZCBbVyTTy1fkj8b0rOPBF7rmGMMeuZA2l1vPVBYgecCf3NYmn
l7bcRek03xo+Nl8O/XeiO1YTM+eqSXpb6nO6iH0IojMirb6Ev+NBVH5DeR9MWX2GAr96hKHFoiQ6
UtkEucCdWloKpPfsTKeKMEFeHiyW6hybJXEtW8VvN3ZQN99EW7z/JYcSKQMa4z3wzTx8nBbsqCc6
YNKzf7PK8LsM3yCE1fvPlqCvA+ZfXFaQer8Ad9wEx1WMA8Ibs9d/RspVv71Tr6oYOxvG+TnScEVQ
zu5GOhohJ+VF7wGoZHry7qduMWzqzS4vC7PxzJUKchk1cplkwot4+gekRq/cTvsIZwTj5kGRFTFe
I5/d+UFFDuemJrezgbp5XDhhQxJgUQHNqpTTNzOhgTKTCI6G8AysX2pGxu6hUSCqoxMnXxzg4zzl
3GadNPddVJLlKOhI6zjZ+pqPEGlAdyFEZMBZv8LaSYGIn2Gif7M069Y2/5lZXVFfQZwsEQuzgO7u
WaSIi8tGLLGjOTSq7wvWZhq1Df1v1ocIACQ3zopILqRUa5MtF8Xg45kQn4Y+hnemfM26UPMeQdR/
KLN3rmDK034jl+/ODUYUatX/Lrngxmg2xZ9/o4RvFfgm3MmWNQFVMe4vrIUPHV5NgotEW6WgGnXb
PDngJbR3BGgiEA7yOSG7b+i4wkPfyDeqEA29A1nyg9AYk7NOD+5E4kZ9RvA6zPlAhtIr7QiCiQnv
tO0e5Q1PXLOnrPsTMRJuRtIknvCEbSTB2oPntK+p0zHhEDt/NwjCEU17e8dF1/eiAAvlfbG0mzUM
Qgg8LUOo3LuoURAiBXDduOdzlcsPzYa+iiyWOOG9uRo9TBHgb9gqBYINZoStYUjwj4SYwgzQw3cN
/wG9r+VQkniBbhcrPpKyehq0E23nVidWjPes6n2yo2xxXfNFueAY+5cCBpS+gXj0ZMm0eiMgQJM+
t6dQRZE7eIKcyDj9I7+7OdbyvRdq5mPmQRNxr/X6JfoHL4kJnEK+8kC0HlJugkOUaJcCwMwZADCx
aMUjZKVfuwMwfCfCdoKoqGHmntzzXIzjF2vHeotwKsZP4XmLPZWfEI6UD8+sEcgQ/a2+BYcmX79E
FvlYzaxttU49eSd+PCsmZxuzo5MzK3A3pJR4jgbg7tgfre8WjW8MMUQhsHK/iX7MeRtYwfAqW77h
fDxTDCVrIimYkknVBns7Hjobq+sIE98HSnqQEXSTeA64uK8mGrUjXV5Hy1qgccd94FOwUt2ZFwlQ
1sBQhxVG93eyXQlu4QABqE+kr5njUO0WTaNmCkTZO7d2wyWlMBOXYq/GBa29MoHbNxNZkCElIGV8
IsbyktaTK1Gnk/Sw3U76GUx6S/7toNAHU/FfzirF3tjgHodc7I10ut6eDvpEXZh5imQRxWhNT8lE
Vb4jePFXpstMXnJTJLMPEEg4vkZ9eEnX44iJ9vrcU+ClPovYv3JwOn2Ug76DDjsnUfzucHQW1ics
Gzp8gRLVOdAy3oZnMgM64K7hXQ9eaWcB93QilQ/SoXv0a8scAy6I9Q3O0I4mxR4Bic8UmNHfpGA0
hedXrQggesIXhbE99Ga7DJ5pMb0WxzT4cdMpvBpKtJhImJ7XhR/cFE41FnHz/bAzJFY/mI+RhD+W
nb08WtZ1V9Ggn7uCoEjp4Zx5CU8XSg6eiaHrc6WpTnlRVoYIHCkb4Tj6+SQdGAKQ/4/ssbfQsEls
Ynuf6i0HGlarmGkKmkNwd54ileYQg/qZYBKsU3n6kVt8RPRp/e8DDHeEeZ7FxDvF4rrNEvPrPzhk
L+Tw6y9EzNDRYu5WKxo/PPHHZv2FI849VwhHhOgRx9ZJ9YMBtKdzWUihZlAACyRTi3U+Qh2z7YEC
oLZSOofB/oPRmxndbKbYXurdjM+GlSjchX+792SAG+SBzAjA3pB2yJWYurZQi9Pj3Ukz6Gj+i6oG
ygEagzeq7neUisbL1+Qcn8LDeQqBiKpj9XsqUOirRcEDKErWYgx9caoAgY3z51X7oY36CXF2Rz3Q
Lwy4QLwtrh3lpT2/bWAOricB60B+2nCgpAEcL+Y1SS23sAqSAMzLXEOuElN2Zzk4AdkzbTdXqzcx
KtMrSxJ5keKi8NVqV2foEGetsAsiatUYdRZ8TO2WC2Td837mDBw73epMWGdmrRQMOS74IvFNCkpD
TjkW78uHtBsz/ZS+L/l4y6D71GOqMz20+NxhprmhE4qisB7a3dFN/nZvr/B4LrPlR+U5QYw/NHYw
GCUFnswAJnxQHtA9Nbscg420VHB42d9C1PHZsenw3gZa47+Ples+9ZbPyEGRkBkNwAxNZofQZHbC
CWB5ocd02Otocg1W1l0HJzPN8EN2hs/bC8gdynoqRkb0EG3od9a+h9g/xnsQK/Tnv5BXo6FT4TMN
Gc1bSLGLBkzf7kVkJIQId5ES+oGLxBnbTamtU9mBPMwU5tip2TwnpZ5XZIi7llaX0Q0adpUJbjCi
RluX5wMJWQW+8PbFT0+NB+QcNmKWWlIYHX1bWGNHgXsc1DnttrtqKH5aLFRjYcNS8Dlmr7m3ybNn
/zsyg5ZGcSrl4YsDgFX7IUCiArp6jFNr3mkRZcFS/us8XlB9EmNEkemxQWjL3JxM3wxzIX2HE8Rv
EUHnwrLvBKth6rRuLggFFONaU+z7Wd5g+dgKKkRy/M1PvV9VM+TqkYmfYz47miN7lI4sRjc4VV0b
Fy7hN3D2FBsx7PnEjN1R3S281B3L8PYgY80TJrWRRasxJE1+FA3FrV/rHF1QW9hUFNgnDfNU1+rc
uguAR7a2IGH53+1GDoBVPmBhzVbhyCr65I7T8wQScXN4C2m2Lc65GReA9izgevJq4IiMWHGMx32V
ZNJ534tXyxUzHz4oROe6o0gpKUCuwh2VXA2Byts8WazP8ga6qU2WzdeTXswOeJQkOGIoXudMfWy1
iRRNkVSGrAyZH9woexB6B03stYvcrS3AMjsJJs3S2mkA64ZQrsE6FFoQw8wxHRiA4HkDpqVqqcDh
kmFywmFAeRSybmKHZBblq0po0Ws/aPNVL5qtbahqcUhxLjcKO/+0Rg9XuMJlDeL/3D9K6uTUffCQ
EzZCaoVmKPMxoYUNILAhvDetU7QE8prayGZtaE5SVyrgq2C/N9ZUUenPu7hIvr1eXXrKdKUG3YzJ
mEIesqWomtz+iJiHFoVNEdQVSQlUhYrj+kQYc/PCoEFtfqONoqKpsjpceLDYvJAGfIj49gNJDV7C
Q1edpkhrLa6bJ7ukdJ5J+qIF82a8oKttQMrYxGHWtNGP6CSAk0zPGrzPei0yIQ+QC94/Bpy8KXNM
FU/Nzcwcgz6L8XpkeDsn9z71oyIq/YITv7A5IJnH1JhZeBh9VXNmR+nBVSW9nr8uYm2JJyQQX5Jh
flHiMjSmvLpyEDW8Ev2OwuJp5za1HJumXsTz75n6Vsu362isd/sClbVRLhDLXKWanyPC8qt/Ie/W
QP5mZeaVWoBRc6GV8aP9hs17MgThNtQTc/bh0fHNBU1YoioT/VH+Swa+Z2wVOwnaJmVzdXjWaYQW
NOcty/lfJjm9FIaZEHXUsH3Tlz04tufsZVljYPJix0Dt0JnwKA8zgp32daYj/R5VVlmW+MtQAx0D
Bcfn4NfJ5SotB+xP0TSaK0KL32Qd1zaPVkp+voPLcjpBtWoiNDSeN0/pO5Ik/XSmeGV+mrkVYpNk
BZwtS7TNhdbkLGnvccCyYnb2qaFlRL9unpSEqpbH48CXX+soyuwh8WCp7hGNKJwlnm1nBBGq9EeB
g6XLLThRhU3bVQXVlK10GBbHGWO5plQ7dzmamC9UqjUipjXKsqobjAFF01Yu7sEhZldNr/CCXyaD
Q5HHswzjBFvLnZeak1FACle+b1ZSc2Bz4TJGN0INptT/1ZnkljuVOuSkY6UhlLeDv+ocaw8JBJHO
gOgwLwHbzRK4bNUl7LkS0PfMv3RE9UqoeumQRvCamPTzdmXRs3e0ukMxH/sCfDSPXFvrDsx94n6r
lRfK1qfMUCRQ0zHBgt98iTPGmxT1nXtwr5NwwpYGsls8SuxSFi+ev+4cfktP3bK0iMHLjQ7VNmC6
ctmx3t0AsLmVup/Kyw2u+0SrgibK0gEH95+AjA3uHpPvdSixkXyRx34a6Jk+3yD1ogt2h5G/+q9F
JAnOQBSYHaxb5bAiMboTcTmZvtBY1mu2t7I39vcWWCwyhzyJx/Gm9weJ8b9exgxSU0UJ/gMvqvw4
Oyt2gph5y2eaC7P1E12vAw8472/cTNn+RI7I9ZG/QvvNRrZxNAdU+OzZg0aXNiZpr/o8DlXYneDC
m/Amoc7HFI2A9v3utSssWxqk9jPKc+PrG0v/FjR6vYeiaslWpu7agtMoihHJbQSYDWg6jCMezcXS
xcPEuQlFNRss3OWFTLxcprkUnvCB5mQvrcxbrfTj48EZ8+kNAdBajABAm2BVkZ7tw8NSyUhomNOh
D3s1knIybnptB2FCviwJR+f7+kl0zc0zBHmbwpb/zbxIL+4BJKvadBmIjC618+laO4gvBigNzd4L
UWQzK3Mg3f8vLviznAXyMX7KcdGd//VNHk1BeWto3FtZWfue2HjcpWZV2pdZMi8oOaQCc10uw1j0
uaSxQcBpT/KlEEXXENnRsaVGu0oI5wFR/jrpsmobj3zD0phI7DrS6hqFyxHgymKrhTH0tyuMKT7w
l8ZbVpgz82qjbzv2XPF58Ndj+YNpObm6dCUvX0hTj6a+z2M26/rZta+b0/xZLWIdzqlKfTSivqnt
0Xj4DioTs9IF1+NJmIU4s/QRPoyQMo7rEJOSHBZVuHNhMAJEFaafXoon9e5J0853fqhUFxMmpFVk
WIn2NnyMcbYtwo6TG+zl+Btlv3X8Tr17dj+vBMUWNNkueXbrri1As+TOy8R6sdZb/SKYNIWa4s8n
sTfr0YKS7eVAIORU9QcfdgG3H5646JZ6efH7TGql0kVVZptuBA1sun108p7qGaHLOg1GCPDthIe1
4OXQaS1TNfLUMEJENAsTrEjRQklCEt9NE8sx+UbybLsBTdqYotqIhlzBBn28uafVsI1zUSw3W/2w
FQs6aMrBYYkWuVEudG5mKHb1r8vC2/pu+RPtOhFwA0qcN9TCvSz/dHuw58De32lXnZDpWRzzLgSi
ZM+Iual4IqEaGGfFNK2CUHxogfury8rLPkQ2zkD+DC1W+zhIglqtvD/bNNeNBj9Sj5wI8Yf5w4h2
Ux6Lxd1lmecaZijg7Bnowhp7yW2L5BGTFHFNaHYWEKVetcNZEf151RTZ4bMhIc2uF7h2oelng35F
7MAhy52xER/D8JP7U74f1Z9Oa9faHSVQstZ1S4oAXcgpBZs6GtFxCIi5dtBOI4yv1rw1GjCTfnST
lhmCRlpoeazixrWb9/BfSksQHGkSWx85NqdasWgTSFvj5Dxg5Z+o+VaN0uzJ+i7skcOkaK3zmOZv
5/ipb+SjYkYRpqRUaRmMt+jL2oMgK6Km50+hqk52xj/NqpY02VGMUztGZz6TR5p3K7vnG5AXyt3/
Qf9ogcWKGuCHQGk8fWJoHk+AC7Q1QYF4FaXNQttIIPWW8DM3rkvMMgKSC4od5KNYfRpEde980VWW
3H/okbIK8zveL70oenQA09Cl5Csd+AYX3ZPu0zLPrvwc25BnmsGZ87jcAiK/Xq2JIIRlHKq0UTmU
L0qqcMlaSnwvk2c09ND0EaqkMFudLxRehdCsKsHr0v+3ZgPQrxzRn2ofjjc0lghp/uKQLvT9lSl1
vX+7jHl2lEPCu8AEvFjYGyrpinh2OmuN1kvvP2SaKL0VY/MMhjL7/WaxuSex+uduUQTEFpXhHQ/8
dTVAeFmgI869FZFXcrmcqC4+JAil9y7c1jehf4k75ibHaawIqrTOSKo/mRN+X79YkR3qrfq2aTfc
7wOSFZL00QEURB2ZhNZ9pTtSqquUI1PUisUCdEqVeZ+5Ud/THYHbH1OHmCeYQmhM5bC6m1g7+s9Z
fqQJhTEm8KmPjNkKrY4khYcFDWwquQjqPGHy9Vl2AartApvDG2AfdG2xJgBg4/cmMbUhm47zA/+Y
RSz8vY6PPuQOtI3JQi9n0grfGPqa6MjMgVNsZlsZNt1ga/ZpYqdn3vAlvYupawUO9xD3e+ezUmXN
mrcV1dm4lvbhg0s8p/ovVJ1Q0dwqqLoR18TAufHXK6vWe+A6rJ+rOfuwMJvPKUCmY/UQHLMNR4sr
vlmOik7H6okELu2aKWlhNu9dW/IiyRqhfgcyXPKo+ddm+IELnfnjAKh2ouzOqDZfhehcR7W5jh7Y
auOgycV4SEK4RvMDydIadZMcUcS7HIr5ADcW9yZtIxPUoBupzNZgAgvVMk9TLrx7q1GIl58F+JYj
oxwXAF/oKmCzYuBd8hjiuCCeDkTVr2X+soOZRwK7iAEUfPSM+ZQ/qIv+gZzrQbiPixzLYmNK2xwg
DkTOHxwddtW/L/CVDthNjxV57bBVlunnDg7eWJaTCDioDH8gAYM+tBvsveXlP9dLuWOcEAQ4BlVa
FqDAEKPPL0Lth4SYeCBxjuVdj9pdEnvvtHFxiwIgTvXOVx0yFryVfWXmVf/v6QNsS0J1Hb2CzYhH
PAGnN37ODARuJ8BEbf4P3SrqADdcB55QychXp5LIWsTc/zF88ehj0TfqTLBszBnQC52mRd754jhZ
TRutG60ZM3fhCnQLytAvtiVaW3JAy5hS956cAOy23YAYYpnfev+8Jif1U9RRv839Ywps7WTcicVx
/QQ3XIIwnohy8gw2ex2yJdSomHj1rVNl8ybNsDHtsx1Wb64AL27Whh19MNm+bQo5Jrb0A7ksJhr1
Y2XHNEKQUFFC4XgsNkRWugf7Tr4GI6PlmnmLbeTjgUJ7OeEuJbKgsLy8irnvQDR9KWHr6fF0adBQ
kRIj6cJGZPZB8kfPSGpjy/+GVl3NzX8SXBU28cKrdd04C/mRUhLCLzZLw6MC9MKjH+iKXrc6fzOP
45dfzclVnJ3HFZAlaZv62bk3reOM9uiWl6CaDG41MYw5BwCIyHguJktsBIiCh08OIxRc4ECbLwYJ
YcnLo5JbC1ClOCbIQ2U9fOTkgOcTt+dojs71IMT2NnuNioXdXa+VZf0UzOeTUMkw5pj+xl6AUKhz
nxyHektlBfrCmQ0Txf8VFqfb/DxgkLQmu6IGQmIemCeSWBws/f9R+rjwfuhUhdzEaC7WYqKJuMHr
Av8myilTR5VzkCeZzlsamsZLeQhk6cKreQBnAdlyuMxBQ7bWmJozS5LLzoIv0NXyY9TUbrPMkeaQ
dvrAdk5GuUwzzd4tXpxDn4WDGJmUmccOIuFTRdAGyyQVx/dcld+abJtlQ5bMUwSSngmzdle7E8v9
GNpTuz7JT7yXisV27w0DRjZh2S/sWsWsywtS14tcDifMnyx3eADeDse7t1Nc5LxkJAbDAUYCtXm6
QyaWAjJ5pkajRx/blB+hJCzoZEEk7PtVAcIZC44L9PzwpZRyiZPKWnYtAf6TH6AwfktSiSgPQ5Zc
aP0Z61EYYjppO8f79pYm9eQ9dzZ5JlUI3MicF4fQO8R0FqBoDIyiH3NwhrOGFfTlp3+PcXleJmpV
cI1mCl3y24pydQX1KBIby6pxvtBhHr4Hs49uJZ2ImJ+OsJl23VJuQDoY2lUEI9TnAt5PqDv/IuY6
kvGcy4MMS09uZmts8VBaqGochBwJHpFqhsEXLZcQ8SGIvgSrVLN5CCw0xOG7RDwsvW8W6gmH9e6x
hTEK53VWyNwoMfBTKmggcVMY33UpMLVVq26dYPgUhwBaHaPEx1wK5gesW120BfTNu/+c81ldsK+q
Tq4PpIWAdVPQmIMa2GC8rFE/VNXSpgFWVhId6eNUSEWzSVjAVLcWvLJKCpni2pdgDlfa3yuOefas
nXLaV8pFKUZ9GCvplsIEW3sZq+9PqvyTCWhkLTlCE3SiSq8zy00OtpXxzKa/sQTPkz05FtXd1cx3
efCGUZs6q7SiUKqNesUTF8Ubte+kIl0yAid+8mAFAULfIQnDtMk2CBhy042+cNTN1zKcq2aQt0dR
mexEcFz2ppadZulj8N0For3KW2gW+Qvf7VTqS2Yjv6umnefnUNUJgCLD8aVVcQ6+jM9AgOdFhxgg
EBYOLzaQGkQ8PGRLQFHR6T5U6483xTcjG4N5UvnLOirptM4eM4XHJYjTeccP+lGcVmVz4yWOxdX2
Fuq/NQwKMHMxZr0foz8VUohgjphdDlSw7Y1/uZnLXGIhSksDVKSDh92ZLykGqsaeQ1swziWvAeOs
Q34c8TAN2Iovm5S9m7BwX0IhEv9qIWli7KJW245W9wttDD+SvtKoXE5Rbma1yWaTxWrfolpWAujs
dZ0CccxvPMv/5IhwuJD27+ljH7ho665TZgbi7VQe0HLwRVCCfdV5iL+QHSe1ax8VQbFOXRoE6Ods
eWfkAwx4ONE42PPwNITtAAm5UQ1J3B79KfFK9BvHlQgC9gCLVtKHHFHRoa1GIXzTSNDgHAWfWxRT
fTwcLQGhDhbfsMWfikHtywQP+abS0PrvrKMMM+i29rwGwiTcLOK+QQbC5OM/JaYJ+6AnspQqTUdV
Ga0RQxfwdVFDfl7mWP7HDa+jH8jPOZ3vqeOTVQC0x8+6cuzgS4mxFHYA/9RNVF8iEtExj1MXO5QR
/Pr9G3X2i+0hgmzxvt3f++IPZKrYigZGJz23G6vaEbOjbQdGVE1hi/il1QVsj5bw6oEaLc2PmHCj
8w4ZwsYnSnBkzdpluEzoRTR2l8P+uoxZzvC+S9kzCnreggfMoWu8cK6GeepPmjdVHduQQZiAfAwy
JqQ5ltenGfa7Q3ayjRfM9oPYgE7gzooBdYWVwqPVWkTxaNzXRlvbLV6aGhLqPgvCudKcL1HiSYOy
Sab3ugM6ycnyYUjZ1xltH7mtwSEQri+qHNThYWBBOOAgAsPr1u228CfRnEHbbimMgiWMG6eZxyqY
urK104MJLAz2lWjI4Bdyq0SGCVEORXZ4KIBq1sVTSvcJbQapUmmRMcIV3Uqb3dkcpGSyTCEoWgV1
F1Pu8jkaD9BxuFFqDXEYAgiYK6cl0axNrWW1znxk/W9EZmlFTM8QyUqLjrwughtgiu7ZhQM7BKYo
3sw6ZPHLuS5Izm5VrYoxyjx6IOm+bMblkOO3DuN18iA9dNeVQM5CAoGLpumExvxvCTj54VrGSN6L
NpbbR7ErWGKYGQNdefJ0G1Nwhl+1dew+KmwUwtJXdVlRgTGVC/OsbIC3Wjyb4BrAn59a3XESr/Vd
hK0MJgtkOsT9qssEWvwUMofbYVBXAPEEY0xWwW7b9IMm5X2lOFeODmU8/cb1yL4gKjItZ2VExkf3
a8MOKx6DPEq7H41gjuLGLI1bD9r49xHRgDVh0TBtJgAtjS/b6yLOyTg143zD7R2jVTYFMZiayh6U
aKcXNov7QTq6mey+8GpQGXPwPLOy02fg0hetP0By3QpRKRIY2IW7o0gl/sGV94bk2gXK48WsM+WO
ArB8+eFWRtnARNNyEczC/k75vYm7yx9ATtZDMhHthmC80TlxLgxJ6akrEyMKeQzCuKlWw1MwLeFG
vXEl4Bp/Dy4gIUhosBRXvkAy67OEzoygKHVQhFRawJRU0LFqT4yz/mOVUlAIkDmuuWd3VOi5fHvM
Hf8WcgvSW9GAQhRUjUOAdMEMIimdImgIKyt8MaoRq+vY8GT7S31urAkITc/97ZK02LzyDmXSem+k
JJ/Il1mEdykIFjZK7MHfUmgIexGy0kSrAxN1iWzJ71NpjO5VZJuKZj3zGzQxzYW2RfekgtrZ5hmw
eb70qpXaN7z+l9wSMOqM1WNx+06JdzP64EikYLezGDZinVUCyeR9GHxqPn+ykY5YYPXNwgDpxJL1
Y8xf2ThNsl6wCK6e9q09hYvbxfX8OPXCCxcC9dQDBq0V00w9EzcFSXyeGI6bLXMfXgVsuIEDRhaU
y++Xlb6CJ9m5STKj+1xz8G80nGh+4YaSOqH0rw56hr1xdyawD6quXlCTVyo15nXtlpyPTpaoz4NG
dHrLWM1W1nnb55rIHfsyBDhYzfLfn4GI9cCJgJiyYMCJWHAzH+YZB3lGRX+pJqrlwnkIdFFL/yBr
4HyBveJ3KNnI6XR2oqrvugmtIPXhr8RtMo0jfsI2b2xsyzNFdn0gE/2MVWCm3dd13wGOpqLLTR3B
PsAwJ1Y4bV4x827nO/yaIT+D61oa9MVo1YjpT3W+G5lo+HPOHf8t5ORbOEh9jsz6foI9+niYMUA5
ByJpKVLZ30BRyjVoIw7536HMxvWzJEJOgNN+7xFGrqiJAEOIzJB1WcjNswoEb9yRgj3DGwovvydQ
slqyY2R12/E9UobtVbxRY5V2Zchwghh/TpTEl81XEQ1D5HWjjv/bT3qM4EDhMCVgmwbbFBmueSD6
1RUTZ0NZf9im7oZ4ySwPG3VP2Y7oTWvdn24nxG9/R6RIbOrtmPr4JVxd/7DqeuF0ewWXRO3j+PAE
040Vrv+Get0KpBnkTeBRegNNFQfAxKaqVzXOyW7Qpc1W9TTr9foX6N6m9TuD+lHaX+7aRPMdhll5
0Iy3gVPaHjiiw5sdHdHnMNfCZBYDd2rLpnU7kdV4lPyPJ+94rgwaVS6wBixBFl7r/XUNEJdnTxpW
ZwMvS3Cs+Jvx0LN2VjR+rC5tSZuUremwsnLVFOHnYBnh+OOWF87RTq+sliErPSkMuSvmuF9HVfNn
Lg0nVq1M4UW9V1JaDR3GfMU9LkZ9sNDjflRLgHadnSpXJ4A2LnGpcy95dyYFpYp3Wyqmd6c+Qvzm
J9sjKqL4USudIbXeVkiYPcgD8NG1uPstjm8zBXoQ2Ai03ZIRBWC7bgjzR/6rDLakNtwgKlXOqB6M
ZSWY//eMSg9Zf/XCKT/4s8xc4fRa6Ho5G1se9fmmi/E5iySIYTwvOG1C+HgSCcB1z0RRXTdLW10Q
N5FNQmhqEn+NXDc6hWg56mfi/kPjA0sLGxFYgefj/EDAB5Er+KQfnHdmUdoSs5FapHQPEmdOUOzg
TkjzMmjRCyuLRZ4OC/Li3KO6p46bS6qRJxSGLDNwP/Rj8SUaJFlC6eE0wfIno2dAXeXjN56b9l5t
cLaDmQ6A1zAJjglVsOyxJg0/WAjjbSdg380EhMQ/jv293a34PXJb/XozK8q/GTUq6lbXclM+v0f+
jfoFiyugtuGfOM66HmH9d1K27+9JUI9WzDr30MCLf/hyMb3qs2IU6dSOgws9QP82z0L7oLO9ZuUB
H6+iMG8zwpzz+kB7EPs+VNiWRaW0mOsW0rtLI5RUmHyTU0MdYh53YIqxCt+5h/n1nStAKkXDdXRo
6AUKSQuuVuHoUQ1Xhv5LPVn5uQllp01KtLSYUKZ+QNVyxEDw/rAcxhRqdz31ZIuHks7NpLRlCEzY
87ZTwhyYl966TPhmwb+zK/zsnNUa0YbtxhxZsMNj95skqssGLVhAhzt9jCUAVHe1ZdwAs2fu+6aR
pUyRAIayj0g1ZCX6q+OueGKKSivPvuorpfoP21lfcFl514P6RENudj2L7cjb9bEbr3evycL9Muhj
q0p2s1aKARgmbgYrIOTvLB286G++SZMuLerlhhu8PtmfvWIPzK56eUR0ah6Eg3rGumKMBoA8bIXQ
M4h0+e4/1IRmIVSITTe/AYA0dfWMBJazEi+rZFEF/LLT7ayrteIC19pebPppUXekBga8SAkDfw1Y
QgVzJUcZkEdx+P6Me7CAi4BvcnAU71uCcTX492BP8Z7a2QGcSTHfmHXs80obkizGOt11dV3tLdYJ
mcc5MM3eK/R3H5Tkdik9k8c4+pQd7xC7aClGwGybu4ujyqacVzj37j8iUDP1NQiLNJ7svU4s5DEY
xpbruCwpfS/xSRHNUd90kp9lUaD3rvqAuXrBuwzYGmUU2gzaoNSwGRwhfJk8gIjOMn4xKkX9j3iL
VGCw8v/tlgdldpX+bWx5U8V1PBcu9CtMjUJBB0qjVWexbU3y8Qw138ABIBaHN/nkiViLCwo7URlC
EJa6+Poo8EUqKgn87cxvTMfYhMezjCiySPKQc79JSVd3QKS+JdxsUhgEV4X+7HQTbentp6FAg3Ba
CCooQgIH3TDoUvB+Vm9RjTthUjTOlL7XbklJ+u+fmbGweJtrBfzRXtvADrGR9MCptZSoVRzK6HTn
3acs7Oq3jymiw9xyPl5gbCaC6ktL+p4l0rlbMNRaV8OsgLSdau5yZk/n+afLv4on5xmGcc0fbqy7
Xb7hgbnJlbtX+gyZr5lQQ6xJ9et+ZscPQf25qm2hQK2k1VORi4kim5K8pVyQ7XRV4EFDDgmlQRHP
BBv7tFmEFKsOX4CJmOvJXroa/Huzcyj2pbHhq3zSn3SoN6UADWrLFQD6Lw0JhUwO81bsZMX1ZQS8
x0/EUqk6Cq5WPfo9VMoaLXxiDNEP9ez6J3fUuoTnr6V/dW25PjCLOZSNidYizRM2s1uwA1PASRS9
qG7ALwxyKKoTD5FpycKtZgPWqVWWALmU5EXXIVWssAkQ9g5X4aMgyj5uft76D8hqvkUWLxTnx+q2
TZ+tYgs/ni9VBlqwhtDH2vYjHYNr8l6x2ChS1PCGYUeDdOakKXpmu0hb3ZHKpxOOwdk2WqoZJ9XT
ROmaco1snbqIspZemIU5nVRq3LV5v/+sg/dbAXV9A3tJYGEMIxmnFOj2OYJCVaHsYf4oQgwxImGt
CoRt2B19iVEEpDGrknozFsOCXC10XDvQ51KKNFQnAiI2H3Izs7bNEI4zEO5iKK95WMbAcYcmuMK8
jkcwZJ5ENG1eG3ug9kh933KbGt8TsXj1RgAOxLJRVz3NIUKxFDxkjeat0Cc1PWVMfUrNqxIvcZxB
UGfcSW31wikhkC+SCYcT1w3ES/wSGoWCSVf2q2fDlCUZSB7AfaxgiXGsFIK1V9QqO+EcBWRJiyn/
rpXBQtFxFqIWwG1jB1MguJPtcDXSaO79Mih+ZyPSqkQWJiFso/EQStqFU1XO8rO0ZbALQhLQlILF
jcU6BuBVk0LZhcI9zYppExfJVnO8eH0xHtqClEZMditOWxBlxro5RSsCZ914P7flYrFCUwT14TFW
htADbMsTiSWtNr9jeLCj9khXc5qC8AOtFhjuOEH3JlhcXKlmKp4zRnJ4KSX9It2b/5YFSnNvObnI
Ojrfsn2yKTdW2V6FAHMinXO9CA+GSbkXYiM5R+qNmPFSCPZZuM1s43yOYsdh7PKbPyZx3JvJsRY7
LOw3sZ7QFL1gavVmpML/jLes3XW9Uw7ZVxHbGUdumbiMeIzekuPhapxEe6f0073wyByCrh5/EISZ
/njRdLlUm97H877HcfHq4DenZ/ZY9po/Al042B07TKlwzCd0ZiED+6SSXHrGAWOJl37TZERN17FG
rVQMBpVUvdNeTmY8nlU6qXKiiGD0T4bIRuZr4jsQeiIS8Yet7pOsG6j2krJ3Dg/dY/8J86gJKM5I
OnjOh9RieagGpDGUbdrC3sccKQY/30oEigqOnw7Q0HZM3Uj89abZR6kWFVN54dFm5TBeaJ1bs3JK
qAXoT33j1sIbp3sBxpVs7g+1axqMVgOApCpkgBWk+5DI3hqSV1FsBsLCbMKH11EX2FQ4Xx9XVM6+
1krLvlE/zVMuoVqwzSV6jMreorXmOmZ4FejRMIZLfEO8iXEL4CyP5Y+9E80enHWQdH+N6m5ymhDJ
O7Ljp+unT78KCgGbw1gZt1qcD3BnjsYywBuOecTLP7Uk1F90QLJOv5EgD8+2VMXUGdrAOMEte6iT
0VjZY6fMhZ3hJzgmsvLQ1R+UGq37oiCsJ842WykrW7oVfJxHfBreu9MerDBwvNs6IGu2k/XuQX1L
XpYYNH/j8k5hFraT+nw9Cc8cij/LpSTKt8X9LfxTZr021lHOO+g/ZYUbcfnN+ISHivKIMQybrQGf
BgaWBLIxiMYdoi0AXh6oImS1dmYw0B7CyYHwS7QX4sex083sH0i/qGEH0gqY5AWkOruAFMA5U9gC
cWZDB8GZJYCcUeBvqzLQeMdDMT15A20lND5IvRalw/yZypqJvWW74EriCi/fzIutwQ/0ky1B/hsy
D+dbxzhKJ74A1/mzjaL5qAmFQtWqNQQNaIwstAxJw3ZicBXPW3SC/9s4y44Fz0KiNu5ekASkQPP3
UUTROmg82ojZsePdImWIF+1tva2dyCkWjwGRGbmHFa570eAi9DAniv8waipwMJoVjPmcndAe+UEE
ZqgV70enUBITyjxHTt3vGF/eXk56wtd70ZIm4lWL1Ilchs18MuQyCGUdRFiBJVCfqDkAVC8czSxK
4MuywWdeYjrCSD3c5sfc57MZt/ki9l2KEt6mgdqRmeFVZl4wXY45ILS/jp0baSwuUtI/ucdhpgQq
UFJrpExEz+1UbUZkUNFBzwfsLjd1b+JVZFa1/OUBy8BMdTN2nWKk105z/gY5OWIZl89CqdGqmpl+
So/EcnR4WADzG7LulWcGawjE56hfw30IasUv5HJuHDEpapZBrn4ZHJYCPV7B2iW4RGULGhMnSCuh
9IVQ4sQjDQ97Nq2aqnX3FAXaoAqAtKucrozzxwTLRJ3BK97eodj7xcEf9itTnH0T/TUjAltqhW5F
35b7mI8c2LMQEYUpW8FJqZV9RajNgGsa+HZ9FC/y7Z2Ackjw+j4VrQJEL2W8cMgXfNwCr2Rril8S
RBqPibcXbWQV4ZlrEyUBoQoa8QlFaKQejczOf1vV6hlEIy5S3LFrCdI4dqkjJf1ccaA4EOOCD5Lq
2c1H5f8NvZUJyqKKzzplbAg0Yp4a2fecBgE+oQXcwezvBhymLbeZjERZtAT8pz1txm0nFtB8gs+q
jHuYYkJpFShwALrhBOEP0R6TxIbgt+AHVTYRPXWCXmGP0mFbid2vfReksdSvLx7BPG8NOnkHlhZ9
+m3poKpjFGbIXgotRyvoSXB7YfbuQz9PTIN5vfG/IYvkBlBzx7Vo7dQ5mGgJX0lEmU93B3AQTquE
G9r+OaVpLpgpNZqNgiRk/cit9g1BayKai3kxc0kGXrfAJ4EvYIG4hPMiOLywo7vWZtWYwxnQTxCf
W1bSyMkJAF4MqbyspVGEaRZZ866mDpdUUJKt2KcD1KvtB2Zw+Qz0o7H9atF7SnvhnaHK3/knWgKr
1DW9WzCMDYkzXz2lHYPSOu/TLP2nD9Ce9YkIG7ij14K4k8+Ny6JJVuLJlwVwIzcqJpoYBZo7Locr
nTOrDzC/JNIdHljR4uK+R2pDTe94cyUVtzaUhm32NkcqXlOl8T2DnxnWb2oL/jCYizV9fTMVfg0f
Hmle5fGjZO36l+Z4BKH9y0C4bkgkENbYtNj0/u8WnSqSZ9lbSegq1URajQu+UK7OY8O8Mpd0DWG3
jobsqXeDqx6Zy071lhChELba1bf/K7mpxzXUMODo23Zx1rWVaBJUK7twnqk0ec4R/HWjrS0FHh+O
kKfPLkdJ0Iulu2Wzw3Dl312oyYk3GDNW7+hvw9icpRieaarTUv+vt9yvSVOKemGJWdSwjkzf2/1R
R5/t0OZAiSj0GLGhiDjRc9zGfpYswjpO0LzFWbD/5xwQvOU2ebGT2HumaqDoCx/sCu0wau2nFyl7
vqUmc//CBzA4nbtV6+yEZLdbNMrCB5isSXGB+nx53Eeps9qUXAzB8Xl4lsmhUowKAwbPaXQfv0wr
kIXGDx/rdt18gS+f1c7XGKEILirGW1fHPb8H4WRQ3RcvEVeOb4DXA2+AvA7y2qEcas1dFu0eDbA9
XefoZ/rxrfd/tAvaqi5uAOqLD6OZyFUjAZje3bGxSjl1xvN/YHfBIfbYbJ6J0V2LSC4EIKrPRnKp
8CwVQXpqGGxDqMXdOQMqMPnOPsaLI4ThOj9lFX5pV3HOEQSJGr3ySozPkkK2GmLrcAmtFBLPma6N
1PIzpKcNWtYJKDGjnUo+RK0KQqlCPmcDA27eHxthzQ9SxxV8FSFvVqyyLskZ7l5Ge7HdMvCx8BqX
oTWpfECQ1bmOQJOQmsqfVseoyi9+A/9Eun/KU5U0P8WymPSe6RNSimntXHXOAQTcaRt7CMVuVJon
ycKBd8L/wXcxy/O+wUnxPbsWhKueWEDUD/JJ8IKTvlwiBQxlVDfoBMQbGCgwC5ykl2CPnsW74GSe
XFl5jVxlD4hxMtGOKwPugQ79bYFn54YsiciC/gSJnAgnHJnF7QAJfqmCarsesp2LQL8Lyf1UBtOm
OlRaz6z3QuS3IZjEP64cg10Uv/Si7vhylt6K7gtNOa5CHxHsNTXtgDi0dg7RNgdvqHuZR/kRLal0
rQgNk2oXRdiCsFtOWq0b1CFSFCC+xGyu8fh9LAcgoCoPeFWp6Pmp70r/KuQoDJDlytRTiaW+ay+l
4H/eJVxsmr97/MtSfjjaIrNx+Rf/BjCmVwizL2sQOIgiKIfAQCRM+6uIerNCq+R7y3USDkr7NkNS
KS8eRPcGivOkTCbUuM9XfIxyHtCGEaGz0BRVB2zpUU/UjBGSLCF8yvTP4yNG4DA2s3ZPHhIkyG8W
lTv74TE2O/vRT5fr3eL8Ehez4VaPNITRpj7H3tSbGAZOIgOngsyHcNcE2Y8FaS+12zurGxGCUEhA
/cys1PmOTXMQBV38tTlP1Up4CrCr5o6wMN0UZIdwhjU05rnlCGyJdJUhDYr4BWiTjgPz0AkNJ22V
hi73otMBjtMintcXiDEOLcN1hqY4LXq6enE7TUN79rvlyUtt9Pocr3Pe0IfLv6dCkY8N/sD8+0Js
1qEyE62yB3qfQJ0j4KEEj5M539izFNMnsjt7Rrx0BMW0/Mhg6LU9e4zaDbbQQmQ2Im6lYOWFaP3i
+aoHU879e23uQW8o+ecxQqZItySHGmhv45wXSZSa7J8q3WFztCskEfnT+Z6vAi1IZWToddmpMH/L
aQEjgg/+iQD4CZuQCZCPtSaIcYS6h+6JPOLR4tnac8VogkmSqwWijwPFtTTOQy2l9sNumfh2uXSS
ZEQ02/lO/8NbEJ0POW5pyNk4asBfCDm7R61DbN7w9IuM7Figh3S1Hks6qAICPyYd73EQwWT4CHDb
FN8sErvfCRrqQAwPAosTeK0pUG0DIToHtS+jNSq7KpuyYywvX477Wsj/i/xAoGWr3dG0oYHN0b3v
Nfd/kZOEVU/JrlJJPF4FF7/5TDnZ4Ju9vubB9+t893Xur3S4wDRrXfcSo9OfcngjfvQJd8f6pojv
jRLd7UL6gdDfBACLkt3Z6MruXVyBsvaGpFebNVkESTe/7Wlj5aJU5rGo/0ZbdmWjaIkBhlrJmfir
nh07HDDcPQfm9yr+oUkzqo6mnuODpQfTt/Mg30U4xnqKIfpgHNiizdXmnb3N4IcmBwIsTY0K1VKL
bKSz3MPciXibpzevPJsj3KYNH4Ji/F4Eo+oHlGejHRRjXsWoDFFEZpgsV7YONcQHxNZDzrg8p6ln
SmwVfr3WgnrbOshKlRaCRh/ybgkXX+UEpnNeSyCp0P+hvg3vV+sMfHaPPu1Re7PpNCpw5IzYnriy
2AGPLiuUww37/GS6JlZ0XpQdJW7puhFEGw0pdRF6zBPpHcmG51KGIzEoHo1PqJrkPPfoNNZxsKn9
EelPKXkKo9N30L8IaxiF7ZvIR0VcfNgpq7FOszFxzX7GcEaQfU+d05BaykCNoQz2afEiqaEMnu8f
n7AVRaYcA442zEuA/JGXdrpRR/ifV4yfc3bIPblcm70CuXG/j0ZyUzu9/qtCV9lRw55Pusq71FGg
+TSF+7EEA9/QjsKyiE7EQ1cTuv/SpxIIOWAV2eugel18oxwwC/UapPEjighM+OOIFWvzM4i6DQRD
clXYUlJ295DrbAD7NzH2UySys9DLhHAlQT82c+M7jM67RCnsMHtGmcvs9CNxP6CqNTewVWI6TaP4
eGFobTYkr1RzpnAsCpO4Mk9i5t6x6l+gbHgmVi9xJ29hcbI5dt0zYsz8bp8iJTzyAKSDLf65mIPM
OUaqvA+qVWtQngJXaXPgGR9wM+9GY/6fktRFX+2TF7vK8J6DG9n4cowVPPoqiBy33HyqTZeKNpx6
vblKrpItp4LUWTrb1xk9eLvUv1EVKRISPDQwdSbifpM5tDnoukx8i6iJ87UVKD6SYvh88BamaRzn
DECp0aYVnwWdIVQN6lkhXHf348xHDrll2J9MrPOvanyckABFERYALyqllsR0ov39xOBiH4lURaM7
fRCX5NnSIgNmHcKGptYCEc2f3b1/fUbmXPA6BBCMOky3vmCxDW9B9Ot9HC4uFFgmbYO1dbur7swg
e+vGhaYk4znQgdNT/NisQIZALpDke3qn/RhfTVtgU9wGvV0jGKprCe8XFU1nXr0l8aoPCyR38Ba/
UyvQ4u5uaz+JuevnDA85LtK3H3vrt2TPceRuX2NFY5LI0Ks75AKyEDQLAXyNgMO5la8v1ccYTd1t
vt6zsGHauUKnxpOwk+BnwLE0262cusE3jqbZUwSG6so57lTxJgQkgI1rG6WB6j8gTRu72EpMz7yL
133IslF48+WDmKplqIB2fvHW4135gAbPpE4SLI1taOjEM6XIMZaHh0oNfObDG5wd5OtvBAknPxM6
aAno6cRtaL4IAxLbzdWA1WRPko1bT9uVlbAxNR+bK6R77H6gxoDGaInRwNPa78KcQ/m3+mPhgR5f
cpIcCpg5D+80bWyXvUuqgr3ApfObGeWvbtpSHuZJFpAZ/8o7I2u0Q06+LMTHxaQHwgbKsH9nQrW0
WmKIioUSlJ3DGxfcblBmb8STewUzgo0fc2/IWPImBuuGD1JtZIlARl3xPIlYQzKQlwMBYKpiOJ+t
7dKyAfCwiHWMX+zXCpbkrlJl0TQTqe8eeDrUgnjUiyLtXQ66fvYAMhfGFeRtUE19Zlju5OV93Spg
Zr/9jk+jEmkBK1SN4b9+uitrtsnnrkMEqtXllHeLP1RAXPG00HfpEMCFOpx+Nttg/+55K68QPDOd
6cUVy1KzzBVI8BFPIQaty6Ag5yEmjV7knHacGlWYLxOoH8pTancRxMAGyUxEoBzK4LWyQ/NEZ9uf
Sb2Wry+ylsEsIcVGTiYDLp2UaHWpL4GHRwtv007aISiAUhP+lM68mm8l3uWhtYmZ4Hr08qvsPprZ
MB1RYVR9quoRYPwC+NgLqfk2gvv7+WCMLWHIIPEHemVLcstilDQTH/vf+rcpIU54aslRj0dk4qUc
OygToRTnWK9+ABGrXRoPSVCs43n+m+kEgG1Jau5p8ocw2317kyEq+WCkGLN18iwSANuvnvUdkx+m
9+Js6YjQDyEToxByIvLqZ5N99owW+F+ck0F6YgBFyyddASm0Z+Z7AdxhJPTef6ExjI/CLvn1aKyA
7QRHqOqk7VaXBI8mqOIbCUIn3dcR+FYERQQ3Uu+SfB9MN0YFu3qrYsemJsH+qHvXTnby9QJ/2aea
lladjZ641qzTn6lF/oZTWWQo9qP+1gCDGMDvuDjDdMQzSt05PADox74UIdv4EtFLtugD1J+SbLsZ
tx/JWwYHCwfztvhuDbuoCD6RA4sd8LqHMB2nqfwtPhimkotkPVYij2ysvzFPMA6aOw99d6qxuYGL
IGTqEoJ3DplQvVZiDlNVSnTxM/lSQzCCXUxSF111cgsenV85wq/USTTgJsbhHa4A1PczlYgcr7aM
0XSzf+b1F3pkN57Vw3UoWTt5O+VMoVMU9ufnOSDQV0NtENBU9Qnkatib9/rCmOh4n9/GNfsNIPN/
xvboUwzcxXxEgvFd/win7/aykrYFRPFHypzYHB6Jz9NGFwKHdp4J/QuRkxKdOQ2ji+PzILOzoaQ0
0xoEaMzTfnfiuLPOgLCONCRMgIoTiR7r8MlBavTim8K2InmeY0coBe2g6Lye5fPFWDSnQDeKDom2
Qf9nnIDEiECqb7zDTACt7p6XIMnqyftgY7ySLDP8XPNawMJy3nOthNxRQfpwjWqYNFLsmmakgrdJ
radfLYmFERFYTakmBOdJqYCZDJxd2hORjhCUtbwcWkH6a71qP6sZF1o6ww0+K7SMrXPpamTA01jS
jYXnva1YDBV5OE2jIrizUkTSIklsWTAfeduY94AT/Vkn4Np7qRorjsgeRM6vWSgGZXfPWPTqJ0JA
ggPYGyU5xdDQv57lymUdcpA9d2TXsRWKHTEp2PGPU6DPze4nLzTtWrc8G9qVenLsY/E2kUA1YO8c
DzDBVNVGspr60OlHpTcOv31zQX9gj1br13wxpekipZmYFpH+A7ck2Tr74fU6BjAk7PJazjUTa8/r
BTAcKHM74E2h9pyeAAeWdv6wuXCT/9y9QfX5rPmKcjBssjEiUSahJCkOtrJEUpySmRq/AIH/lt6d
/wXg8Cuoao0DdBxtbAM+gn/mdkpij+6Ft8mziKJEsoRq3Sv7+tc+oW+716xwt4F1aVi9II+emZim
slmyvSd7+0/ovN3VvL7PQHMJ5dUzy8W2jmXWfTK4oZWuiyAXbisaqFIicUxJUKxZMhPVj7DBre7o
h6yZOJ+3ljzTRMXLMjAujEQL0lLhotDbkt7/V5kDGgP0rdJ2Frix/Buojz9MgpIAJV5JA4x66/NG
RpErEF3Et87HKclIMDCNvdNOt3PZiMTlXFu/gr6owDq0J8x3gZmZ+J46LbXEiu9JQXHD8arhQldD
aUAJD8knTG9W8bqTQzbB+yemzTqmK4MKjNjq5VRc4IFXdc9+u5UBPMPq2bBSE56725C07t6dD4DZ
qC6qrhIffMfYYehXlD0bgR0xBMixtblFA2UlFhBP32FptX2UivlUhgEBNiHFuXmJUAbJ4wUmr7DT
Gk3XXwSLrJ40YHkHm+IOsx6h6PnJ00PgznPwi72TBO1D3Hb4LJkR4IQahtkMhHzY7x0Ur98UTW8v
xufdy/mOlPlTcwFq6kke2Kyt8VO4448HF6vsfIDMsndYUMuXXCaWM4LSZlJj0Jk0gJqO2MXI8AM5
bMTSRZLEuSqsCGVO+MXSyudqzKdXJhClqoWp/gcwNgG2haZfWYDI/czQIPT11vDNgyY9uUBY8gO5
jYE5rPUq5EDpPL2J5wNjD/TaYfkcShvRKgTncK2yOnQcCXSkuYen5HOOgh/nukzyId3HIfPCT++c
5JFTHkZW+svgPb47HYVpjfrbOkfWB9POWKAlCvCjLcOGOna3SOHtdAp7ruFHWqEkMgJ2+rd+0M77
XEGVjn/eqwmlaT0KISVLU1SMQ/tTDDs36HGfsQeydS4kuAcdUCFa8fsCzNTGegT7dyGqJ5l9fCYj
nqkG/Ou1rk5v3f6oIW9e66rkPq+pun/v1INqeeKHC5Tx9Qf89edEiAgBHjnAOGoOT98MjAgvUdFh
o3ivZqeliPqcDth8F2pVyKMG3/m61d7XFkHVTsjtkkdf7pITXHvostlOiLxM27B5K/PTryYYnFmq
vEffBf0emziN6fuF9SaOiMQAuXcYJcmwomQqAUhSF6/8J1+HmD9wGxe7wyoWUGV7YSHBpH7ZK+H1
C0i8gm+mtxjHavyhuBjTXyXADeA1cE7VT7Zx5BzEidTZId3n7HYcOLJXsCSkDWXFE6Wrb9VwBXEz
0vcqnTXGCiO9xIPbwGNpMxvcqARsXSEHc2DexaWpDOaM2zYI+PSVuk3mnbKkZEOyUydin6fVtkJv
Gk+DwnJqiZOr01eCpTqdAxSM1Tty0JHWSKlavLtIQL72qYeSTjBMKs4ydokv8Etz1oyVqeFqdq0l
UiMx9Z/aHnFTQjmtssV9Iu6lnY/GGIRgWeYPN59pTYYm4Ay/PVOFpslYr1at0CqQkwE4RrDpwvnF
1HX8e2l0I/4tsABfxZ5I6Qk46PldM+utgE+Clv69jLLQwY0rLiAyRsOdYvE7gpE3mXIsXj5q6sGX
vZNtHaKQNNehqPpdT/uIhl0QQdxn52JKtaDnztofAOxjssWqK7vQE7q+cM9MsdiLUb9rQ7edMW4H
Awz08zmfw4TFMibg/Tj4Nb+PE730ARvkAX+EZvLVQyCkqdhPPk0DGjb7UL5nb4/24eXPlnTIjzPK
8bKNEbFFzxnIWs/193cNy6Hso1m+xko90hOdQ9It1qX9jlhEFAcVX9i9UAlBk+TKNjImpYF5vs8j
7e50jdkPYHhgDx48API6EJQNjeF8uHcNesw/KVcsq2BEFb6B5lpIdIxeYsxE0QRm+UifoIB6qT/1
0IXsjFI/zflzvYq/GYNZ/sYdrtWxpOQ+SsZ1zHk/hKukdC6dfffMeu55d4OcaG7yaAYVSHC7+Urn
Hra2T/1qBmSQwE3R/QZwUJ/dll9X/gwRtK0V0kgloN0PVRKQU3ZxNka5cC8b4XOhvtdbvxBbxxOZ
sNSHwFX4VNR9w5Yoc0YRTzCvVME+auh8y6WazjcYV+WGi+K1HbIiIysDJ82rBuIIbCtXxUv0M0dw
XfYmY53pv3gOvGa//9IeoD7PTT/DZ3FKn0znLrF4L4vemTS7CUQfD3d2NpsHI/UxW+SA/qE3Uxsa
Y2DDQ40FsTgsGs7lXg/PSXvSa4thd6GHMhsNGAansfWoCb3vCP5NPFb0P5wLzMCs7/uYXzk6wZRh
CUZklWDqH4fI9D8rxgR4JFWW8PEh9Vjqp3cqrmJ+9CKCpIhNWe5ihClORyVEJ0Wl4v+fq1l3Yf+s
E9N9dVs4A00isRey7JMlRbQnPH3tBLXhruno9K7DPeqJXZZ3BRu6wpXQh63gKdFaZ/gQE8hUcfc9
OQsPffhF+nPsylzVUzGkSRIavpM5SnfoMmU7ri1tHsTBeXcemt3olbrKy9kWHKHLrKwbsf+7kBK9
EPlN3uhXk1j0YpAf+y/kXCAKIa74+JAr6kYlPtOKcOxcybVuAdDZsJyXpUSGaqcMHh/Oh6Hgj5q+
Mipi2mKY1/CV0iaTfMjNBQwSOmGQNCzjZMbYzDmn6QNuxlwa/t961MmK1S1brkEh914pWZZS+wly
zLXAI6B7PncAYn7cPfLUSrqRbYWkI4MnVT+ip4fNzh4pbxrYw/z62HZ8TXHCbahBC3oWq3WOPi7g
wko3O+fMKM4X3Jawlox53fH9RoWlNmOW8wtZv/5mpYN4QsHsACpwhqmV2GivH/q//w2aMjFXnxW8
2HjaNUnpMshIwHwhhem+T35BHZiuNRKNOrYTfn07Vl37CrTOAi69cetFF6U9EfrJWB2fE3nTQ9RX
/SeXB9hD847EksQv1VAJgvWB3wouzOTe4LYzELie4Nx3AS6ZSe1c+zyaefY0vtgttMQsuq7oxWel
WPPG7mxOXGNTDHZpLUnc5PNOkeYj/g0H35TsjyvwfIU6/yPkjSPWCn3fvKdqM8y2HTQiymI/6dt8
mWHCbxeSsNx2JtPTBnw0sMJvl8yZqplrgdIS+0AyJcPDufZmKGtXBsSrvNTne+wEirV/hF8hyFVI
0eIBXsavICsM9senb/QTjiLAFc0MjuFHe0ZbigOeNcuNl75i0IEJ+03hGSJ27OIeC1g5DcSxQhgA
zZnyGyTd3ZMvnVXMF+yZSMhWvY3Zr7BpM4p5OoC2RAYawxUKZ/v/ePXy30kK8m7D/aUW4It4BuWt
u+DY/oBN4xw1Zy/X8KuoojvmtXTv7a5Ez3rcjHQmATNztI64sU8bGMVpJDEFv0Euy9xVYdLwQlds
Koe8AZ2nIXaUMHQAkhbi9bM+jEAq//tjNAT1LVX5Hyw4cUeMiXGHKR7FDs1CcxKNsGE2KxUSVPEC
uPJhF1qYb9v3RwYSQcDoSQQKSi9iLGDbBndJPUEF+rs6HeSy+Np3I5vwaJ42LRHguBj1a2igreo9
GRqDJQ/ugoN5pJurAurXDxkj0C67M3XRflSuESEO+mZZbQP4t6VJ4ZcvIvygHdCPc5F/0JMnHMEk
iIkxZW1ZVKnmKQ/yiBc6CKxeewxwAww27+v/P1alfv7zUvmHkt78EOLsXnCXEJyxxQ44ZEBmz27F
uFNdZzyLquLqPvsul1wBGmRiO6r19vTPqVLoVr5AldWFv8sfIzJz81K43LVXTfqRKJ4FZR1V3Y18
d2ndJaxfHWrQ2Ir729K862kQotCpQ/AEDQOPad1715AkOODooLL/r4rzgOoJD/a56lXNEkTbHAjO
hj/89Z3UBVMeGXBUMz1rOx5CCnExUdneIZydyxDGkpFNUXRMEqddTRuqXrjaa+RTZY8MJQZJkkgs
VBbdcV6ZTLNQkr71kj8MJ4PXYgJawvd3Ojpvu4Eaw4W9IgCUkaR5bfGWytiA4YyxFgo3u7azgPHI
bgcLEArhomJeH/KokEToTTNSoxRhaKD6MyRenZH6/AM4AkkAkogZNvtGoPV9xJ6lLx/V36vCUGau
m+DwcAyM/6Lp6EDUh0HRELC9nWlQrrdYTBWpjs3OgWDVmwcajYS28Zwb4dos4mZkxLBn6rVKJEli
W63ZQ3+xT9DWSS6c3kZxJt9YSKhzM1pjK7rTp3ptWRM3hl9ml7jqBndE8aa3jwwL0XgPFjgvMr+9
/SUzu10sA6KVRaYmSJiFisNHEHrtPLn9+gBhLiFtrfG42EOXyxKa9beEfCeUtvvB8+hABIi1FnYc
GZfoe4qJtYcpIRWGaQX1nA6u7tEoBmIRRwZ6/XuQDxqRqjzvXHJWsHM9xrRv/Ah1PXt+PkLcZy9j
P+CKTEd3U2GmpnMTy5N8tzk8YYjqNzpgrYOZyULeNpWLj/5LYms8KznYHcoj2oqZdJLJymOht8Fw
ZYXpBIHF0SN7ZlBKcUaXUs5f91CxmbalzvZXPd4CXQDK+vXi3cy8NzfK1GXmPtSjJm+6lFl69Kur
XS163LoZA3iyZIto3BaMEpPA76aMIZUV7JFQzrng+VmVxwzbakSL8z4wRlNbfzaUPifar7s12EuZ
L0sHRppSffuE+9U7Ut6p9udMlR2Y069MVQNkC6mhcfRB+SoBFl9KplyROny09c8C2asZYp2AVHVn
SA57bAo6RpzNDnvoSmITMmknmzBMNW+Z95zlcZHq3M9RUCvEdh/YYOoyB6Q3DYP+ZPm2L52DiAw1
fSyODnj0upw7wyic574bz4XRNUA7UhzXjWJiHC8/Xz1TJNHAyZiLvmcAzImsNsVc/l5IEY9OS4o3
DxHuC6HbDbA10sDLCti7NyYlM08t2EPEbqB/5J7F+ljBwtb/jqOPt1Gj0haJj7ew4O9Aj28Doiey
IcGJyFjcGOhi1GDojh3aEvF3ssVUqudPtQPu2VgpmQWxrfRZppdLTm9B9G2AaMTS/VMFi8XJWKtG
ibriRz/P6y/WkDoayiIEHMWObWivCQgqJIHuCLxjfr9vfWIHJnqaiAISZL0rn48x6DVQgOzAP5A7
2QlVd2C5Ch0/vsBBBOqHTucD7OIw4jHE97fOJ4uXiTUKHpFRzqfItHBpbHyDWvKhVjZ6qzy3lejY
TATuxcPIqfBCmtQ+/QG6UDfRuo5L8ZgNYZrlY5Xv9w20h+1HVUvSIQJsMi5krVdMZ7eu3z4RyjVP
+nqObZWK9wnySsfagmmLKhh4B2rcqS8XdmjKfuYU28hj5H8T3MKLxIVXSPh3PIDmCrdQ11QfvmTB
r7+G5ivUsrVLa4N8srhq8O2LCkjYYQmndCCA5L6LXMVIYo9RYTiQaKcBYR0nPQWfBGvoqNSD0+qh
uR8ZML1EKiDD9adX5rJaQPB3gJzB6oQCk+PNK4SlJjyX8a+2nP0QLBzBPM0ddc+KDUlWfGuwrsgT
ENiL5U/Bjvkcn3K7gNNn4vzdwoN/ihhWsEAoUUVoVGqQDiY0R8s5ZuYeJmz0mMgoAJs4qv4/TEcg
c6dnS+XvnO9Urp/uPb4Q4Q3GlFMVwRqVuCug9HHEqCpf9JaArOvFJPIcJQMGazJp1XzlZEVaQ7xt
V8x0EDnrT41OA0IW1cuVQlPyy9cRnnqcd6qpRwxaNAnzUKzH1O38GWtCM9MVdYyAYC0nNa/D2jJY
oL9HWzRqkTFhwXTAs37bfT0ZpxUECXtJOWCiduE+r1s2p32QwF4FQRqnf3WQFko2zAasxTHPb5ev
TooLC387wxqCBDMoDUHk9SBwM07z/68CnGBpMPOMv4yw44KMEoUBDfsgoas9y2O/w52iL4CS6DUr
aMNQ7QFe4qlVG26S/p4KAuS3fEXfPOyZgIbScJkxaXrSuvLkCZFc0GRTbkAlyPYnQQcesPyMPhhs
YcPwusDyI1U6o7avtCYaYcfSTiL5QTGyq7s9y+x4BBQHRS/VTS2bnjzz6rzcmg2qk2jYlHQ9msys
voX4RbyPeVRTGfsi2Sv8dxHXB7Fpc+1rk0OyjwZUIiEjNCadvr40JFyVKUl8vM6L6h9Gnhw7Oe0v
ynxeQMOgFbWVZyw27JNvgK0fV0jQVsQmQE/o37J4Ba+QRWZBMgvyy0CBh1QxG8+BDPjtPNq7rP0T
fWuTJd3v2p6nwDWZkcKyiChQzeU6wneMynUAbj7dkPwTqoPgdtBNTpRldaAsg1XR2moE02+MMlAX
v87CQKm7PgAtoDutdi53ydmfZ2rx5lbXnaaR6YMkkUHMimG2KMbMBHmTZLT4LnFsLy8hZcgkq1dE
WkCY/ScwJyFp7eTryGIhuaY1d0M4rqH6UgvYYLY4dOMaP7mfg2RHA0cu50TjrR5LBFVjM4aBDc2s
kBPYO/6vZePSwN78Vcr4EisrA19n9sORvm5kbYo7QAedfhJQZ2t/l5haHcxhWZ5XjnBkpIATXTvz
epZO4hD+52nNMXgs569OTg+qs5u01qGLsgPg8Um3DXvO3KU2+aGD3vOSOXDFiHYktjpFq60QB2Ka
/vpmisQII8gEl4jY6QArMY4JVTyIsio/JzCVSU1nes563k9r3dXOKuYhhEwhHa4kV5XM9Hsd5XWc
2uJga4Yekh8BjKcgx9uIrp+6y2FHJwARLp393shu49XN7CV2HDHYQVM2uHY4sBXLNhSFPIZIDUWA
CRAsk72gJa57cCPACuCwc7yW1/ny6yu8xZ052v08HYqFVRG4e037ukEeUY+X5GUaTgZfgaK69Qu8
Mf6D/TRb90GuW58QY6GRj+4Um+OQmPaVXGl+l+TDpRflM0wUU/Qo0iKirOICvs/0nVltCIsraiQG
XYqYYHQXj+xWfoWRVq+T8MNr9AjFOomc4vels+87rHoFj4MRYe7RYuDA4YmajuE+dtTZ4Ss+jF8w
s567c4aHkarta9Zz/z6iAGNf58UIwojHe872NEteCm9Wo9zc5L1dS6h6FOVXdxKniqoZCOJR2UlT
UfYtM64DJHPeJDuEiXnbtAgHL6+4mYDVHrQYOuuhv619MIyfoe1lLKhOZdCa4nIVId3PMXCaxul+
8VD5Dckrnfusx1pTExjRfWBitNKv+7K5QpaJDsllrwFq+oHYUUW8cyi/dt7NvSk/ypDkcIkusFpC
zFAAXLYZcnJ1CFyVUIaXPjiBEl2QKB6crjFy/GcVTsdcam0+573q18sxaZrXRaPQjvq/o8/iS9Kd
GeeRIuVCnWjtpeUiEVgAqRdCckg5tEiayYsNNJrM/2hg6nhR27+aOmc1B7L0Js4wAcmCglD4xW0t
S0ZUOh44fc3TK33PB6rVkwWz8A3BC582WqF6pnnddaQFal7htDCG2ma+1nUCUDDASfMxwq17h9BC
It48pYJWSv09Etu079ifkFyibEG+pUYTAKahbHGt6zuQhF7Hrv/LNx/4eBASIHgvo5tRo5AomfBW
hgTA4JO+Bc4IfmoOtIzBTYwDTIsy/nVwnktn+FFi5iTsDkLT8J1ZA4rbUV40cf+j92WCjxGWk1LY
JYuL3hn8NFmNc6ElEEKpw2r0cH+N766D/v+KqG1pYKAce9LAj6nyJNOa51kdG9QxPi/buzcQtE0m
yXmC9M5GzzTsdFceUR96OA3VtbJQ0H/F8ilJHT4/TILe/7HxTYb38/mWEl29/YdrvtxhTTw47Xix
LJE6Scozm0IKtJoGP6Emp9vHlnGJ43KGfpQsJFC9AsIyqEmrWcmuZIuurHwUTqFHs9U5S0TIzFTH
NmMxmOOkEj8g/RJxKY2cjVLeawIPniv28z8muiiXJol5AtY0VPoI9IGqzHnpNo3eVWuLBfiuZ0Th
9ynptPhWv9z6+f3DOz1vOMUxC9B/DSDjIIzY1SZlw7qUK+wIRNc6Aaw6pgzeygdWPrdmyhxbLeUR
b0LKQN+7tHxH94tWKAaVxDUlZcfFbxx+XEPe7uvLUrhfcStasZ2BNFuIeAmAAUw49uQP/EbvW3eJ
oBUsWug0aTCqGDfdiEd1Vu2Vu2491pKNC2AaNsBbnrDaaiZzkcZMtuVt9iO2Do9Ml5xATfYXxxSP
JGNeeCDlARMtzk9XdmT9rxRI52SHudCR8CTKdszynxFBPTpKFwob5ImqcfBoHvMQD/i6DDeBSiF8
xZzs6bQ8xf+vNBLSpDSIwu3LxW/uc9ww5sJvtQ4+yZ4ZBg0DiZG5VjRFlcrwNhzxppcsWo5Q8pGO
egMKpugF76zimsywRty4FRkHTC3Yq6cDUfTTQ6G2vGAKgiD2GW25D+3dHpf5Mi7lOj0wiuSVFwYC
YGK1cN6p+5lZydQrBtzNCKEU8PJjvGcz3R6cITKm4QTny8itxc+TkYOhiHB30/5Ez+j0h/ayd41l
h+w//L+AM0AN1JHiNT0XAXNtMjdnslw7o5kO7McqHw1RshSlOty6VhaF/myIpKcpOF1hBTZU+BFt
sVZZvAWVtSPY9JCcCJIOK2asIlrYVmHU7NGqWejbl1xt1aPN3GajrILiEml7bFi1v0+5D87VkQB8
jAohu5/TpXFLseC+X7q68ftzpFXb8wh3yOqV9OdPT0aFx8JRZo1tvNWqVABz97ugmPH394zAlGNY
y7gN+4lARPUyu6ZfYbNrgIPBcjY69XQHSv5RBikIsCZETIELIQP8QqjSG97rrGoDbwj7vjAqs6pc
DbzlNO1DK2kJWudN8oB7MlrORsGc9fFEZnPi8EUpXeTDk5TMizlmdNG0JQBrYITohhYyKy9q/Z04
4uXB+INFnUkyaNMSq0CwtCv5YyHmugij/slTzwq4G7qdrcuXzgYaGPZ/P86nBxPeO+/48ddZec12
sJVfftz/Bb/z7b2aGhFKy+Z0E29MZFW3TBJU0lLxQwlVS+1vH+g5Hrvt5TMyX00O9upbS2rt6RBo
Dxlt3+cGvfY613uBHj9qwL+t1x3dWUxaUNxdeNxMcBkJ7JtwMTdqo89mpu3+2nltYP08tn7VXb5N
h5Q6Q6dkK46RAzPTzL6MuKWYxEl1/QmjiDehAm1aaw2TiZB/tB1BOdh+xDS/aTV9a6vrNtIPJaP3
Z7b9etCKae0tKqinL1XurE2qPNl/73EFtzehLeMs3CGFvS2nxY0nncBXOIrYMyZ+oF94obGF2lH6
aZr2EehXD4Oqoc0qNyltmAX9H3YUUw/vWz5WKQ87Q9eGXMtXhq4h4ZdAp7C/6b3Pi6hNHZhg84kd
9OXj9oT1+d82zs0yDHrlPHxtfv8KM2LDKxDcNcXqzZ2oodY9hUf3LkN7GUrwUdoHMB67Bi+Cu3q9
glYwbS0c472P0RYxMDoRVxmTgbyS5JdqegsfXJJE8OH6NL3DomF0wIwGbweGOvCrpHq6yu54+Mb1
/Nk3ZEdLkgBVSZg51oBZyRV/C7Sv4O07hyRVYaPwa4ZmSKLrTDWEJV0yEC2k2JORXnoc1J+qsYIo
nwe1df2lqadjHChO8kwd68MIcSoNoaBhh2DNQQgm+1dEw7/ftmUa07Kkx4DD6e+tEl2rhk8e1UtQ
Y5V/YX8i3xJXXk8KzNLmO/EBgTXCPyPLehu+HuwLA5bbTibmCZyL2wcZ4JaQEWfsyByomNZnr0c4
ujBDTHlq+sLuiV6e6DM90d76egHV1qz9tvHG2Zgn5E7u1Rv0AaJaNrHL+VZHJjnvjdYE4CUfcjkX
h2ndSIZp1FI2ry+VSTqu03w9mDg0LPgE5nezXYYs68bNx6WyF7R9ANiPJXMAcS3OAUZkHbLwG+AX
PL1oEYYCuNc4Xo7sz9W7A1hwk5pHNAQwTuQ7PEaaBF5RLGaXo9p/qxWEuhMUOwrt4YFhZD0zbojH
kggeueBRRztlc4zSe68TmjBJBmx2Bahe144AigRXVL3vnM88u2WJC3WEERDHYw/LviPGcRgIGIIy
cPdAB1tzcmmVfLre8FVbwndVKj82+uaf13uweikhqKwSQRAuguXkXvYe0Yx2fICTXXX8Hpfvd8+S
rA28rcZVqLX/fjX53AquhbARuAt/iJWGbdaS38Xe7iXrlGKpxCwww2vY5Yx4GlTxKOenSgRvYthZ
LvVeZUVPxaDXVpOO5FrBwwc3lkSyITlvHBXBaPa1F0mJedXNqxhKHOaX8tgwusYnztAmw4UB0eZb
kXJPd7rhT+Iu1N6Jx6g5PF8YWIhZObPEZM84z6lPNctv66Pd4jS+9SAwUzQdZn8QIUZqF9tEvwzD
7+iFNhvbED7780YRr7hYWysBQ/1TOqzrN5dCTQxEMH7F6qUYJstqrNy3qBfw6dEjyvhCwnPM38zs
FyjQ8f8UYq+kYug6KoQXxVTmQEZYbR6zVOAgbWptqxaSRJax/ehNlBK2z9wP82umi/b7AlirQm8y
Xuf82qy5VIRddtvvcb62fe8rmwPWDCJ8vY9C73Vz2VlyDMg5Lcz+qKZ3mpvgRTTxXwayix83K7Fb
gy4428bpb2D5o7DQ1N0P90395L5uuTjlPIzWnr2zHhBip+b2Eb+OtUMAaS+s5rl7s2ekhGN39h6x
Ry+Xai5kPDzdpHS7xRcR3UnmZwU5/XwpMc4mhy+ufdb89KJX+mDRQgfvEV6DvhTLEMzrtVqdRT0R
FBIfuHLgkvNuA+fwk+FigLTqVrkLeIPIdygjTZY2k/0wugU8ugxC8s9QPUodmKLDPs2/71HDyP/1
a8x0N1PA2yAXL1kLGS1q0QH5h9nNmXDS7vbhCoO3UrCIRPONxDySxqc6JudJxFvbCjuSRWpMitWK
vLHd3wE0tTJqa3Yohk073pLRFgjUikDUWERJWU5LumuWoZ+eYyBc2m1mV5HhZ/dJ8TZXU1onlJ+W
kNWF3ZArBihohb5B9+BjsGvevmyJsCQbZjpmxEf/jaUY7nxirSsihHDHLq3IaiS7c/vrGVUnkkMv
Dtot1I/FJKp7vIyX5aibtA+WvqsAaK1QL9ujcRSCes0RvIKu4y8fCvhqOWkV9sfXai6/8BBAY3Ha
b3/nSq0W8VHRPl4wqU2L1adImOr4xyYF0ANt2muYy/irqGFDaEkpWGhdHGYvPOL2uNmjHYiNXXl7
hdi6w7sweEYuqB2CePIWLj0Esetq57OmM/MM3CfK8VgDU61LXWCr97ERLb8Z6gFjGp1dNjiU93zQ
h2j1YNjykGTiGS94X4ruI9AzMfHsazckjCfo8PKyWyYLdpyOwFAwEb33pIhw7IhnUC7fUylphSoR
AJ2qRR2usK1bJaY5xwdzIOW2dcFbbBMKuvaEl6bvu/nuLDLLxeYKVr0JoCUItFcYh5mD0VqJd4k8
SkKu3RpwU9w5cw/OiqFHTZlZLXuAZjMWXUMjIpNwikpxqW4ULdquLAuTfriiyMasph1J3VsHmWqr
rUrqEVIcDSRfl48T2KsD5QHS30q4TjQFNqGLucFqSgfvWVQm6HWI8zI0pap79iYZRiASwJx+MqOx
FKjZXnfe0g2TqBK+uTTq/lMFefBI3dxpXiGLlQaIAJkj3iYM+dw6xbxYsxefXStvhFi/WTxK6mqw
7W8i4z/kGLhLKJkPmHcHrP8Yzn89SSKiuZumBS52zN/+JbPZA1UE9lMzHxHFmyrZfAO3uuWRTh47
A29t2ir8rSF9r+ZsIrsZ3r2UfwgiMyay/QEAr26h/czD63CzHrWZiy62kcAsGZnQRUoDB5Hh+nIz
CoZrWNR5mZdAKAqYd84WjYrzSxR4zm2+MlFcc6tkyq64z+9Lse+GA0wnEAle9KK5Igsp/52D82k2
cFel6EaN+nF+UuU8/ZUuFOKK/Ef3lCnzAs7Nte8PEu5T/MGGALmMo59nUTVRLr1H1Px4fKRBNmIo
dDLI+j053UYGEqPwjgbmKI3njaIJnA9nPNTV5o96ygde2j7Rp/fr/ELLxdMiGkVgKNRsuT3kvJVl
UPgh1Hqbw+ujzmFrGP19mEdnitnC/3X90hlbdtnvyPFrKGuzu/ayQC8ImImOVP+ZEjoomo9y1Lu7
7ONBO2M/KG+sOMzUwvRcglo5Hyv10rvYw0tJCcyhk72ulKSJac/DHnDYzvVKWjOJw+wOs3AKhfo0
39SXt4AuyNN0co+nnJ2ENDkWXl5nFxniNmifyxwtGxXIg7doPKpjlU2SWBGYU/h7HyOzXO2+XzHM
pMjMzt2jxWC7FrXwMr5pzq/3mDKDQHJTBYBD7MyKsRTyoA/QTvbBsacr/jVQ2n+ZSDH2dHSubvM+
NP5+cNIYLmiTciSR+0gyGzvXcHm4o+nMquXo75f7HZBvP7noG1LJx4Ze9O7y5b+eHOUVidGAG4Xc
baBH2V+WFhCzKWK5GVj80soijZXToQ3cc7+UaqppOWiYi7zozFo5xLb6EcvI7iP6f89gX4eu0FDw
8Wl1qnr88n2LUb0aq3Ujy5JRg3hR094bVTnrNin67UXiVJBNWqY6uFySVlb3S9yiUmTRdlKPrVmf
drdQRAY+ZZZ5k4lTOP4vUn12eKZzcaKXKR1yBAbxdFYyKiuxzlWMiO6W6wdSCEnvsB1L7oC6a9FS
+WQIE+rXMfkUJR7mmBv/hprH13NqRLKvyeF8hws+pIDlbP/xyqz33QmueHgp8Mnn6zasBn2v7SZZ
TlUDGZdkDyY2/MzezrCrtkRdTXATonytSz9R5Qudo8p5gAn0RO/uCnA5W7wtH4k45VpBXQfVqsJr
SRTXk/XB9oDqqT0KG0vu3nPKRXVs8qsrkXmrvMPtwInau6z58QbhKjFzeDJONuTKDKAvIkUFiaAQ
tOEA9Bjgi+evH+CyDhvPtq/7IsBjXlEupqmEbaQoNe78tb0OZsT3Gd7lpouIj/ONK9tKZJ3K0B+n
6NZW++KiMJzdA+eRy4imPWcnDhDK7m9Fv8Yean3vwuW6ScTH0fb6HmTFjGcazPw5dtCgowbtpfwG
XrqHaxoDv+yZxLizH8TQkIkir6LvUuxfpIOo7dANL5WoFdbIDtJwgoZ9go9GDO/enpc4QkOABXLv
Os43Ch2BwPKxxJbhhuppzFZPvmQzSWctNJRNNq7TT9ue10CDGQHW2QN6FXQPRY07GlaTc7bZ0Fx7
BYpm4wKEHIvNxkBQ1MxkUsIWp2I1Y6VogWfmtecSC/d3KHN+K5PUjRXLH+yVpY8NqhG8FSKl6rZn
8eRvzwQfgHQHAxZdLv8D9YLxxLmJZg/HVBu+0+o0JyobN1AzfagiW9rCr/KQ3nffmlf2+skze20Q
+U1VehX2/OGI/+2bMycH8qO37SQJwFA1cCFKo82pEp4dOEKW19GocHBVdp+YAQblXz63YlUGaA8W
X4z+wHD201+2WSf+SHiOkFgmX9J8RAOSo9btNZk03F2DIVkHNAmu3hoySwq03EjCoaGD1DznenEN
3IE99VYDaDZPvKrEciTBhZSmaAldjSRPNeJ9QmcIYL8CXuD5FRLTcXKzdmO1ENjCTMaXcb5Zqf6K
iAIiuHN7OstiHtkC2OPsqc9KPKY2HJ6Z0U1XgJO5rPoDVcz0nCUKfXwlZXcC67PZlxIzbj4lj23q
DlZU4naEX3WOT8itYAVKkh+PnxP7m+WkTO87p5MD3W6++8AqmJQJ3KNUqlfXpPH/jKD/eJq9JpnM
0X0Fake9PVvF4OoYC/dWKcJjAvgTm9QdAbctneVFxEwMt3jXb9C1m/3prGSZ9db7mE952VL2Qi3z
QL3Ldq2LqNdOCdtdceNzOJVogbAwMK0RDcCE3nHKRvNTssiS8QSnbsKwA0BaVZK2gHyHlwQf48NA
9pERXLdsaU1yxgF6Tr+k2AhqvQGwvck4txK6YFnenvV/X6aIqR3r2SMpmW5x6dhbFVgzbBc4Cy4/
HZp6iEzHglTLBkJUC0GnsY/XhPlZ697mmxFowlhWfFGipCvjDo5kYUrFm1Z4KI4wkmqsDMarq9D7
6nfFd9CPZVYCLjIqg/Ix6FvmOhH1Pi68RrunrVp9Y0FGMd3CZCpCvZdereS52v7yjdqH1LtkIkXN
W70aPp6+7E9uF+uGLKumMVPPLZmY0Lqoj+NeBBThKqTwa53Ci1fBzDrXdk2s6Mt4c+uoJ2XFIoE2
wZjTLomUNQP7zzn6xXEZFpo6XCbbiQKUB+pFgNKN2bnZG9jsLYd9CIP7bxWZYRF8G+kModEhdRaH
OtY6cXUIsqs8Usz5rCD3Vpq+BGh35ArjTCSL39qyavRCaBblWSr8D1VGeh7V8P6Y604IPcpeQNa+
KHHHW5Slh+ltAuL6rA6R/PKSZe0Nl6D9i/sMUC73bPMmU2mv6Of2YRgeqKS4q1FsBpqLAdksRw6V
oDZ/cC+EN/J8rfB7vMVs9Whe327MffkRU5Ojp1z2rCePQysPc/T2+H84/mz8gekU8TR/FnOgHNPG
+cZTB8CGpiMYBaWVYdi7rQVAYuYR9wSl0Kw+9p2m6m58gpcanPM0zN27MJX/suN14gkUulTuEL/G
hG6kYr+OKp18mHU6KtwMnAXlHx1v3ms7gsOUjNmnMfoiATohz0osLrdg02RrQqEBN43tWJ97+Qkk
Y3lOY3vNA6FM0Xh8+FVKEFAR/85bPf9LobNbx4+/dzJrOpSdX8bY+gXgFTSbHudgjPk4FnrSb0Mo
76C20us9CDF9wm2MMtltbAjCWF8XThN6JMkt0PIdFf7fQ7dUC4Azvc2/ZcXkHawBHRkJur9gAMuf
utx/H4tXOcZEHvFZnteqmTZkFt/3VbTEq7OwWgUsvCGdq+DxMx8RIPmro1u/3YfwNzzhDoUXP9Jj
wJgYG8GdzmiXbbj40PX1vos16HhPLqbJU3tW1DvuX5w9oBOUnJRfjgHgesyNZxXycTLZsZiZ5I+i
h/3s6TRjjkDBSG2WRvO6h0f1yR9b3Kf81FftfTKAeOlCA0q60UsNSiv86WP5vWGNYxKXWDK22DAl
p3/u3h0njWOpuRcph3EMLL43c+Zh2J3DTjGxljWYFxfAwnRVzvMsDu7aQvF6HRT004G+kd0o5zGO
P0HBTIscMwK/kkvEtbTdeQnx652fDWpFJH9KD5Lb+qNos6461CK4fl5hoNCGHKGovBEPLZoIAN+s
/uZZ1xk/6kjqn2n9pt9OwteC4XLdCFJDulG8ReDcBDY0rmDqqVUgGfBgigyPnO04h4LpAnFMXABZ
1YNKj+G6aAVdVxyq3ywQO7tE+8HJPhjFssTcxpM88r1m0Cw+SHisPfUmzv0opE6WwBS06tfwFgKF
MTvJ2jXSj68ExKd1KhhozXuFMBrhsBDiUIXc6GS5UmdCDcVcQ2tZIQVOm5G214Qn2fI/x2+ol5Qp
dLboHFkRl/s1YOmFVtW2wnTgDIfMu17x0pVdZZRRcSXUxI4Oz10fqkpEeuvpI6Q0jL/O6NVTDGZk
GUNovojJJAVDrQuMi5arXU32RS2SfJTICfdIVds0suFi9YtknyfyvGnVot7FYy7gUjP2RuGARoN3
M7aEN5MHfQsWQemfQmXa3ZLhlOLr5Mz7uQ7WKWUc18FbTrNw1wx395tr7PfBeUmi97I8UOe2WvTv
jp3Dtru9rIkZWIgEaO6Gq6kGKcXDOKzz6WUCZGGux5NTSNWeRxLRTNiiWYwGVdhVzVQVVVEhGF6i
QIu4XjYKIhoh0EBxMm66q4Bt0ZvOROHwwVOuYSGglMXdUEwPZvc5FfwJT/Qe98x926Ik+FlkuQiK
AzhQ9gnKnQkowRP75i5bXHezfLM7FDvamGNc/Nyt6Mc7yjr2d2UgYF4VSd8R/DNUuT6uUG7OFH2k
cmUmx31pG7XuztqmqfFXi0B+H03zSUW9s0/UpWzuNSX+LN2QFcBg4JMP3flzz8ElNF4jD8zpUR2c
nx9CDrSyc0/NvXoI0of0OjvMoVPyJ9Eh+M2R3LF/Ubt/aNHI8g3409C5iUqhSECn/mSsg6qNqeYO
D91T62HNpFw1y7OfWc8DQb6Lwg92HXXbEKWmmczEW/4RL4mqsarnwmYCQb/6Ce6NjgeiE/9uWGss
8GtTLv+uNhT7UT1byv66vJFsrDBrSQJG0h9kj1dZMlC6hIwDWuXxrxRcPINWJz4XUtTZnzKR0OWZ
LQMI1QoNV5hTT+UXQtsPX59Z28Hnpmzg2WI/axkT1okIaPJUz3SCoEWsFeqqz5nio+Px0Nw1oGuk
fA+U/DhJSXGnthPPXELeKbVopJ3lT4E1vzLHGu5GHHiYDX08xVPJyd0WT+hYkTErapt4gpI/uOK3
keeIIYA6RkpQ6oA5pW05LkRzFaG1dYvttcWGhQcx28tmEE08tF+tnV+D9bjd7mPxZ4v7zLIqjNRL
rPyW4rb3UaoCxS4bhW5ZZ9h3yJBuJyFf28Vixl9FZztdAa/T54iaTQE166fg0tQy0trtAYEoYdx9
Wh2NpxMCkSBDVA3D++ROfkjksqEiKxLFF4JnjG/R4bIHTBPhi++mBZ3vge7wuRa2UdvGu+E82kBV
9wmRpaprA2n7DM3KwzCCtDBzpYnASWlK0lU/dctFYUBD+wjV4ViVlqeOYSFCOGnML7tV0OuSlwON
+eEQrsoDu2fG4tAws8uazxK6PElEh1ywb7SsOY2zo8oauaP1bC2U5QEwiFkBHLVl7Ew+LVuRe+YK
BifX6Ehwm8QxaYh+YN1qxetos+le6Q4ESVZdDIdGHnQDL39rj1D4la6WOe9olhh5Q4vBv7S3azxj
9HtnCFQbh7+JUvtpBhiOJKcuR1u9mrlNOk7k0i/nVND/4/PvKX/qiRbyeLpQDkbe21DlfdMazkT1
+GCfVAgPCU/zNWys76YVMNdFd0fQFsC5P5kxzp3b6UyZMvyHSfJJ28+gAkLb5B3zEUYN31srUGFo
idMH+a7db5+cEZ5/2PB3Nvdl4YhmzOmOnBSvnW+MnUb5ikN6X+WJ6vIgYQ+zUYWi0r/5ytUxtMqi
LTIlb0PJHSRpJTtEv/NskYBP+vW7nCWurApdHySBmZ2tCWy8ygQ0+AHcKMQsgT2NliwPoe4qmgxK
WiUL1F9lOJfmmfowIXrzL9Bm7ibgMpQ0yvybwS1ZJKEDwfwxQiximFSHdcYOa8Ot2voXU8CMcq8E
9TU2bTpgiIVVvF7uodWC8Xb9nPsCkOld0nOm2OsA7zA03aMTGGqOU7bTjp8S2dXFRziZ2R1tCzWj
+qsdLRntK9R2iQMgcz0mYemFfhB2d7UDp5H3hmYdJe0oEYmNYTvFMKVMmFdP6Fo6SDdbr1EfAG2T
vc1xXBx7WgCoSAC4rFazuAx8YWR5eOHtt1iupGjK2midwrddGY7R7sPhUcIf6pF9wtP0PSjVW6B7
dLnI3Gu3QCX5NmN3950Ousx9YaEPnMzxYQVLHerdX9Xw+A0cWC5jqVpwHsV4Olu4XKxT5+2uhdSA
xsXem/ARsOTTOJ2IkH6Pp74UKD01D94fahHrA3P1LKEm8Ty+Qt70kpvVIpovU7P+4z6JAWdauOJU
Sp7o5Z74KHK4Dl7G3eGy8ytk7WHneX3JVMBZx9a8riI3MogNtAzVtjToPUhvrhQcXjNHmZc8VUqL
cn/xVvlkbmKKlrLIZp9m7V1665odw/2VWey/JDBjn6X39SSNgO94xUm+g1HzDehvUpUFrk14DiL9
Po2yT2EL+HtXOgJecaTaXb61H34LfwU7Yitf/U7u9AfUOx0xMZnmPcudXNAKumGmXT6DDTGk7G6Q
wAyQouDurTvyyNorWL+OqlHpRg+J2MXQWvkAHJi/0eHJGwqJY60nzbR3wkf9UHXjnOZIw/IhbyqQ
XfHI9Rmf08+VuXviQ2XliGmxZXVeFCoe/hjgpG01c/J5U/89zY9pOlCWonUzmvB/Fp9sCCDJu6xm
4Cb1marPeVRmw+W/8erD+zefb1rdJaJaPCNwuAJ+wEUmkV+38J3mcHdNYOQn6TXDRt1MOgV5aw0W
IjCAZ1ZH8OO8qITgM0f9FddBwSE1aHndT++G0H2owW1fDGxZqFmb30t5Dzr6FZcXFyQ0XCZGj9bI
HEmiqhN1CutNqRYX9ZPpobFvsl3XQX1qTaAUMF/wBWsEUYhqQ2cZjcc6nR0G9Y/1DM5Qgn7cFSit
aYnO4nuQxM1NJuZRh5RCSXe2TE0oHoY6s3Mpmnw0qiVeEUVcVPewDq2mZTWHkw8AIH0jvMcJnXA8
tbLdQRsahht/TzkxueQBtWnTblfEKP60xaRaZ94nLOuf6lg+fjuaDfL+xfsYzoG4nPKpkPcR53Cf
xDQBeq7iBEKePnxAZ9hsF/qhxyY/EbIxyNG6pEaMkpF+HBjGtcLcpFPdHhBLBkBog/5k7DBW8IAY
zAo4n2OnMI/MoZT7Sv07tV/lmFvnlZR2CeNhA+vuyDzdXAJbt+DszQo/0esPPmUsqFkzf4B4ILTK
NKwTs7cpr/wVgztseKcsvVK4O+ga5eeRAA8oI7AbvuHvXnMH/bA2zm3FHm0qk0ciRa5NKylGOLIY
xa9YLyuH0j48O+jtBqskX4XSx5NeyMj7wkXnQrCwWqCb0pY26/m45zvIdbaIUtguueTIXVmQeCaT
PpKIdJqphreTrSFrHuFvK7sHl8ct8v44909+9Q4C4qVzvja/2RVk04vIwWZfC18jUfgynUEGeba/
89FvYaXe0jPJrVAywksEujUqU84Gpa+395Nalj1ZY9DOq4m5DmjPzZ7ZXu98i74g1V0ewrJflqg/
YrwpyZsC9bVb4g+cEWpQsTbVdFee+w5ujwc+F3Ap0l4xJjpht4iflJwXvZwfJoDiZvImQS/r5RYm
6VGMUSOFd4+LNB9m2/UdKN/aauncdgEu9eLUyD7oHGzqlFmtxXO8tDHk4p2bPSOT2Dex9+46LtDp
zPSYItAm1JMFGLcMhPuU3cf32ASdofL5dMOsZsSpteV2fVVvKdXFf/sDl2emG4tKuO02/RY87ocD
xIbTC3ugNND/ZNNpvFlP8L5S62DxH/o10XDj3pJAPWJDIrv2E5dcfGV0DadduG1s0ySVR+0poj4O
4GUuHa+BKbCR1cEoQzrUaVZV+oL7YH3TcTqD5OZQADNHPYuD/sRJipmNA/AB9oP9Mv5KNnOAalsD
tS5obc49HarXWCdFLfR/q2x6m5+Hk8l9w4/cKzsq2uEkaEu0xXr1ls7P2UVmrHXrk7QtVIK5m/NR
EOFlpAQFxhvWPJNBkds69QAgYHJAk4Hb6PX1yN3acgAnWhe/G5WE1Wxtzn/Bj4aeEbLpboo6z90x
GrVA+qpEltFbRXdcfEsc0x7E4pqKkyiRRNF3RpvutFEVm1M3aGT9doGYLCFWsTgasl4t1uviZ2Dh
nUP8PVRA2o7DOdqfMEnrNAlVicrBDasM1Xt64/MEU64cGsiu0X8MPKSnoLc5+dppCkV/as4RxalJ
g5QUDUA3JrahsGeugjcX+VSCrouxfs6BB5wOJzJ+Iyzdti/4kI2HytP3MCsb/Bd+pRwdb1BF/ksG
0TMeaBxahS81Zudvcu/usWKUCkYR1LE3hseyaVbFew7GsnS0jwMwEfYQW9MQx5xYthf8/yCYgxBP
2DeSaq9Fjo6vHhKQjT5PTJe6OY18dUcFmOVhxN0GzD25XCrtBHtKHurstHWw8rWMOwGEGsf1KWWb
q/Vb7eK2a2ruu6mVRm2BxC0Ke2fS5Kp+4v4DnR4bPfpasOGKPGEkjqhas06axBNPtNZETZnqTLH8
TcqgmbjipD8WHoecpaP557v6FC6llDdG2qYRuKG8HB+om5dpxnXxIwsJaSRotjsxWNLd3afzlwUA
YFtxFe8NhpW/7gtVLeDLGu+deGAZ8M84TnbjLUnnwZ4x+WltQZr5NesSt5UuzgOUI5CoUat7a9GE
tcETb6LkzBLj0UcSvS1O2VfqaioQdmKKgdtOOlEbgNjzGARIOtr1xP+e8UZO+nP6yua81EFrfaFr
4uEUM15pzm+c8ac+qqR3VlMD261Vs3mqQ1yT1kU6C2d5Q/bitKGfMBpW9wMqROgcb/LLeqfCOy8W
s2gcwcutXHKoNKdhF6XbKnZvj+RxFdKkkLx7b5q3veAjm2ROIhdvxeeTMw6aSLKTzKOUEp0lcrkW
p7C9jr7Q77Ae5HX7I9FUxi9pplNp7s8Ne/gnPc5052LHtsB8t+HJQ1OW2BarDy1pWS6ZE7wKKFA+
I3EgfGb6p/oiiuujDhu4HXJk/1ETz0RaPTSoa7CqNWMVgyfpKgyMITBTYrAeH2A/1oERtEBN9NxV
USUPWbFz36xt1cvVqlhhPN2THmV+GULKDpgijEIoujPAPuqMZrzbuJP6y+Hl5guROt+AV/5v21sw
8B8w/OUtOCHrF5nxUxaq7adeTTLC0hc70YRah66Y05e9YnzevwjUQu9rCZ9zlVVI9eMjPbaJpixy
WYJhSEqvlwdk8lfPMUnG/Skv4G7GOqnUgXXC9Y1hKPeAauK9Moqf5DRewcnuG0uzqV6KWf2lCdgp
+Tx5iHHuKz9Zu5Au6Vmch3BY5H/QVDq6xUmdVt5aAuD5AebMLD1ipL6ka9UQJQsjITGyqxa2UXCG
GfGbMwMZ1ZBpnfD8G1hMicNkG7U1Rn/JFQN5URZ5FFmyoTDCrn4m8mMMFnUR5OK6wclpcL+Ie93H
Gk5/NHwTTaNmUafNSk2Wwoh1ojWd5tIvs4r1a1WIamAH7Zoghudt640xqg5csv7t0vXqyIheuTH1
F95696fksRwHxPgw5OSO/YjteLt1utyENa14+HzC6/Kn8KjNVpRRFj95FMJUzVkMEh6AOPlrIP1Q
g7NfffuLyKxiq0T0sZvfFhxh0xBougtKHYA0jRzoQRcNVGRx1bIy9pkfYmblFrXVEyBqMI6BYoBN
JbKt7E3uxoMKQ52XCQOFZDZZfU10isJXJjtqZWRkYhXiKGmpQwdh3Rn+X1tB4o9owGRg9WBxuqSs
qWeoGarpPoh9gF21+Sl0B3Rr2kDA6gt1PlNSZaqGC/yRlc7cEpnElBVuUCEXQhRLidGBYrPelqL4
0ikvDfCuK73I/YeCog9XmfcGIhg1W2Onoc5QWEQme1od4go5l0hHh0NhPDymilCQbiBqU67c2LzH
WTzpABmXdznGA+4rf0OQALQsg20bjdR0dTHRoLp6fGx8X2vZYRd5K64pDhC6ZDhaJCfZdTU3W69u
yle+tab2aw6RgzUd5ha549CLdU9u7u9/8DA2UNzdLfa8f4F0F80YLyqcejZ4mKc6+S7pbZBtUZBS
H4rS77MoAie6gBzs7TvdScTsQAldcONO3QGnYQWybBgyjjqAQPeZBvCAlhYyGY91du2ePpKX3IIX
gnTXOQAOaSHaTO8h0LsnphEPrFkfBm/b/fqmSwnueyTDcag6b+jfvlnKpmUfKaJkOH7ZHhDQQXHe
VMad8NQM6pU74rldK3djWvQH6RzK877Rpov6zCAalMjcEtG67iNelz/mDfPAwcMwKhXDg3j1HWOT
i8zUlsyVbZAp+SBW/T1hyme5HTn2aaCJwstp4sp2ZfMce2XCAua2KevN+qLOv1FhFNwD+D7twMDN
qGtPXs3HkjQDQ3Vrd2IMpcas4xm/9T2cuLTqCqvK2DKZgF+3Kw3fv5Fsr4nRsivv6mJR5J5vZOhm
hxgPI3effB/clci36TntyxOXCwjWt58d0h2ee7qKbjVhFYDTD6ePFeXyRyYxdBfq/J/Je/I5GUGl
7I2rq7PD79ZHl7xmyIqRbA/ydb55lYP6FpjpdTxRwT8pWFEPqPV9af6ONu+GtXIBWikAdIfDNIQG
BJz07bzTp2KkQv+dgmYjzef4/JdIgcj58zalNKtR3URNip+bkOlz1VRs9qMt10LdhwZ899Eh4sGY
T6XRuibvYBGwY5pPoW3OSNr8l+H9SWn5ZchMHQC898q+BL8oewuBuow67lWMGRyX0vnor43Kov/u
enoncXPKBdMEUxnn6oePIVMbYdwky0evDOBzuykXFOXDTQGCTFdzUckXR3wfUcec1MLSkj9Du+To
rx8okQjGPXm/C5ORg35QO3kxw2IpvQhQIC2oMrXbDgXxU4BxTh78z+R/jfhMpqrb+FBWw5b716Yb
mfF5Ut2qG5LgeF4Pnt7/6AtLmqDjTAGaZmgqFB85nUr8+KGufPOvk263V8SsKmL5Wugrpv9D0cnF
agXzeilzbQmCAvLInEIRBHq4wiKxPWS1iBqmoKSTHL2MrQgPdMoYdAeMRJTa+hY3avrPuCb5/aJG
r+WNWTW4LC4T6k2wzjLhWKlLSM0aAIHlCI/a+HjPWmsoD9gezqufQqxCHIkeXbG9pk58Yd9FKX7A
x6OJufqCuIWmPEangBdQ8RVjb7+ZNal0Yhryuze9i3b9UHsn4s3D1ixQEcciBJ7au16d/ziOJqfs
CymY2fbiTHTNjxmItjG7y3eWrZawR7D2/Y+pcV/2qCYPlgh915D5aCpx2XDic/xyJr+ps4Aqb+Hp
4q9t1ftmDEkM7lE8NYCSBfhWDSeSrucxi21oWMrnthNcJbcDfuGeSSyQmGfO3h16emmJexXP/VC7
eKyKXp6WDTci6xvw/WAvMkQmqrrwsmf7qBpV0o+a4nhADRko06pRhfokGuBMR/lCwvccomMwVj5K
VFStL36z/hxM2DNwPyLvF/O/lpbN9pln3wyrOToBQPFYtMwg5+pniYV/7hQT/Vt0lg5KM1trfhyH
MFUiohHxikDEQK8uY+KPoIgEFS7pO27J12OYcO0tiEV5rRNbDflYnDj32+wJmifNpnhJk/P41MnU
I8Kok/7ah53jVq17GPOmVtmstYJn4uEhLsvOj153PmNrFNa8wNuz2nWnBe1rrs3WKXixvidNcCuJ
p4cl6GgMsMoubbYSY3d2gznATRszIJKp3RN34Yjupwvhc06KzbGdS2jlyoRMV7ZBh3ZpLlJyB0lq
RnygVgz5kVvso+KJKIAheq5Hdh+OfGLPvXzskgNOHg5EUQnTbUvNa7KrxRLhJwIky+7zT02QxDld
OemMyQv5lg94ZNy3sjOIemnS2tuK8yjcidTU2otlKehvQx67/EIMHstdEKgGSIVKPIlZta7I44fE
iEoJqJIIk4unu26+ic4iKl2LQ4m5QH8dN/smofOAo6eR70aU6WxPOGQym4qYN3Tg+ugvWCy42ZEJ
WZHDlOwVjDaa33qX0V+z0jXr5iibQiHatcfyKp57dS8upOUlcn59YahjP21IuV4ocuIF/WxoHvQr
/F7FXVXxofQijTV1VtyYBIHgawbY2lSK7jvsmHRjSVnjPeRUpk7dT5+r//LecghR9dZlM4fo4a5j
K9K1UVfkLpyqjIUWv+JE11lQ1o1NQL+rKK/1207jCo+o7gzmUBpAW2KObiCzuWKUGsmuwAlhY4SO
+9U4AT4jcOwD9OrD28pWKDXdel9wVcung5P1Ir5uoDNg+QjFVXaLlwVKMMENA0vzxCA/4wD8cAWk
GekjG2XPdh+75GZ3Xoq4Ya0N6MB4zdUcgSswNPzc1TNnpAO0mRMJAmrVqAEY+fTOeSFW/P23uWs+
i9jtic/3XgkUKfh5Yc6AaduD+SJfw55A/8PXEkzfmDFuGBk5ZGEifPzks9ducvcFmjnlJM4XNaS2
SjRvrHRqcvhd9F2F1IA/kljmOpfmWJOxvf84lK8BeOycLw17fdVt+f2mM1zPjoRmgvxHrwIT/8KW
jHSPgzEo6pvNEuh3n+ADBxI0Qn+zBYoBleSKs7wdH6ckT5minNDN0kT0KbZnUpZ77+IkkFsTIBs2
IV3EvTKhoWDQBTVwwKzQhFZhh1/vEiLdNj+EuUqw/uQd517MPz/iSKej+wOOPLq334uSx+SV5PWo
8JqvK237c0MrhF+SV+GlaUKmBIs9STLHY1IZ04YWOGh8Ue+gYmbmFXJHP+EYpN+oDh11MOcjMAfF
o2WfKQ+bW8UXB1HcLL4lnnf8bKvuDUPVTiKjLhRS+6A+hZ8vVDo9wOLNDVsgRH5oYT7NzTIUtaLx
ArOPqk7uv4cbdpucK6vDRKzJTkHhzcTivPWi+3rU61FHeHqkhLbv3Psme1pvjaG1CosXWXRJigce
aEc+ldkgK8VmP4DfjYZyPHdJyYcf7cD4d6B+bNAgI9Jab8BFz+mrAoOQb2M/EpcJJ16KArSI6kjN
VSjYtS3C+AM0ydFz08XyI9LlcDwXrZnX6PMiFx++2N8f+IKa3CsUVBIEqfa4+WHfOOVpIfKgaUPG
xmduZUjue+EoZMVXVOx8y38l4b89jeKCrZcIuCDulH+F0cFl1snLbvx8hi8pxWbbP7hdALJ98jGb
MeZ7I8yTVQgtM4iUJPavc44ILlDNEXzw84KjFHaALph6uTRo5ewI1C84EMDwbiy3CmvN3m8JiM1z
gVmSGOgeg495y04iO71EGCMx8qSIag+U3jiGG99LfEgW3r4SfvDtLFjHpaF9uK8d/l3Hb0CPAaOM
OVKfhZT1v2wcVTwKkWue5DC2gNnTuodcpCEyR+qKOLyhnHDlcXDMGWSByQy2LJrK1+otJ2k9uKSQ
lpdfvvibxaYPWROnraO/D6+9wVzMDasHPbvtpbRmlCuO92ncIs7kv0Mvce3JuIJ/IbO+ATVSPjv4
/3nJVlp1X1xS853PE/HJS5DjdTYvTef1rrWAyadGMUcZ+32R921WAYrr5h7ZLuFsz2hZ5OXO2Iob
eAXfcKEquNYvHCMOjU/rxj+fMBKBwriS21JwtgLubm8ZAhcJ0C7SZskbTWFu5a8naWACycr6iJsH
KxH47ExaTcb0/e+IBinZ7pREqx4TdME8mirjSKMqcgvV72pk9mZ5L3I4l5+tXVeiuMl83C8yBz51
QFtG/Omi0wrtgQvcxPSSSbsKHZWC5zA8UFb5rACLHqBN/wMQXKVzl9b+cB9mDiyRK4hgOfFiTlhc
PwCP1cpXUYHnOVxmYKg94IP7ASTDuS3Ai8SPm/VplLtlsdOoUFRUlOOZ7rrftLRpqn4z+UuAGavp
fmZ5OZfi0wC2Q+cq4msXpYfeOWmfiJaxTbwGgER18W6oVKcE+7hHU8lEg2dwEzzkfvtBxG4AzfBo
dfmHaejQuJyNNQhk5C+jQWcT4rG4i03zslV+Dly5ceTP7aD0GH8NMWnOUyglRwhIjjwqfjqIG6iS
6wd7huZXrS6T95joXhzKk5G8fOFLycx0dY+p1Wi8ztBnMTR1Ju55esr2h8AOMDMfIg6kbNwKM2QV
7g3L208LskLOgUohrIIyUl2+h8Ofl0F9sPKIDKlSQP0p2E62DmLtFrG/HRPseLrXjb9G4FJ1M+m+
3++NR5La2rcm4VJz86yKDv/66VolwDD9+sUJyf6QwZ1c/RZxCVQ5VptESIhwpbgSX6kMXVHJuPne
V88PodM2cBXUh9nYFNaO2pPGJX3TzimMwxll97MiH1emMVYpP8obLkXYz+7R5Amv23Z3xiykcn4/
ocml9dwSeCikHHqs0/Pg1fNFF2N2/O5B/bsxTEerxUSNe/H2nRZIEC0O7ZeOYWkEnj5GV9kdVdrE
hn5alq12zsiau+lOILi6K0Fu80+1drsLaNoUrLdch/CxKaxhyTZ3/YHQS/U+n1UEM2JBtDByKMqg
WbJXSIZcNqgb0InBQeGsy3xayKQSSKNsddciIjLPj99jQXA/xMvqY/26ZDIBEUABlosD0RnGxKhn
AjPlI30jieCT7oalzwobVx+VFaSX3ATNwYGN/wyujiTgCJxjSaKJRvQxga3tx4Dz0oFUfHuPH1BX
HHlDzXlNSo4UBxngMEAvkN6cuE/hwwQEIs5Nw0LbaMztK2yXwPyOrvW+RxnAjJO5IaxCph/JGeFQ
EtPi79h4zn4C9NLIjagZ+TItSMD3ddgqfh941t/Q0wmBJte6Qh4ObwlqkrfdcQWfjBdRGeOWLSgS
NblZVyXoJyCad8INbRk3qVpHh5VNTmqw+HULqqVae1+rR+i+G4yXEE9dvMYZCtW47oBCJhvaz0wN
2cR5Kzd62QOhvzREsqpjeYFJZP6MJoUP6mobv9n6r8B7cE6YA+lRQnQWk/jKpvavKVEtO19SRFe3
A2MhZDp+PJI1tVWqudbZfU61nNq9NikuSyXKVv2DVA2qZ/IwFdS98fhOyDrElaOcN3BY8JVkZRgJ
6OG5o0DYQUxbmlw6IaMYyYCkL48oWQg3fWlq3+jIDjdc0t0su27GoAuj/6GJso8fwm0Di9Az9ACt
lZsIpLr1ereypuBXmKhxbH5djqtWYue3o475coBkZRiNiz5ySKFpijcP2rlWt/hL//J25EyYxfik
2Mme9YLFTV2RXLmfAw1eHyJoYm4FS0G6M2/uzlgMSK3ksKoDADdbFOyb0IviLC4JNFxmI7VhYypu
ObQj5TypzQw81t8IuypCfvGuwKIhxNzJCaIVo0HmdQn4IJ7R7reNwb4Bzul7g6n7z+FztO5Q8P+M
gvbMqcfW3scPn6wNkONClWt9OYZ3yOAPej+qNv8qnZTjxMcLFGJz7f7yFs5eYgLgJ+XM5GuaiXeB
W7WuIlDat2UYUILVpwllziy8XLOWlWb6LyJQXIu+AXwafnqWO1dBYSxaeqEkAPKzotDmuOlvXe1+
2izMg4UziHikqtLV0m1hY0/oa1+kgkP5rnZyO6/mW1HhA+jp7xT6gTc4jquiD5xjFNmL7PYBYuWm
18YWfbsamy2GoAh+zWfkY+Jkme5foD/g/NnZLIMQMruVqxlc+R9w7zTUXNaOjzwKqFnAqZbvr88y
Ds7nK0PnmPy4B7IFbZD084XoflWRF0AjVg5l5Fwdn4ez1GVP2zu3Z4ZFfib0brH0gOoIjDslw10y
iEsdBgcV3yPkKTvJtaXbTBO56tSmos8vMFiw6pFNqkMvxboJZfqbYnvQ4QlJ1v7Lx/jrS7CWW/rj
vPU540mF3X3y3XvH2uEG/LV5oYcIJCcc94ykQ+GLzi4sR2+N2Wn7gT6oQSRBUrzIfxlQ6rEc1ujH
4ZoerUvwG/A+TfBo0nzvqLmp+jiG9S6/eYXJAIMfcevGX7jIDB5tGVMkHOO8XzIZQfki7bytER0i
b2IFW20yDzROI236msL7lqV3hkzgAmdQBe8GAidhnIktayFbEuWBrai4K1nDANlOjUDAZO48TYBs
i3roYOf1g+Eg2ZZf0l9XfftbxN1WGHbrCXXeSSXCd+nTusDaMmH/Un69liIQULGmPkLpaHJO0yr7
4jU9OwsRTQWUS26CjtiIkXNNf05qmoW02BwnO/r6tZrBCW1+clVUcoJMSorzUKi0kzjD5Dvh5XKZ
w/Gs8GhQUTsLh4bavoH/HBrdc8AwphOpSSv2/+8NEY76t9VJRQw7EYXeFGg66qgAadFcEpZ24oaR
i+/xUN7oSUCUnri/s4GiQZzDiGqhAB/wNmfPEfsmqpZC3aEw7+lO2Hb6NlD3vkvHLgqwR/54AvjF
tUeVhJ8SunRpEVJ3lpU2c9pdFbr0dt0pCR9upFMfS6ieqyQizmAKQsXYk33b5mPoNrCLghU5LPHy
8OHssv0TJSIFZPtmyCAJ2oM3T1o9q3yet/nfLgSXRBm5C8/b54u+9w5X4oxJnzz0J9O+0fzziSSe
o4uCWc8h0xZ4jbN8/jDiJl9Mg2GRFjQvxVSThRuM1nsaUCTAHE7JxE5uvPZkcvADte8Yc9EGawcY
JSWZUOYauECkIjKIYoNdrQHf5V+jxvW7Q3xT7gwxPXrFn8IsnX+mQLKz2+Wpl95Kd3KMbshJwXxa
kA8WU7A0TtOly/+tCOs4QOWjxms5wxkk5dS8FMNGpdQhbNFdMJhHoBlnd53XgmTdl3ysXo5+nULb
OfjGlei0sRUUbLZpP77AvQ3HRu1EoH3Gbcg2ew0kJpJr8ut06e+UBIeqVx6korkZTjE8Q6OkngwM
WEJxm1OwEuQXG8EAnfUwfnGd3oIM8EwUzNhx+LUV0hKxXyGMXfLEFiZIPd8ZDL//AZwSBodBgQya
is9xMnG/WBzI9Rwra1u9uB5pcYHucZzgiEySNXnPbLyfPgPoJfJ2um2ACyxguNrvC8zMkAFvq50x
qoYnrbWTCmfbRvErjTwMfvCHWOfPiX492/X815hixpbY1R8PERZiAK52W49IV0YMQvg0k4zDcuqZ
g//vKUpbaSITY5N0GmoRO+lxHtO4wgmzEUI/CKMPUEnc6a4IJbXjNbIiUrDmGkWCmSABWQ8G3MvI
blOPM1ySKzsq8wiba+Vt+sIKGPhJHY+0dmC9rd6M72IwPj/stc/PaM31zUKf4EWL4WsCGL+DDe0r
QXhuRGD9ttZNBEEEu8mXGwM8nli5b3yHzAW3KJDpNjY+6r8Y5ycBGJcblKl4qbyHfPvyb63JjnXT
gnKxASpV00uTNgGD4JiywF4ct1fsSA+1wB3PRh6yP7hchU3wrPXZfCx9V9GslRLQXWIUmYK3SA3T
UPwd2zlUxnAJ+5xZEWuBo5zo+mCmnGN2OL/D8kYa+o9Uzu7kFWE6dermIxfRBeLTVaGKvu77Safl
UQnlFIs5gJua0vf0WzTRmjRNG1EOqrJgV1TXDkFmf2ZhnBdmQ4fmK52kpA1RZp/PLAW+Z480EOAJ
vL/cX6WUI0Lei/hks/P9ylo4L5OBF0E5WMJFgb7RAMMH4Q75akaj8q2UIhpAP2VHP4PzjNb+X3Ex
oYGkIRA7aIZkVk1uS6vejM/k5PuOZ4OPqRMVoeRca/T+l5IKNGtz+CBuKpLsRh9Tpzb4O1lpq/yY
duPz79MY7/vTFaIv3b/dzmyYbXowj0dcNH/nefBdp+tyeMo7XhgQnnefCrNzjokd42UUC1/vsdaF
qiFwOv11HGf1uWE/YAXVTzfdgIfZQ8DRVhrHPjr/aQqjIBA9svk7jpTwHCGTvXyjOtjleiXublN5
arOWS/rIo5C2QnPWNpL51bQ2wiasb8iRuzf5/gssXTYqwzgt0+qmyJu1WjyUGAWsu3U5FQKUMNHm
lt/GE5KOoE4ZOsuR+3elVk2xd3ZxPbxZqxNtynmOG3RyMO4UAN8mpm8xhlwdjYg91y21g2CjLh69
AcOKLwrNu4LaKqxov4+luZM6oE1BMWKybFczq6HyrGzkGcoS7X1rWN2Nxb5eiw3WdIX6hy6DokJs
qBM7WAUtlg/LEY1KGUJfE2qHC0uhOBWwtb4HP8G9UuSPkHlEBUM+0L4JCb+tI0P82Q5Ml1/qYvsF
GZHR1sAzPRc7S7oct7FBvWdwiEsIK7p3C07OdGEYAZSOzJLPhZmajp5jhXumGakvggmY1iS9MYbM
OP608Xfewu347tvjOVh5n4BYViX4/0euSOowSc18h51Klwuqk90wm1FzTEjgWQeq3VmO0lpG7jBF
pPwRgBVE691e5d8jwPdaeMqx6yBkTkibxl8bE2al0EAmDjVSUD5qXcamTwPl5Gtc3zy1ILJ0MsLf
zxI6Rew9PNj9I80kOHmULitpa6d3RPtaYLA5A9Ri2jeoXH1uSxmEM0LLnmA61OMkMi+QLmEerIq6
Ey1OP77d7VHLkdU9sHlSjm+HDXW2S1C9802RCan/Z7dPF1uCiACetOhFbAFY0O8e/7eSs0wpeTUr
0AHplWRh/quXgS4xMVgV/JTriJCnMXH2aqQA9PmtsYqIRVtWD0K3bjnYQQtCT1RmEYXG1FzcJbn2
NV0IThB6VDla8zZJ0AwGDYhKLwFGy1c89rVL5D2toZjc0KbpJW7gduU9Gme3fKPa0L4BHY7chhXU
d4dmIS3TwgBCJU/LwaFSfuLsXNEeFsnTdxWlzi3q6s56bo/fML7t7aKWrHxkFP/FZY0HCn+2tqi3
de9lwQuC+EslFyNyAu1vNC9dIpN2e+7k95BWu5em+nuXtdM863HnZcFSkHMJSA4SeAtcPEwb6aaV
qV6JStvL4vF9EDm/crDDTXG5XVuzE78HobyObH9c14B5Bi7MgJNS4wlvZguQjT7CCSeEQdGgmbtB
PDy+MhLfTTwhVDl3YpRcPinH8pmcMq70B4mSVbFKJYeIKJ4n8XsdJbBhLVzNbKF/jefrb895Tv8m
rDYgzKPAk2O+BBQf2T+i30Z2FPF6ffEV8gTgBCyEX8q7Ecp2VCtsUNQNdgedh5nJt9I7AbDavmuL
29ZVVqnSo5aMZZGSf+KhczD4NqRjbfdODH3D74goWyhTr+7el439MBTEDrdu1M6rG0Sz3HorVnyD
lv9QFrSpytaondRhjMxKImf5thxQpB+3jF+AWtOeBMkwC/HQUsFp60K6LiH9PhlJxOdpmROedMyv
rc8aG2Sbc3GXxPllAdtobCIrqQaAk438w2Ey+2zLTePBdzyuZjD+LCyIWTa6iH8UH+tgg+cAXmLO
q55wx1cIq7fSU2ZLfYU5nkUJM+Euapvgyy9x+LmjTsy/0rb68W3DDRZm3zAU7d4uc7rgSrhK7Vgt
8V23kSjvskmdO6sVEz/9F/VMvOXwfPpLqG/bPq+gKfiLK1yTJqviyomv7ZPvDTsEXjckve552nXN
L/VgbGiRFWZbAws9TA1eqObNQ28QXr5/0eWa9X7Z+hmURJQAViG5+XqNYrAcs8HCbFpJ1Y1fF0ZW
Tcys0xKIHXlMm9OiEmmAozpTvxJpO/6iET/FEgvjaZmDItlys19wLXP9GJFH9whizaujlmNzOwWA
Eqn0jGsZLYLmTnPke9itdx/Bqjx3A3VbKnKhF4ReuHA5kDKsi3l0Ufi+gswgHujDrneB8ShUxtYM
Rvj8jtyVVARBXqOp+jwiq2BWZEcLq6bj136qyCf+YKIsEU33U9qSTFH200g/VodBHZ+n7ypl17AH
4ALRsGLIvMdSEhkNUxr0AulhqEz8b4fdhTYhjMTKANpxJZZ5HOzASC612J/JBwBOGZ+koLu3iP6Z
Hm+vcuVQyeb2poXpNZeaz9DytT1CIZoIsZ5QYVrIdp9Bq0qjuhzF/H9UNHYefA9Tkfi5ntCOqZSO
v8OPLKcWsWWk8Wam2k0kp8clTMHVRp07zd9+tVjPQbbisa2/L7mpklEKpmxIE4EsGfo79mAqaozY
KLdB15IP6t9HMEUSjvr7LSgE+7n7a4BH4mquh7a5SYYjJP6WmGID8HSpVZX9648spin8e9uJZpYd
i6L8s2dIC1DzmO+EcS98pKg3T5wii5/LfLPlczqJMwN5VH1FgTWu6TIpaxw/Z8u+vvLE3rkOr/YY
dO1zZlXdWVh2bklc8ob+yaWL06aaixpZN0J0lIbsOls7puIJEnrN/lMutNFBblIU4AIg+iX3ntGy
PMw1EH+ym5ezuli67MBCDp5rJnC/9ReUix8XnU8ZQA+wkUHN5c4vLm2MgVg5kXhswMWrdHy11ilz
CM0pIbnPKm3+DXRemTsQZxFC+4/RpIvA0vORTG06AH7ondpXM6OipNIRHJJ0102VjBRoaapjpmbQ
0ru6DiPLo4tTfCw4IN/NqyS/jvyOXPym5lt55OaJJ7OUFy+P4SUCs9s92K0+Io27x7qKPr2GoK+m
qMBzAIxuETeEfNspBXjBI2r5lZrccYCk60ZPGlKEayqXk/5bvcHUaHfK142HWEtiUvrmWkGlU5Zd
PVcb2e5W9VTHS6NMlf39y/L/uxntEqY44eEM556MnptTk8TuS/hL/DBTPun/uUrQ2KRrS0NbWBlS
jVVU4s7+MbjSO6FTSUTHtykdJ0npOo7CuJI5zjG4R9aFyoxluM7VwoNJIsiWrtCPc1R1e0lijllw
xIuI7nmfTw6F3gdbE4NpH0s+JBC5aCzn85irg+eI+o20EIIsoJ6MTWPS7JYcqFYv+OeNY645rL90
5IJxtQ/DQRgr8+4zdO9NTMQXs3CxqRbyVQ0XYmzm3TO4O/fDiNk7I9pCBrta6/DH4KTjsNPI9oQ2
WQoue8ZlaDnjg1enGZZGX3ke75ThnnuU7+dFQG+JcKl4dgIXvBX5i+lIeY6p64+AlPOT3V0Wpgnz
zFWNqg4diu0SVYYWdOqspy6QYtD0uczBT/lxUZqlSc0QOe04eM6J0ccC4PSUtwwBZlfHO5lCpv/Y
tw3nfK2d2tNKbnxaof9yWnK4OyxppTqthOAV79EQPnIrR24+C6zEYhUrIsy73ux8oQ9tmQ5IpTzb
HOFQ9WzVn03jhKCDsSgHU21LeicukipchsGB8m5uGtAD6HlDzZqeQXeFT2veJDRB2P7jNjkJFZFq
nzTganFrzabXbHInxlw9NNsJ93+OhdYPiVsuWR19Zno+k3+O0XURBZXnH3FdROs3UaWhXoJeOL3Y
fuLtSYtTL1hO00Mz8peeM73k+vnyhvwcnd1CB0Kh46Q0U9/VD/diGPgwpEjDKe8UH8taFMYhVjZ1
akq6oDdUCAnUJvE1NRccDWnYfxwNSztJACOYW8hwUZZYJrIKD/FD8ANHU6PyP6GwVSHFlAjaUygF
hW9HunPPzkIyIfkBursQBNbUvO1cJHZ4+nH/75GPpE+9P/SA6kRColUBnmeY0EwbgLisIpoiEV5k
/4UVcCQPdKn9ZtguP6TnOPJ80VL7hg6dTJXmwznv9UIotKzNDyuNoAZUQU7IvA39qszaWICfa9Vz
nVX83ambhGsxaI6ubtc81Fiqn/m5xKQgU9hgoiXfaB1U0JX/Xiq90MYMPlrZ6h2x11ZMgqBPHuYS
RQBQENIdgd+UzTJFlVcoSuadYBcoRDVQnBwfrWb0yclf8RaGE7HGWG6I7IN001ZZO8aVOVCA93ds
IMYKKHFubgFCeoUdEJKYtKrw9BTTlQ78vyXVocpRgFE4hIeR1/NLg1YFA9VZ17I4mvYsjq8hTrB+
iJnjpKMVIchDydNDKnASEfg8uAxPaocz1YRrr37Si9v+VtdPofsfNpdwxqKTxYgcJl9TtJATjaEv
aoTtBbhgBEDZFugH0A/mVRcvYYfTdC5IWNdbKAj+EnnOTuYNXQUVbD87kYdjKL40/tg8tYHkqPjZ
Y9Y7mzFknals9r5XUnVjQ8ytkM16By1sxAkTQLD04rv8BjBsoSwn2NNQM5pOu7QGMeUR6x+BN/kV
gUn+sHWdSzMcldb0IClnC5TjLwrlPCsLfLHCqeOxLosB3wEctxK3R7ncplHH44S3XMBnYt+eCZds
tpjcWVvYP5H+1CM2U6+w5i1sxhQC6MsP5VUKJ/iPFYQHOo4Rih2c/LdgsIM06g4cdgoa7N/38rT7
eCj/8p1Ebrrn7JWF2k8B/IMBoRhtfErU5RFB54TY7/Q4x38iC616CmEiqUoNENuvN/o05043GOtE
WJmm2xoySrdh9KnFggz8pU6I7m4BdkFp0u//1+nN1LA59u4iS9nJLEdQ2p7doB5RwLge4yx9eA8C
mjXMpJF/pidzLc78I42XxjJuGgrIQKncqGRkG21dzlOleKwDHS0i5o+07qbI/H41GwRudH+GmTQ6
2Nhxbnj2apmylD1Tb4E3xjCYSbSU7vY/77BYXDjQK06f2C+P9qgmO39893eUh59x55uJS1NwdUiy
pC7A8U+RpBz/xeCky3YitVMGqUXtPd4Jry1iSo+w7Nn93gtqRa8D5I0DeOCPshZE8vrcq18cP3Mw
ocOWhcfg73H8bcFR8NnR2/ochB8krmLRvXRo3jbsI4XR0B9ac6GWPv+rznYw3Rp5D/r86PlnZeFA
Pxck2Lnk0jOGyPz4zk4AoS4kthNgKjkSahkWztfX2oIdQ2H2U/1r/hi5gRry+5S+M+0yRFR7fupi
HE8UHs6rlmbSe2gC90WRmCNqQ1V579V1GTazDwF9amaBBhPfn/4LbM+mLYeTtgaK2MsRH9oSlRk0
+95HEPt+ZNbSbmvSGxjSIOJKLlCDuiYCoCY16HkZuLvW6XBhSGAq5e7M7SNU14y67/WdDeC5lYjm
dUn7LfZiZnb/Ha1wRFDuKNrJqVj3yY8ZC7zxwD8TU969JouXLbk3m0gTAFxWcGbmP+I4DxoZHq13
apGmOag+caF+oXOj4E0XmpYW6JhblR7d88EQcjv0YSQWpYXsHQ4agp/1IjGqumiDecjiNaptXetH
jN9Yu1W+WY0TbItCP68uazSQolZ6YyIX2ZTANk7JhLPTgdONC9XEWYrw4tuI4EMbBagHA8R6d6Tc
cpGbumLIvxkd+krZi04rtHVMPkNULkFhzH4UyI6e/g0gCfFnOosNHiJkqcbCf2zHi2LLeEPHWcoQ
kGVok2kWgD/AdXN8rBAyHwnaro3aBPF2Ly7+/ASdatcvBqrXH6LMD7+IfpB0cVl71BNqt9r/d5wC
F3dB5DLOZPV+PPv8BelWWtR0lRbV5XiAzxCHUMxk2/aj0Jmvp/lHm0YCkO7ohILBosSRMuR//PUb
GtBr5tZAPgfAD017/kkHi/KGgPGeOObQCOKd1sEcDaq2+I00iY6y+urRB5OWbLl7X2ufm33elOHS
BCU7WfE8wM+w22NrbxHxvy4ShLsDBnDe/6SBZRt8IsqVdpSUhifrwLzvV0tFrVezgo2IR3RjEEfm
ksuIIDsCGp73NURGVvJ+PdcnlidUsIjFRFVnuSZEUlGj+FqA8z5Lcsale23jlHvAlthFrUFQqoGI
xK5DmFax1RTxoOPqTKb/6kn6t8xwXVAflRZ4J0/fAynXGRe/sqjY7BFHw+9xYhXdGX15KaIt9CWJ
x0k/82zel4tHmpOSPL5+w4Ode4ZFkjcx1AlFLhB+X8LhLhkux4/G6K3o+daXt529DLw7y3Xl3679
taiT8YvLpI/KYem6cJO1uCTJgzSs/Csaz/XrPO8bJw7xUcobnaiJtuAyKc5BUhf9Xhs7xIVOvWX7
JpCXV6gppV8ixvtJ57hjTsT5tYDMrvUpjsLQ/0TUo8U1cIfqSbLkNRR0Ipnx7ALy+CWP7HNYfZWK
r2pUTevJ9WBHvAoE+9pCSNmxR2gitN0O7OdvgXy6Ktq/6e6zqPVxcvAofRC6cPxlaZSj9sdpXNcF
E2Cttu8osRapCAv/tUl98LiLc5xdyakSUM4sopMoisFb1Hm3NaQNJ+UCFhjFP77hUZDErCnIXIm3
X1xmuuy3abY9fkvj8Rm4bAJ+n8KdmzcXc5z4L3PB9gbEMaJGdq3QTiN2tb1J7IGI2rIA39USSeUC
Qi0ESdBqyosAEwFsmb3/cbUuWOFcD2mWrEvAn06Fs30OsfIq650B3tkW24PVVvus7jhZH0DvMla0
toAPGTnwR8/mNg0h9unJZJjD5mx2Cz/4Sy7FkkEZDoEG/q+sFmIDAVBKUlo9/I5qTqjBncc08uhR
8yeCPpxjBJ1oVcdEEqYBGeVzQHIByRQvQxqBc10vBPXYe5KiPrfAzD3/UqsS1bMko8JHAlCMHtkj
DOZd8ngBPXVSk3XwRweQHRIP98ttCX8qzUATILwzdr8cFjmi8HCmt6LKtir8kZ/pX7WvDEO3Pn5y
vYDHF/QFJXNVaznPDnqWN3AA559trr69c7IluTaNT7mPIKGFsCVRbzhhL5I7TDkdwNmxfv3461tO
tliQ+y8DjssRN6W+GMz9ECSUmG8qyGRrOwYP46RC9KeOH9UagmJXoA8tGPpfVY5zJnJNur+HXTr5
PhhFRyq+aJAEqEKdZmqyeaIJ5T4eDVCJyAOyvwPqbVZCo7fuTYV2H1/IqVoqNA9EggORJEOmEW3R
7/RGWUVNoZYSfTUBHFH9VCBkhBsam1dd0CbAJ/jXqAdq3kQBkbfm/HhrPyZ+zMnlCs5e+ATeLf+O
zvYjmpwgKwaami5SSkaxRC7XZNwI1tJLetCb8mYZI0vYn8SGIb5nNbSvVyRHqSP2NJSxyxYra/fu
IrvPsQ7g5y0E3l86vdNko8VEWgRVATxBN3JXpdbAdIor3QoDDPgaEBJ+e7glu6H6l+yVfRb7xnAi
FD9C8aURZH2HyqODNLRbp2WutMs7v9NueGu0Y1Oz2A8uj//kUz8pb+wKPz6+edvwY7vkkebDNG9x
F04OznDZ5I2LXPXlwUkmPFl1L4eXT9NYj34mjKKweZ8oChNwnGnUxc1fqj2pjDoYlxZ2MH/1aO/s
vnNq7P2zZqPbLt/1G/B8Vw9kR5CZJol3rk3xUZrRY7dDof/tLWzLKQgh+O+SgV1ja+P53nN3qffy
x7cy/B03t0QlzTFgVBj1MHrIvmx5RA8FMLDPd3e6Lrzylo09cdFMA1ElnlGX/h0q+2ACoMYDDZTf
0Xbe8JZmNzJPuUdKMjKkiYmdddsm8+tRJMUG6khTF5FXtuLQsANCVFswFOdlbqll7A2Uw5uzFivO
Qjhv+QsggIIfbtSIxmNXzY8BSGaJqhxmn5nV7w21G56m46Il5LUCcuusEzZ0m5XRkWipLj2AkfXt
84+AoI4SbkGPLmjKmk+KIjCik2uiYPjNi+MKb6rIpvVoh0POJKSAN/2O7OSTLViBHCeAKOZg57aL
nWh3eWoWjxYOE/JKF89Vokd2VvB6qnwNX1J5lfxGz7+C9BpBZLaEmMuLTDEu+cudNy/bijK+XuLE
RT2fSuuKsOmr4RzedDY9OEQcXbw4gIrtKavO2jAHiXiwJ5fUHikZzOI1upcJL3hpOR5Qdlqr+f4c
uQH2hjFyZ7DZdE42PgwobA+rDJsrUG9CxOdZiVC/ncZH97CR+OqYCovbn++LfMEgYUyl7hl6vHw1
l7D0Dni/8v2RBeYN47dwjn1TPKYHAZDoEr5gNGnf/zgCD08G20nSoCqxHCsDp74rGCA9FoFRk0H/
zePgp6pVANOGj+H1t0g1bYIIYwVU5ZJUCqsgXM7JlssmLU5lVU1SalXiowf9Ro7y4xU9ibGsf1XD
iE3oPgAix+nxUPgwv138DdFe0oCWWEFtGOXRp/fLDa/79p7Zf6EItpKPldfWYBj6VYLrZCUhm55K
HiOAdjha/YYpWxGSj8r13RJ7yaUk+Hoarw/9XtYOhWaEwQZx1JvCBXsDCGDFDHrcGRX2GIMjQg5W
b+pk68g4qhgddOsW4G9PYr2f8Qr89Dj5JNNCIgkicHZ/HD33Ml2jtdsFpB/gXWZ6fhRbA8csCOJY
plqWChE5WxVDi3VplZlPbkiEq8sTgB15l8r/th3JYNv6S/uhpN1+vYKLb827pRwO1meZf6h/MAuL
qQPkTdSeMQ9mpBbeflRylYy9pRO8qRSgmwllVG3iv+WI9RI7QVvzy1dDShmR5UxmeR3BV50m6e6h
K0yYYxmN9QqrJM0i/nUhsSJwhFX0UP3jbYvcOE6Wap9QUsuB4j+CMFn9/rD4Jgglwwj+N1wbAECi
KOLMzrakKgY6u1FJ/lgt9xQZLXLcyuJbi3bGmkjPP0CcUTZkxCqJaZIe1g0CwGqh7jt0LFh8qb7m
juthlQEIo4hzte8HCadjUiPDGVDQVryxK08CmWxvi1VUI24eLkDsKmbPYHiLz+TEfOfIPyw9x1dw
aEtbx7ENOVvOJ6WZtQ79ayf9FOvXY8dd6xd1KjpvXqVcJ+uvJijknMSB4lYq+wv5f1xi4UM3tZ3S
IzTKvpNBZGf04qa1ZsgA/eGeitALRHn78h8f4/QeGVTOttsTgUCD7AvXAsICg3Eljuf0ed+Zvkxl
nlugNkMyuJ6JCjkCt8WcMEAtDw3bNKnS9rt/4Nwqkj9xWKQygwHaPC11t9f5y4JAYGGhULAP7nn/
zhFnwGBAz8lBaOkQcIWpmJ91XOqTV2Di7C3nxawF9nO6Q8e85FZXPHdoOA6/yEFinKTM+2UR9WD0
qyeixR3ut9xJLtoQhqcbUhWB7++P3qNYDAxpuLc307p3oLAOYmodnDRpVgrwJwppLui7tB+wFeAm
dY4kzlAl06DSvHHyB/VnPBQhNmH4T8vP+efJfHFrYgFvK1n0wGamiZJ8m7F43/c6P32w1Ey2H1zl
ayncDBHiVNksMGmvtAbiGoo0AyZxi9akhFjduG0FHWMQgrh78GghyUiPBhuO3b4Qkub0gsOxIADd
t+wbI4bhf2c7BLV80+WxaSiaFWxXo3P+nUzNL2eJBFGWpDhEfrEYOlTx98EtlYDXpzjUSzvyhLSn
gqcqXMVgO+O1Q3FBba7BvWzShK4BkovDeur2673IvIljLWe0wWmSh0NgQarOwjm+c9NKCYhWFzQU
R5GnV4G2/3BKauZ+M1t9pgP9qJ/EjBCYvY14+ZgbwGsODgOkvVoxJ/JYEWwNbTZ2h/SPlLYCQh0C
K/gYANeRW2/gFBNKhppZOU7Wja8JE9+L7fLXsxTZ4mjl0gMB3RgUrF5f2ov97WFAdlpQ0jwfWNDc
XdkEkCq+8L7VJ26S7TC/MGw68fZ8ToTPmgt+NnmK07URw65o3oRuxnCU6xy4zjmwqLaXnrOkihAl
B+zzGFERBksAif8bQkSscSUBxET0ZhUfb1r03t9xRx7OiND8APcb74QWfRzfig1FP//ptq7sPkxr
v5GTliFh/ppwFgkk9N0/CdnvqRcrVZctP6lGxDFpjFAOH2z+MJbZC2pLJgKy/ZzZNXXkn1ynReVO
kIJ443AiY1bH3NDn+ffDvs2etEZRKYOvOiu0LmsskGxSojXg2KLMryx8ZNL5oAYZEVvWNyZzcphE
Eq9y5IzaujZqWMfvv6rIqtMZofwiOtvy7DA2y4XfwWpbMtHpXYrAufFZXqlTz0hVqwJfiLWz7ObY
KwSJa7oSRiKHrhd8lo2J9pWp2rQWajQjDlvJzW09b8yQ9d8F+zxTkgBc7IWD0FQELTH/yCkInlQX
2+kZySmGdgS3UsUjtYtH3Zy/c2Lvhok7g6L/nzaex55ppBiimkzBuNRYjKD6hko+21gl1iKpoKKs
gaywhiiYg/wKBxuEgHeC+1Bj2pBqMNpbx3IBAeHfXeoO9JgSEDxvY7kYfw7jxFnAGwAX40dOdiTQ
FCQgowreYdrVLF0c5XO4xDh7157tCBuFkeD1vQPglPlKLTYLr/tE4jO70VtoGNaTmPEt5U61YiZ1
vwlnzgVDANfmeDCN5Oa+iz31KW5iD+QXd88gELRuygi7VTpWjiObwVMf1YP2bAERjAUW7KIKtF+C
Y/AlQvQaUv5w3uP3x8LhMVHAacHIDNUZMKviX5as5A2P695mfn8F69xA1trA4TGwfS71RKTUdp60
U7g+MRlmpxeDdKPCpVOAibjcaFE82Iccfqfv2skfU0D9rq61gpk/GDyqohZVfHyfdHbzLqljBsEN
rxub1JJBPbZ6S8Hy5NFbci79n03g3RhO5YHQhbMu8+HA+IftIGYX2FU/Lgdu0hOZHTEh6v/QOXgY
kTlR6WXD5cW3pAECDEzhPmGDYRRjedB5DF+WMgarx4KP2E2G4yaxwloTB5E7rSC7bygH6+nEApI9
ZvVMeQ6jqTvfd7jQ93odTcKytkDxUBTd0zLZWN4eg9YlCDPvZwVc5MDqTPMwepWDyxm2Phbb+9hn
GEV5iMevpnBLX9QQY8p35LsYT8bVLeagcPyn+k7m8CU8DPJJn9uw9kgQFDGCUFR1bu9W8FcFRZk6
xHpi3+LmgbFVO4NfeY2AyI+sZ4Tn7IPjOyObRB8jXhXrX5AmBofxAe7GNofbUkCKrj2MBYe+nqRp
+0xcLXxIKSfTC/h3ZYp3VhetB/bokXKroLy3m/sXVvZMgSkoo+VPZIMQJN/5EQShD9aA9kjIhzKt
KcmWcvHFf8Fh13PlTn6LoovcEzVOXzM6Rnv8pw+HMkfvkFtPx2Iq+XJpR2rfHLIOVW0FGo2n6Wmj
ODM3e8/E3qybJxeS8Fzb42TyaWkhWgw2voTTrRy3g+Oj0/D3ebZ681CVUlvZBnr8ZZKjrbcRQYiK
1eIktqAYis2W7DoQp0107eYtHzwluQZxOchTbTyGgzDOHZQPNbk8xMoF2dnDYYR7Owuwj+xdsipk
Fdd6y1dAaER75WJpXbV0j5kg2wyBkckkuzhOIgNOFI7sdlaePwxq/4ZJsswuIXcsw910bDCdg5d6
lw4fuiRYnE7usW2c8N3kx0qglkJV8kWPcUKQVArSvR2LFTOWCPKU9OnJzwHEtrdnkZkH9qDKLsu0
c0hwjS8B274Z8LO9zcNN2lBygx/TxD/kCshINZjhPCxvjiNx4IeVyVtSlAs8T81+qAwymLaslcd3
nVGDr9QLS5TdCzWMSeCVGy9BI3/nR6/lyycEUW4/Ao1RSI+IcJTYZEgrCKNzxIJ9y0nLaxbS10II
3jej5q8m6olO8c07+q/qBukjPA5p8gIp1rxV5nAk48unhm5cF3lH2IJCA0oorLJ822kmMWOY25zr
vrdteABUGdk9vZ3zvaE6BY8HyqmJw/97a5VhD8T0Ldepfs/vq3FDrLMbEAvvIj8B6vXq9t0vu4BB
63vdA3DIL2Nx/nLYlW4h1CaBJWXaqV5zNP1BFIXZcQIgYROYyuvTD4QPfh+VTqMKv3LJGXiiKaqn
RgLLQbuFffqNAW+5lIuRHXDcjjTIsIiTdI1a/t7KQLjjrGwak3zD2eoXt4BDE2PfRKZlx6MJ+qGc
WSZAYroWUWgzKrHrkRqHqnhCduRI7lgyIaDNw2Rz+wUpe0WauCxnugsCO+lzBRLUgGOmg9jQXIrB
cevrGkXJZQmb2B/SH+GJMqLxlRCb+T/BKdOcyYW9L9avVV8OCNyNSv4R9ReY+Vks2wBPOQl1yn2I
Ij6ReBVuViHCx73RiIvfR2EbunIKp13IaU1Y31ZvIVEYUhZFRAQer5uQaVtTBRx8qZOMG7YzTa0M
PAO5IT1uKj1YPy9v3EdYJlQwRkQKPgr2ojExQ9TQwUtXpwdBFTnAFh/JNLdTF32gxCnPGeNMRwNv
yCImF9JDk0mKq2rtCFVcUAl1sD9gjkKjggjXUibRNNciF9UdOTHTTEPQM5Rr/1iTBJdtoB9Yn/EN
EfrC7BMT6Gn7qQrQmbWnR2hAWAE+ndnLOrs2xtGTqjOsWUeGPMz8sQjhSgx5pQz5lREvA+9zjscc
5AAchSM0B6LBEJhHx6tMsRezJjF1csqXtPr2PqFx5kIUmQQ7iiJviXSlsh/q95X4E/3wDJjPbozO
s9k2ztaejkLKIvQMQrEwLYkPLLs/jS6F7Di/xIGUtfarWRa08rd1hoM4JAFzKX5VjJIF/SP1ZmuN
Rn5UORNiRFi2lOBhg7Hq5emVZuX67zAllFqhwuikM6utK/PYIRHlELHvdCKt7EITNDeGh+lf3+5l
ztaaZst4NGPzJXLYFv+eAfMCv+XdEMcIwOtjouljkeURK9lgKweKLSmjfjsX23D+JxpWC3kiLhaL
E4595nIZlpD72RSPDjgM4vbxveKWRDQxZZ4Kh/1NuFxmCRT5Eq2XC9AxVzkN5ryHN0ZsLNzVnGMx
EgCYSfmdYZqBpeWETYjRGoRXzg2QgVKY7iZKfa+bJSdEDv3p5nEFLCkjpCg96438W9X9rwKld+YV
HjN1j2vzY3t6rArovsh1dsHh1SXEoHDP0RU2ycukByBz0x2Cn9rDHcQw5jsdyWOgBAJapseph4vh
w+sYIgo34QRKhZqW/UR3OW9n4hx8brPDlpMo4DOkUEbUyL5cwSOm6BBED2D7ogrmReRMhLIJ+j8E
eRtqLURPdJE1jylw3mO/Clxd9yIPJ98eCcRu2GZkerQfMf0qN8e+j3Ri2ceECddjTWYtWBUwysMe
mUPURjeo2tBk4gOmK29fRvM+X6h69rjDaePC46XP+TmEc0DjdD0PZwZQBLTypF+OBNcxRpGxRhkz
ZaBwOF60ouCubptM2Z/ROy4naEhNWBmEfSPk8l0oygAnv1yz9iq4uC6J5vvlIJfFKvXmR/jZdd+9
9fql1vXVKcq/CpPMBDei+wiuZpmshm5ghIvYKta93+mH/yS9MJxBDUhghyGzf0LgwUMuRElv23U1
boMQVNVXmh7C4SoUW2uBWfa2G3FHSvJCyQRvl4sE4waGlC3WPAytV9wCLa4ZnWIeSx04nIoKb+u+
6liP3kQPXhOQ32R1uq/mY4ul/4RFMqTxlL2OincVv5Iwp/lOtvZWRpwVmtANqUX4xvrkDjiNMpnz
XH0gd+0SokDdy/7xp09F9FmntUIIgQd/ZiEfqXOAlVbsiU7m0oGUEpyGIS+v+AprMq9wUX4X4M0a
Z4Woj1JV9B2r/kLX/HXrB9jKT6ZKG/X1Gcwsbc32ynK9ori9cx+YOxUjzF8Qq8g+y/69DNpj0wYW
Cbc/IIJmYJ/xePi1AZzczCcF33U6jBO0sGlj1uhVMJ6r7ekHrqrL8bWzprXeRlcrsTZg+UZv9OkT
IMSnJY93DNrTGXjahgyeqaRNQxJc+3eyqHaiwcFzQxS8vywCkrGbaVazDV+JC/Hhm6nPqKp/2rzf
FtHja68xnB4jsllZnMOB38DuqOSqfwLvbwg+zaw8KheYbdxdLHb4OWEY5v+mH3bgb2l5G3+nQAPP
gUSLbpUzK/vKg6kCuoFXbsQ/eVP/wR63/SrOo99DrtIHsUpvRq+VCpI4Wrtg2z1Wmuf0w7b//NUP
kXdJjnszEc2P8nHP9YoqQAUh5fwfG4Ac9gj84I+yB1L0Sa5Kgo/Pu7nfy1wXSbz0/VHoJ+me6/V6
2l6awLR1fXaNDM/80D/1kBQFBGHaL8MzcP41LFuXEaExQffdDUDP8/myq7Gi9YzKRXL55yHwkFj8
AyrEkANjciKoaiQryNmb1RUULwqyQjP+yT28xyMR28ggahM/y6ELHbNPvTkuP4dRzV54YyJTW8sn
NrRsXMbqNZ4cghY94wfA+p0672mTrsTa/pu/cW8T0C6NVJHHPwWn5BwsVoqg2YGmrK+YSqwNw78e
5NO88Bfix9JAynnWUbX5IzobnNlAFplX5m7SAm8p8oA8anVz4Cz+yxHfHguzEDTtiHuKKrmtN0y4
oUOPpBxQvaA/XT5VgYyczRw+W5PpLRF1qjOUY/jzDU3+/LX3XwJe/oWfYb+/DQ0nfDg5UgZgG1Nk
d0wM2k7rAwPKLtS1YsQAjwM7WVMxgNCidM1z8wl1+llsQLehTxBUZSEu/W8C2xseva/2pvNQQ0U3
O98BsEJx+mJQxx6CevMUx4fe6lrt+DTIok7oIR75t4zSUWEl/JY0rZNuloMVDPQ3lq2C6lg0WRM7
MkSj+lBYRQ3oTIBZ9dxYDhe4/WDKuw6W3j5gduWczDPYomTPh+DjBSrHhe7ImiLW6D2v9eUoTpMC
CaEUhGRzmzRyJfCNdKCUxKEiqs5CuQmgNWh9BLTAl2HWfGTHOZu/+JgAQdUU/jPnMvijXHKoDOWm
WFosCARBW+aRh+sC8Hs6wmjKE3YgqPGo2xZJ8+yyydtHA9V0Vyu62IC+zGRXu053Z3XMMJSjvLYZ
fJBPtb7ybmI5UCDXek0hUOvn9f4wKB42TUJoAS1oTtNHxRW4kSsxRNNX5oxhQyT+ZkayLXCUPQ0V
cXaZcMUudWobv1XyaqIOgyAMzMDyLwiVdpC6vjkQygiE6VaL3EiaQWld/Tg4xJLjPvWK1HSVBFw7
2FIvOjcQnYMu3xpXggmQ9oxzSqONkUsjs0Fnx1nSMo1wsrLEaGFyElc31FmCROdmZAAI6MNbpY2s
vcjHSdcBdJ0AaIrR/tRFuHQQyQYgAEb+AnjlUOfwn7dsx9ejr+bMfkQeQHEIT5VPDl+WY2r8OsIL
/0fa9k5Ooq/zQeV5aFksyJRk+YtAS4iYWuvnEqdui4FJ0mE/yOqb88tU19H1jtrRnniC8c76FNhO
oks4CaVhy+ID1oVAg2pPN6Z+qxBj0X9jp0m8Eimr2RmS9PRKJXu7AgOM7ay15NA9dDuAGqYKPqC4
XDGBXjEkmv00xeK/S46VApmNt9yKkbbdfENWFXhNmHGdrgwFGB6R0kTZ6bKBmoTDZGx9AU0Ez18x
NBiCk7ulT4XsA3dscarEfXILR62vd6qwTlcg3U0fZcGpgFMct3hfWzQ0ZtCpZWGYbwDuSpDS+e+p
l/L3wkbccf9Kga4qPo0ZsV8T+sYcnmxIn/nambFWf6/bmJHwtixM+6usS9ZrFJ3iJ3Ng80HeWeYx
7W0yveOSs4aDJ3XqgtymNEcN89Kqoi57k54VT0P5zKBq6/my++MACQENnUcin2hrxjW6QxtajI0C
ZXUkomvwSU3z5X7glYA4e8CdaYZdY31Tf/HmbTwosIY2mdBbNNeK/sOtf2Pa8Wi5MIA2tua6qghq
3BqtwRe2wDolhpY28zZyTrS84u9QV7PWi8MnTEAmYtTtBl4FRAsp2X7D3fWlXVK+ttk3jjLSj1EM
TpRDaShAZbfyAemUcsoidYe9lCfz4df06lGD/erQ9AHhIlsrbpr1k5HeSD2Ie7AT76bYPTrz/wad
4QFkeSsYZ1DaN7wEOjSksfc5Ha+o7ViroLHjOHAl845VjAYT8fCYjo3SxTha+6m1MjOOwLyYwSDK
dGN9C0/6qz/+aytTq0wqpKLs3NHtpoKJPOv7RIEVK1aopcx7lkDSNnG7egL6yV+vqLkS/XyQTZI0
08DZTGM4E1BRSDnb0pl6lfHF+wYweO0TWX+gVOB3NohQDHbsho9yvvBZDeDraTXUmrP4Weu3nZdY
wkvOrP6yGySRJZdKIr0EXjAboG6bqIEuvuOq2XS7OBaDTM0WD62aGxgCQnjLTLlQXPqY77q2wz0r
fXTsw8MNiKo6Ue8A8hJaAmrUoP2WUtU+WiZA8wwnhkyfr/JCl+AIQdGPpHWqjkDryGC2kb9YcaDd
Hsm0+B7wjTMrt2pfYKiiMJe2Z9TVALhCyib4OfnDMl+AWLqubIpsweyu8Nwzkgah+qxYWPFOIjI0
r+TnlhksF3Exo4wEmkPrQ/w40rodpxuSJA+k3iAmYxOxIO4ICvM9ylUhu9nkVkVK/5L+q74HT2jU
uyYJ4jme/Vf14o4mXbsxMUn9dQzvz07nMlL8tRIvEQmzEEnq2sj5MpWc/SI2igGUZ/TqzpiIUuwj
KW3P3AZJ0Tckx9tekx5mDZzLiPNWNhpDlNukrtA5kmu/58gXqTJlVaJoMIf/YSbKpau7e23i66Yk
D9hqLycar8jLgh81+vKBdKR4BWJjomETY4FOmAfWZ90aZ4PPON0EwDCZmJu/vvq9An+sErePheP9
k43eAswjMA6gIluMTwEY1GllUkj81BND60lMBd1a4uuLTXuhJT4smus9M0eB/jKFQt9OpTB4a5nq
0nxRcHPFU0v69QjvYsGERAJFqjJMEPj5A7GUiC8ShzG1kl1BP4aO5ORLD6/RKjvRMSK4QBpuykgH
PtBzr++nzZLmASd36A0gvnsx/7q8WJIsjb9VFT5VQqeCmuxU4+lw/zK7oJ52Sv2jhNI23zLCO3f1
RrW9ohLN2pEI19XtlUVmaoKDsCM9TYoxMM6dq+0iPdbqCZTJuE1c5HtfRNoY1HWPVmRVEKjVDc2M
yrfqFp45IUuIroY7ydb6jWePRDJCubRkeQMiEJEwyzwSu3hauvqQ0w/+LwD1ii5pdqjBqh/Mwjqn
NXMXXwRmbDD8Pwt1xkWtvAUhPbFcEE8Mhnmpajo+uA6sjNvkxGnM2tgGV0AI4+tEVKwWBkuf2UmX
IHsefPZZ7NXa0czf8EhytHbyvrj0vihlGQf1xKx50r4yShn3C8Ntaz9dpZzHVGWXi1MwEUa+wA5/
3KwYX+48f6LdUlgGaJBDvTU8+QAKpryMI0ygl9ichIKzFpGuv+GM8buhb+Le8hjPy8fL5zPlusgi
nc205kNih3XQ7LhX08NJWSY/62sYfDn4MD16Lsd7kXsimPjUfvZmrmsl6eZALa5dion2oZijI7l9
db/6bePls6/gkUgVrZKdE2n1QoG8nZ+oVoSnswT8KkYrWMiWDTYFQh1zUWJDiUDnjBkpf42MuwpY
UNZo2jZbTzf9ajQqSHbB9DWp16gICMRau5vJME6+aEDwiabHMWoTmECOYTVR/Gnez52XrbGfi5vB
mwER71IJ6gHdPMskIC3cdvthMTv90Fh9FRbAvhM07epUGtmKtRZcTP//xQGIw05czo9DNVLiaXna
kyTGKdQhMqgaReM227fz+JPVv1g/3My9RGTTOArLDESjwKhqmYIXpFPXyJ4E+2N0tPOZhtV9b/M+
/N9O8LjAwDXffH11yQxrn2cg4kk9mFo/M9YRu66xUyY2Ik1JvmS4zI3IXeGY4e++eoQjTjl/itQl
wqmtlWKwOEQXhPMHuef8CPTJ7ub2OE2PKWJsfGgUWBOQ6mDR3Xm9WsHbSOZhaATldONc+MJ+6pbm
6Zw8hTUFPJBCZunh38eKlce+OhbR1BZW1SqKu8ZknLZHiAfb01kjGweDPvnz3vvoNukxGkr3lRIS
U3hjc7qx6rhCfu7SOypmrkGaLKYfe8r5TDBzLR9dl29Z4fMQS6UTeY10Lv9WiQmAg11D0T7y/V+G
qH5y+Wb+p4hRNNqlbrkAZr/vomkDUkSiyy4OqXOc6OQPujEz+s8+R5ZUqKuEdodvey6cfI0nCT1O
fsUCl0/NNSHZlQArrRDsQamu70gRHJWxBLsvcTBm+ewhpnqaSTIk1vlSaXhFiqfPqKW+K6gOFsPi
KzWgZhT9lesOGebFXWTTXRBB4IMNzlnwRX6gStPcoH/NFgi6ND6ohaWCrUrlo7N1VkenkpLkZy//
4gE3t6iYpabajV9pqh2U5VlVDc976mamDyFR2qodRncgJSPsQrCmsii1rWQU0Z6AMXSgMObqlLfK
zDPNOgVgqwQFDqqstJ3G0ZPaM1xHQyUV6BugIr1SunHt4qX0FJ112igWy6yQtWzYqXbAEKCIAvQN
Wn3MJNlvnOnPGOdjvl8VbrXENpfpQFMccfytve/0gplZINRVU30OmyQpDtdBYYlAa6iyGRZZXeR/
i12BLGDjsna+whQdlt/EUwsOtUE46QNUxHtAeVs90dTo9eEfxVQtFTWrv8/BDcoxxVToWPG1a4tR
RiKs2P1xz6tTQt736ZFeVYCcor2O6vjP1boIhXvUY4M+9xHH1J4i2ehu/KktsmjqusSbcbs5PPlo
B2jjfE49j9NS6OZhMS6tA6/jIoPyZkutnAmfoz0Asp6RlBYx1XmpXI+bSmcKawK0HZnDdYh15Vxl
NE2G60xXqSiVdnOahxP/AUdb8onD0lpGLLeau82wKEK22kkQhOzAJ1DSn65ZeXHo3PSEY7ERuCFg
y9IHeX7dULKo3d64Y9BPu7vE65xriAQqk81FqUe1JjzDGJtx9PSqfibhgG0feadxmgHA8VKpHlXi
Sa6sTQ1SnYbsETKOarbIwBk+TiPQmY3jTZXOB/UUYLM4phe+lfb3NDRMKeMpt8t8Mib1B7JmXggJ
gi4D2J6QD7qoe4O8Xl3gmEHpor3fFGqekLBh3O/S/I24diF/LeHQq4uhMrLiMps7DGA26DNQw2ce
d9tiVCErhb4HShDDbGgL+IS0YexG+/fpFIidIHr46QV9pMspiPcyeK2EJtk0Ea5HgpMOJOIfvY8x
D1NHsOGhFx9BaBCqcqTr/nY9TMAc939eH4mr9sclOpw9v9epSPRk3gfoJaorvbecy4OSt4ekZtZv
Lj0/QqLBlqfS1WspcZomGdmuAMht0dzb1/XolTBGLC0yuPgy7lbugM9pGiS2LjJP8ooigRxN9sVw
sy2bQRmRgd3WqwXmZBsLohfZ/I+55+t0ZLRIwLMRUEVMG4Ncz9NRES+yi+Q3phE2TZVh91xC01E0
bOr/R7In1M+GdQTA2WKP+zziiQA3Wb0w3goaoi+GKQLG/8JsImT/vcBSmAGSM/6JegnhGaqHJvLs
cZEWLghIF/F3qf9ji1L3WZdE66kKMhIVpy1BAVjv+JOK70Tnofjjf0JUnOUkwGy8u96Xj+n2c/8Y
jMUhE9jsVj460GznnxjjBckTqlI2XqwQ+vGuRfkNI2FeVA8tZUPYioJKdS8e/o0FjDwsXR6sD/wM
CWxnWSBmJhQ0eovZFpzPV6HRXyFyC6EEx8SnQN8Du8DU3CkcaAY4FB4dP8tVHnr5Pa/1vpHK/QvB
lowRCg1Wufi6EnkdS/VPAn3NZOX7ZGimh+WZNYRjAhmJ3SyPM5qYbycY/RDr7KVYphDjZL4F9Fqe
PFKYtX6Oaf8O8DufuOFudiHZ+Dc6szGoVzNBQlCL9VHDM4KLdYvoqcCp4KPGjCTuutpbNTyZKDOi
+E2VULVw795K0VOjRRNTBvdSaQg7BfBvXU/OicYN2gKuG8NAJseTl+Y8MtFdp9VNC524rYcy5KbA
pkvcGjVoKrLevEuy0D6eVSUDFCy8DGLkuWDvgi8533FjhT4GAHcd0FWudkwcwJRRUeNu8W6qh1aH
7u/TZvMsPZbwEWVRWUCzWuA1yFDzjvWHXtq+B8QhxubNHISXc9eUMF9gNDoHJ2MTJgv6bNnKhA7F
NfNRKFy1mBnuH2lwmF/1UJSOg6i+sBgIYImIbowdbSKD+NRHnnjEjBjC/NqPEIJSLnCpOXiY5ch5
R6yKZ1sEudvPTrLTkYpXUrL4S1WMH2vru5gyfmn1N2JBOEdQLEJDyUZmBl3UrL/bGqbxgIVEPaGT
TGLnRJ8oCh2QCnVCVN2uv1FCdaCu2dzl0CYBrsg5VOi8uP+/GLeqRNcW2D8FHqLdBDCAE/cmJOmI
B4Aa7grTqSSKwXZb3dR0fCnPsYsvkHccnxjVFDTPwmmYVWT7rcCObwgZE7+IWPCjKjLvMCe7bJ9x
9FnsLQJS/CXs/Yq7vu2gg9nLum+IiYZupktdkZgXwDBKVVRtNkBSo8avDgq+mDXDBJh8I3OpxXT3
mSd/tBX2oLHu7wfnzF4pXMtd4J/5zzMLgY0aGgpRr0nhhm2hPsc9J1b4NQhbfjbD5Vd3rFMDO/DY
brtDWDKtmINk/ixSFQTCoKxFQWazVUDm24/wpTPMgokc2Uyrm4d0wHp71ch3h9HMdWhfu8cLoERo
20BtyKUVCv1wICsTRm+AfB1GOpfFpnFwjKtqI57pMeMKgTyNplp16ne3xDWRZ2igZZd6EXvzNFVh
8x0HseBi3Ua6FK4XcnoXz3fogsLrPYWUrkxuCNOqC3Z8DaDRvmESJqYqa6NoEkWzMV72FpNtsHom
xopqmmYDmZ9yIRo5aLosmXEu2qhlJsyN/VmwQzZ6ShOsnVquoGFd8kT1ePcGqueF/FTkHtX3rBvQ
9SFCYZ5Sru6Qj9NyQyRR/rG1jt+sIDY8JrwA2znfwtmqKoKGqcpQtcpvHbNfSJnW23baxYzAZ/fh
DOn54oOmR3Ynb5OORnSPwtMDJ1g6bx0e2p24mSWQ8lft7EeW9X4G1xvu7/arHMvxxdCQLvD3N+BR
cZWp0fKAxrhFVl/Z+W7uBQosKQ9roLI60o0BGoiwW5AZnTDb0fuq39nt1Bccb5gqYv0WdRwbaiwi
QOzSQaH4pNRIjx1YXPiTNUQY5AWN3ecqEn0tE2zB71r5SFOHoDne5KjVMHWRKsxfs0qyBilB/4e9
yK5+yuj89LWIppIiPm2XafRPqXjJixl+gkSNmpFlw4i0nMesyI5NypHAlPkDTbpA0GbzYnGn9K59
jxRcdza8IXg6hTM2P4BZxE7KeBVinfThoQ7EkwqpJ2uBUCDr801e2gHU7C7rt92ROa74yuxlQcTg
B68XUHV5IdkqH5u3yuhVutG/+z/SlwaT9x5DwbDApwT/1LLk0Xqv+JES8MLgoAhOyZ3jwwxZo5f4
vHAZjt4BYk+G89sTQr1LxGS/CTAQTR3yuJtB07tRgj6hd10wizd9cHes90F2ND7IGJXBHcb7uacM
xQdCUd/aJTJhFPNeQVsYv7vUzmyB+Whrf4IH4CM3Xdn17/wC1+OubPzzHHCgeBH+K+blOGWVTcLf
UeS0XeJ/YN/9+fnjUiddW1wp/utSHF1xzzDsHFsBdfSzGHBgP43pjcGI7wAIYe5daZAJu6uS+EY9
6HCGRhRXayI2njiUZuw0K1nunm3D+BPXclzSod4vBMZodiA96Ohn8/XduIVu+DFnZrZ98OipkKs3
qKPboxXWbOW0/Z54XOfUpvMkEsMo7aCLh5oQpRfCehoVMsWI4zmogw14+9SaidjX0oKpPxAPPUtb
d7KEpY/y0htGoJxT2rU7MkHWrmvQxDJfVNBH92c4A8nz8uAudQstZj2ZuYbosRUrOJ1fkoySHVPz
YfcqUAWEVtxT2c/T7vFP5N274mDUc6xeUNysNwJsYb92cu/lC6g9hEi6IGd/ZWlq0Y+YIgWgeZxL
4OCtdnH9HNTqgEyEDuIQou3GDW0S2yD6QXCQR2PIh2HppUVeNoSbkYxa5rkRddrjham0KidXefD7
dIRg5z1Du9I0Pdu3TUyTZkLOvM8sHRfJSYxFRJiuw/d/bViGgcEHvHMFGsB754fQpCw/IvUldVnJ
CwZF9JqTB5GEgD5TDgOMJxdRxxZvY2Rq+2rTOUitPJNtHGJN7Ql0ulQeOwq9uDodnTRNW5AX71UI
p+kDu0CaVWnXLIY0QkUNRaQ06JaGmvRC0oPaEiSoOb31R7fRklfSD2DT6vsMdf6vPBzdL9psbflf
ezekdFmktRzDuwn1K3i53QsgnyFQwMuRXXDrcBqSh2jxQO05o98qAiMNT5WHxAlPTi/oQ1W9Mry/
j8FnYO/r90xjto16xc71MI+iz2Y469U08Ni8dEUY9wNsGyNmJYbghG+YyKlPQ/H3/VquFD+BDaDY
t+P6OIEkrtLfssZakHY8jkK1U1zc7254JU8ns4CArUvyWZDzF6p3oYQzwCrgGRSe3X5zSbg+wiqa
UWnO+/PhaqhdFDjqu4g3qO3aS9NA9UXQmjx3gOp+usNkDs7q5AZP7URtx+xkB4je+rfaLTZz71Th
ybl3Zmizre1XY8Fmcq+heD5hO2lYFuNUYxEF5WeRxWZJUg1X41J8HJWSffIdBxmCk5yxQzSuCez0
Y+2CUFYVWOnrM1coGCshQ8dKXUuBYmd32N3zGM9XluAQUd4hT3tSxNyBaoxnMIY0pBpSRn4BzIsw
e9AsOT5uQQN63EWA0+RVihTUO6DJtzO8e1aL/Qpolv6Bm1G3CRBE9NuNnsUTbZskux7NW/xeBsHd
7ZiN/lUssfOX/pGNpCznsZtUjK8XD3l0jzffvUoanc18H5vR9rX8jZbUkD0G1ehFWiymf7g1WYT+
PxygjA1asi25v6fq5XF12NtwfrV5YoPirKbKdzahm19/frMeYvzQs8xEypS+1DyM2u5qdXUaFGeA
/j3EBGuZ89GkPrYih0GNGUlLU7rHIX2Qux5Yt0buH3qv7nnHkV3K5A1XlMPYHLzEyly92mfFRIKo
uWjY3bvCeCLLqBSIGMpV+PU41UYjkiJUGteMCKbAS9WK+r5LABa8Qw3+cm368oxMqSWalJAR8EsQ
SIevGjmJEMQ4SpJqynTvlt3Vhewn/NTPpA/wEl20Xa0Pt6mgjKXRBIYg3QnHv8l3kUovRZi73eZ/
7eXn8bo+b8YJu88klNwm8vtJhVt3Abnn/SNgASXmsV9bCGcHKu9khpbEQOFAWLVMOdll1gPQa5H6
0PpPiIv8pi+pKtzTAcrKKsN4wncEyqu3IVBIk+xnTtQSomEC3HZNAybHai6k4qQ5Qadh+TZ5Fb4y
etub3cc1fnbob3eip7Prj5dCdFAoNi+MYnQjKiU1ptIAknbkiVZYbAT9Qxh/oM7aWjj1arkiioJZ
oAPe6zGs6QdtbupoSp8D6YopiO6WojrbNErz3+fERibGJ8lHu9dx5zRfGtKQbtz/IJLwkSIBQHpr
mO+OBWmoi/N/QndxF4SB/ORv6TvEGq8eBwdj/hG3rmHEFKVnfs+WxHl+XD0VRHHDxJ4dqxRcWMRS
/xEi0bDnQxuARaRu/JsdTnm0bLlJLaf8A4NwyhtHMrYF30Z6Ixw32tcFccLLCXI5KKGQXgHjjgO6
sB/6AbI99iHTYK7/jRMPxDyGnYaG1wM8VAWSHNqUCtaJJ3AgPG4Au7md+0TJQYU8oPgGBKgZi8Kx
+OUlTRshMqZsOircaQYv2l5tA0p0aVwvCuRIMb6sDa0RVV5wquX7VQ3hnFo7zWAlBq2mhX16dSuK
4ZQ59LQFlw2NMDs7CK45MRR7iosvIMXptO6p3kbvWxEwJzNIqVe24RDSp6S8QATgmZKJOna29QXK
Hx06/O+7gAsoU4goB6p1hLsYyuoatKOAhfqNqd5C4SCfz7Km6G+hHXSkcPDnp9N0dr8jTz2MNt9t
Yfy6tg6LKzDrxiJuWpzX2Mf6JBAV8ugPVnAWr9XQ1sd3UCzrsYBwnmtgJDDiAyd/2fYsuDk7DVro
YtYv5tX7Sei93+RKawvkWW8v/9U2bKbt3r6ybZkP9IyZj6pYGIfg/5myZZsZwx7A7G9DqxZ9asCS
OZflVqU+J2XmSNJdK67vq91vhALiQw3b5yYCiVy3oTpaeBaiPPC4Q5xVepe6lUbqZ86vlyqYKPpo
dj9L782Fnf7AzCMzNoINiEfzBFNMe8xlKMy0liqK3e3vAlUGeP7XHBn5qG3sgSWuPGZe4cfzX0b6
XWV+8V561UvYh4FzW0Fq0mNFLrCRkBGu0JXiNbhfostz8WOSeGNgqfVZcSVVMtwii5M4oHF13xKb
r9FCkHKkcG673B9MTNE4dC3MBuv7v0iH29UpNLu4yZsvG5EVGAst4YrLkO8vSFiCFJ5zwpaDdxlP
0hDEotCOAtbwWhzjAua5yPeYYz2xIeSgRImvjc7+rIzg24NS+h6VjhFWKi4dIPszHQwg+z//X/J/
IVJs597+a2WzxGDlVLa6P3XmNiWP0qaYeKuD+bmPl7ROL8C4OaBwiHXQoPEP4qz/XK6UUY0ibkrq
/nBtOWk9fvrfB3LeaRObTQOiWHBEtBesuuQm0AAlEghimqqjF5Q/d1NX9uJFAj5yucmxcvmbsiEd
qIuMBpbwnzf+IsYvlJf4je1aThr8Hdj9tGdw/KZ+JWdyammRsAddxl8Xy/X+UHi54spcUyyArWg1
R61PE/piHlp9YPAFrOb7zMRaf/OjTN9VNEtCBivWYeoFnyVlFRKQ7gfJEj0OfgTxRuV8C+Yp4Uk4
rZokcItS0UcPpLDSlnGpuMkdz6g83w1OxPjSLTfnrUATDrm2jFK9Q+Wsb+ka9TzRXKBtbhteHBDb
TwpZqpon5UfaHnjuIg9zhRs1HMmFhq2WBKSHVsu8RgpyiK9HcMnwcRDDnwPCXE/+WMixvPMToMS3
F28Ao24mXf66PeDCEx9RWBtFDDnmmbyjlxOdn2kfa2c2QqzFr0C9JXyM+4ku1geK4fiL2ve02f99
yNCfuOttUK1vCB2HGm46magH07rMcgCt6UW58NbXIKnHvMFvf7yyN9N6LDrWADmlTHKsWnzb0tUY
BCwPY8tXKxqHpGLiQWK3MX5XYQriPJMVIF9v5KGmCry233TLBfaoh5grvzOpC0lvXO/+57l5Qg3o
+bDxiRUHNLC15DGm0oqll2WXbqsEL1uQTke6OhWLYoCGRGRgmEIcudZwLCCmnCPSUz8CRbJUWcwy
flWOJk+mYCuWZhGBoSUce00k9rr/Vsr5/v8S8Qj/2TRIbShxsOuvKgi2M119/0vF8g5R99Py1Zln
py6y1Dlsf7KsYChhrFW6RiszX91OSmsD8dxQ6j8vDhgsvn1v5ZzDo6pO4x5iFRWkZSSZ5IL9xgT8
h81lAhpxWah/TwB6VpmD3bBGAIX8dwITd2Tb+pc644Kc3eSzEjIYf9rhc+U7zvt+OwrXFfPKftT2
AIpFRS8LgDz8LdKLaJ6lVuHB74b9uAaEnBCZASWDToj2o5Hwgrxdc+he1vs2rBMxXzFSB+CNckMY
wG4c8rWd7AXt5ZKQf+6hPFpoQUfePzAIwPxsRBBA4nBG88uJ7GWAOJluY0TOrnsJKBnMxOPpFjcl
uH0jBKLP/Ebl2vNzfICFjRXNAvADGVSj5/z4ayKtTuXAk0JHL0EoWIy90G4ptFRTlhVkFkUmA2ZU
yT2aQ6J8PpyqsgJQv1v6iOYtYBwp5kF50MfMUJ2NoIqWmAaXNz2Kj/Q+7m/I1Es+2RPIiML72JYi
5X+Hcycg3AexMlxRoUiqDEGuiJfUsYfknorDopB0cVo++sr+eYnqnd51XBG5Wnai15zEQzFHDX15
toz5CmAIuT3Duoi9lCqwSz/YYue51DFVtBRzU8KBnT6NDv6CXOkV4H7e5ZdUzV69/NJIsCyCEFAT
4MT8hogJsNL7Im7GvcaszfZ2TOGRTIKUb+s6AOxZ+Zg7fK0Du+2+n/KchfMZokUJ3QVvXm/e6pW+
qVjfYp5zVDcSXIDEykHAGtqAAcUMymFaxWmgv1wzIPQfvx/2ZMpOedjeSQgy3VpJ0GpmpejXX0bc
0UqkHmYDzZFFCW+zsfR6/ukj1r3ylBkjJ/Q3fqZDbGH0KoNiKshPrptc1ac/trIjZRH6mHUYywJS
69G+o+4Ltnc77LBfEhj5Wu6TPsIifgtBD6ILIY8SSlJ/rly8SaqGuMeHOjBh/VnxEMdD6QWb0nFZ
tctvAwqLoikrdlS/cxa8gLr5CWgMD4v1BObqb7OMtBylkViMlGQv7oUUCM9RgKczMEHkIvJYAE67
IgTU8PyjtzYLdLBzg6NUKjgFbYt1gPDJ7dGBtF3YIMf8PpMISF406f8ui4RgzjalleqJj/1gn+YP
h9dmdf66
`protect end_protected

