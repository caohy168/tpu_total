

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NzvuEx0G5HwsRW6LabE9tv6D7miYm2zk5H6PW0m/i/QjtjDng/QoHKP9dRkjbY33CGdh9buWzj/T
iTEwIfiPpg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uegFRRymlgiluqMREKLn3cmKVsrP+ARyKVAzvWBCZjZFdPGfyfY1J+5BT3DHkkLkddk6wXmHAzrX
ex9/7rPxn+a96Sl0KbXb2fdynfQE4js4WZ4s30akpkF8OkkOgqy23iNrGN18OvdCrTBqFOvQDaql
PF+LonzhjBYxOrtUwws=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gjd1vqFRZ8aTV+TyahY2j1KhfJ593tIUNpKdAVhQ+EIPRnR2KOwC5rRL8piYbMs3haRMFDq/M3IT
/aem+fv27HwFPFJmLaqjvtVRcHzMFp+FoyAcJ2mxiZH9qUywwXzjLPC2Ts3AYHsuVmpURpaacNOm
cFmCLiN+R+wVCW+cs7dE/4hICriINqxB5Kl0o4ROo7XXB8/xYi7xz/etzt2PGPKbrFy/qH2lBU2d
WiZg1a7PxxaMbHGX9OoSkm/vIR1ccWUUzgxhyxc2V5sGkjZMGjZa9ul1SfswjtT572WnNbWtQe+S
lN3rKrYdh6Gwx92X062U5Gybd3T/HBAdBci5XA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
geKqy+6ber8+msEscNCFadd6Y4er7BUAQDjrZkOBYXPalMttTjCT0+XMYDc8PJKznvwRMh6ooDsj
LZdawq+bmAdqcoz5v/4rkkmAhy0/ncLLCypSXP5X9tWWlUoEnvVbtlwfC6NwKkePEGsy7Fmll9Ad
2sL7f410b6I9rE2IjhJIwoRdTu4EOu/DBmpRZqmekQ8pCo7+WwNVxtdxvTIXxS6muy7qQay/fcbh
di2a+gCDWGkGZihCVDg6775vyIidmBIUs4RCZKuDaNMpUYm9/mvn4/V9TEHX+dBB/h/2zp+C9tX9
ynvTIfmzZkBKJ6f9vk6mvrM5IXwnG2qcHTKIdw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dsuUaPzLcdY39SvSBqgPXClrpHS+X1tsCzGy0CVXwJqaWmB43BH2+kL42HsyYbHdRL1d1h2W9PvB
NeliTjJoWFWFvteYzOezxoQPAKCK6SgqxafIETsM3orD5vr18SGtTi/27/T4Y70CI97FZK29oxAA
JItt0oJqYNVIthIcBKWVAEvAm5ETp6YZ8bqYkDu7w9Rc5BGjflKjMZdaIFkCkrvcZZ8pEKx7wlFE
NnHlPu3SR6Kg0jKzfjb8z1TU9bx7LxEY3kORUSjwx8tq2Ba59wVbVpMd2sUfVwCKuzW35pdVhJx/
EJXk4dh40/eC/1Hc+4WQopogb3oGihfV+iXAug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L+I9JABBUZjbd/CC5epF3i0eyHgklkuFl+d5sHWFIHZaeNgsI+CYpI7zMU0TujxRxfXut/dDvlCU
znUHjYaZoSIxQOknBNW29IlmLFK3vxW1IzTKUT0DFvuI66bCtIhVRMdhW2j7hIggeulPevB2fnaI
YkWXP3KoSbtPRhHzRDk=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IBPd62E3V1LjxCYxudvor1B0/8+0308rs3QbnuE1+UsNAPZqssy8vAjEL4xFi8qCeZoOXq9+LlbN
yU9VHjZDJBurvxM4T0rHxh0E5u5mGThlHMCOeTi6+syqAtm721hpkbPDe4TDjU/6M4uKwh0fRCm/
1rV3ZeaSGS9/RoSU7wzUf0kFz/BvgZ0L669JkBQVFeiM/p7ngOhhlXZvPksUVkNTFmoa5U/dV7P1
QmboeZWjz0j6lpYt92ON9/ofUBtpJf6+WuHFpNxXsPjScFxhnbYRXM0w7GUtVfZ2VTDP0EbXwOAk
TlVDgbAqmCGp2OZBUn7nvg3nMIcXVY0axMVNOg==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YDu4ql3XCT9RyldgwN4GvJ+W4jcRfHKJgosq8hibl1HWZYq8WL8TKFYqj4JqsEg7atYHTR0Mp3R5
YyCfO/2C9da2AK9U+XFlUv/W/ba2Swm0HZTdSn2DYsfeFh6F7zgHhgjwHpr1DnRqd3bIXcRMVxPm
T7bptSqCjMDJGTaEJhy9JZO1/RuXxA8CbNkrfR9zG2Uysg0p8sg9BRV0Dxc8R5wPj1KHbYs/bCxy
YDjiii9PoM9ERF42RFALedlZy6GwuiTb1zy845keOhwWyzkdC5w2ZuJlgvkTMgB3KU+H+6kvnyxt
B1qfyGwWxzQtacrl1R6XexCXBW+tjYwvdEeDbQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
uLQy/a/E8+6bjaVyXYZ4T7i959sX1qe36vlHV/CtbegJUp0TUPWow4hx145EkZ7IRE8EPeV9oSWQ
GgivJugcsgdwciU2KFOBXfnz9+3vfA8i/+WGSgezcu6yvxusI4NOtWzRNs1LfXdKUCu208JDPGj4
k6tVFvKDzqBd3+fF2oOZEyGrSkqkNxuntOe+aE81G7jNLuAZbVHv4H4r2sCeV3UN0NXSzM3M0mTn
hMzYK/kTUQw0alBtbvCpOd6IPzt6KiPugcDWdwopEajWhHoHpBZjXT05h89hSxKdkTCcSmVE8mDo
ohoaDi+ThQXNnqUYI7f5y4CPtXm1m2S1d8nKZQ6p6SGjQnTP2n2FlmbOO2lsCdKf5QwdQ6Yx5NOu
k4UmOR77S0eqshUDuPELLaxTbX4YjfaalXxgJw2PWqwXbTmYzZ3WUO7rG5DrxqT28yVdx6MNzDI1
tR9eQc8VyR+z1OoFzVcAAz+vlhHAtnTOK26TI5r02qF6IjXAxGUBlEGaF1aE0LhzbcoqgIHhQwsk
tV2O7DKRibyQcCkUK98vvtnv1yRYEk2dpEoov11QMFJ7wkK4KtmHplyHUya/ejn+kQn8MgCJ6D0U
55GEvoQ8e737s6WZMhhbUc/lPd2a3vll2A3MNDG7R2KhKdKckDaoK1yNPt1uHBJ1kcyz9wanoc9G
nLgNZXT2mJGEn8sv8QE4oH0LpLOVKKSRDXIRgYcEbkQkVG9M/gTPtQcukBTLuwN4uuLnL/pj6Vjy
IguS7xGlEWa5uTS75ITIv2oSioCacYQ0a/gOWBFv2XvHt5yQlz4npLQF6ucqC8ZaC96Vqcnny+av
04sQCie2Aqk6Gt382+l1mWysyanNQpSOJYzMRAowP2omJMvS63f9uvdPg1GUvPtVnxjU7xA/DmNx
bPsLfhMnRR+7yofSj7paJtLcTAvW2+bryw31QCZOE4/xsVFOS8E+4HlkZ1PxCeyj8zGfjhHG8yqJ
SZfVR3zVNLdaVRnivavKxz0hk187Ggsgzt+JaqcLzrC7lF/aJf7J6VSCfDJ1Hbu2Y4LW9zk/UYeG
WuK3sMy5llgiuc9CMT3YHFdgbqNofyE4NeJHh7CawGa5A4NGX7z2IMHSWFZaZ8weUA40uJ9DOhn6
kZbFbVwiAOXu7kxUVM0+YrH66e4cvn57yMuBXmJCcB8rBmp2GHleAmORw/pwbAqoCJNW3yq0JC6F
WIMrNRqAhBN03AeLmAYl1U3OKgNajFjM/lkHfLMfeFzmFvHl+2sjhQxySHGjkcKFVfrOLFipjqPd
BGmVbFlB6h4UgkfAL7nbyeRE46OPtnxY/R485iSui4wIEiuy4dGHNzTMbvyiOl2S5YMOcI074Y2u
h1bwA5L7/cchRMXk/T5EnfBNgNBzo1OORiGgZQqWrdc2BLrNMsSzPSkRDBNM6LnyZ28RiT5OmfFb
UUM1YRpgTTp6Qs57E/r9hAKjFSsbP4YTFk+a+X6OLw/orUm09PQNGG4E1CLw6vP1YEgdJfNf1ftR
gDI9zmKJ6G7nddEt+zUrkZYVB7ADiewchtGRGUF5wOEbGrJlWpW6GDTAjWKSa0QqSMrwe/l3tvMA
Px2ZKUqL46yw8a3kvgyuHalazNoOWu6eHfKeUDb2Emb964nEEOYSU329cqGG+NAc1HcmIUAeU8Fg
N10DAZip48BnFKRIYr5Jo5mbCti8UjkrthBlMi303RUPAoRGhXhiQC57esAeEHLBTHIGgLJGuV/+
hW2z9ljtNv5ZwwGWnINtmK/RfLYmvmhRJzGACF7By7s5jRN+fRlQcSA+EDWku5UGzCB8aDTycyPU
LhbteNMqel43KXxCF+GitJhgEJUU0jPxhX+w1ILeYc+vUMaWc9RjUm9f3Tkt1YYgShHuAnO1DJQt
CRNn+bgjcw7QEQ3GT6vq5pLi/naYsXFoKRhpWFizZcPjb2HLX9HGmKP2F4xI/cIvp6yNEQ48GrXY
1IM3vak7lqFryVlKb5q5undcBB19CsVFCBiNV0zpzDuUfjKX4XF32T1KK7tAIFbY9ev71LD/MQ+K
598e+sl+OMQyQhmLkk3vD2Q9x9D+V6y0CJFrt/4kr0iOJgcbchchQ9Rb09z0zCls78B0h7F+B/ZC
+K4F7KcrzTFUNetAablklz2UAH2Anqft/n7+TYwwwsE7G+C/hbreuxKUgaQ3HnXXJG2I65JUzsuP
qQkv9MTw+/SVnyDJcqeDZ9jPwOvk7jvEpBNPjQAF1dCHKcsBhNTfk9NQwv+zQmQM0A4ZNqLCmupn
44fuK479vBILril3tBnQORvn12FtG2XYYlCXeW8Xk8AhMpE8YTBNwLWzbGqqKaCAEvR8umdJwkeR
lZp6VwYkOvBbnQvhFiTaWC1PnK6tgc6Y8DyR6hjyYOc2P1OZ/35gWmIbNAteKZDIO42B77AuOG12
i3X1lAQpqBu57Es3i3pn4M4S7wgJVSLNzWHy/rFX1xhws+WMQKQ0x4DbCeEDJInayrSLBopyf0Fv
Jz6Sj3H+n3mX5HY0z+nuDg6JkMWp1KGiztPDoiFm3h/1OdeC0l0C6THXG7GGXtlGk1+xMyLJsMD6
fp7WWdsrzev9de6t3dbvBNrxB6lA73iXa644t6AJ8f+EOJRQC0AqvJqNmzS4KAIyzV0nzseQhUpz
cdS64vmYYZ2zNAFGd7fmxmvguRaY4re1Ej+WX+p4CkAcXxa6NBjidQuzZy2t6D5+5jo1B5MqXss0
WdGN+Fzd7Bl5xWfadhfrpTm78pZEAeGZMyv4cqV7CpjEdsp9MoTlLxoSjA454QJW0iLgONa/XT+2
e7LhK38OkUK7Fa8BtJoN6neAo2yKf0aKVAVngIkdA/Jnu68qfo4aSmzhMWQg2jnritE5eg1aQF9k
9n5cjiXsGmP3y83GT2l1W5p1T2UvLU5IcbRey76CWTNHwmJZeuam90edvXBfLmoHq9Rxg8FOpCwQ
ApZzFo0pXplvYOzSZugzeRWI99eOTBLllvx/REFrd2qOh23wV2JtR1TrxbZBCYfzz4iQ3WePqykw
pmnsPLJr5mA1RNLkdM4qfpfUVQQkenK8pG3AjjFy/eRXJfmGx3ZNhzNIKaAnNm0y6GXmEG55aVKj
NyXemOqMZN5LYM+fh4+nnDUG/zAIEs2vN6+/AscXCQXLtUiS4W/7hT7GR1n/k/4I1jPuoa66Q0Np
IDCyWxoJN7ySPIn9SFWLTLHC3HAknRUR4AV0/vWnIQlX9NRzDZEgpXJPq4F++wcnawDvr5yzO6Wt
9ZuSq5wMDlE80Ca9CRsAz4td9hiYErl9WgLRPxBqUKgjOQaMtN23nknpPq+6Omr/1+On/VqPAyYr
T5US74Q2l6oDiiScTnPuaUI+rVlfjpwpgOx5YKDceYN90IGg3jMfp58lLyIqkDJuY5wMD3QlEknH
zYTTn9RKuT1LA6Wn5U2+wexaz2yS+hJ+C3fQqofbKwQ9o+tNHf7hOdj0Cl6oTuJx6fwd4hNZBNk6
To5mVRx4eVQmZX3zxFPqTZc9j/fo0nxx+R8B0g/x8RYjL3lJB/7lzzxewJ8/o01IuS2yIJuQqwCn
Dhnie6wUNVFRb8U2xjwxL9hI0s9npEH9BvCAaClKkQhuXnofq7f9UkUim7shQiX/sOEvdInvzFv2
wokfxv6rU2oekw40suoDGqlKT3r3o3NdsqJqDrb8AGUePhp4ESFJsM5v/DVXr27fhBjJ5+SSntSe
lbHe9f9FGLob2K6GJsHeiLyQw6J5jF2OOtV+hrFDJtQ3t4XnJ1iFTajIY7il2/kqKDY2hfu0aMDr
0hcBIz8BX6vmcOWCYbAlHyDU0ZWD2B60pG6WP+fm91C5J1YCZqiJ+q4s6dcCQKPJZJynfOamlTWN
TrIbUzSCAMUe2j+bb6pxVmLMzfcqxyBqjR5e+nZ9FSIwhS7VkgOHR+fyBSh8FRiT5aHhIjVKgySH
mQvvvVDQK4+0dohNqm5Wuz4DSway+A4IIcmJXJcEy8o2a5i6IabN87zcj/oSSplRjK+5v1VQMGZj
c7psIxGvVC/LdfSz3tk+tNEr0XW6b06Z4/yriEbb10kwZJnS7fVYzJv37VBr0be0Jtb0azUeaLKM
wJM8V09MLBX8vfB2GCl6S4AhtPMk4+QCeQzff1j0oI2f0C1T9ynB+O6E16gmGv76LeIEuF9vVLiX
RORL3LJhHgho+S6LQEQ9IwQ0BzRbtEgwOrueyBDVh28TVIECKkBlqmrdnL9I5uTcDhkWp6OI/DoJ
19x4E5ifX9F/Gjjdf5DVQ+tm56HgNSNQT524s7eHJncmt+DW9rJm+4CNWtTmjMHJ9hH9uH+SFn+1
Qxd/1KRLJ/D1v19z5K6h7oHGELVmy+VSNNEfOdp9E+qAKvheBCNQ8oKLlwO+JHO5sYhXDkuZWzK/
OOk7eX10CJgxk3FUHFhlQwhEN0y3cQBAoLp1a0KxSu6vZX/17HwVXZ2eZpNjM188sKGCOTCvvZGm
uXZry63QFnH1jAL3bxk6e6gsIEZ1czhMkoL/jlbKtLM74Bsc06UsZBPIY5GKdAPPesxs92qeFUss
oT4jZO4lwN6/0pJdw6rXq/SG7ToHdVgDLqYcXtP9SuwsrYpinqzaw/fv5Nu6pZZnFXVcYG454XCC
P5dL6d5+6PBVqyp/4L8UDkNoPLY4CrYwEauH4LJhGkLBfBsKN4FozgXygC0oLVq8VGhaT+JKlTPg
la4R5drd5/FVLI7SdtZTVSbYEoWCXelGkaceY+7cxsLuKblcIeMmk9z2NlZo5D2t4tDus87YI0pA
+HTIETFgvx+w646A/v/uPoHiW80SbgvxSn9Qu4J5ZJLnt766BdsCUwth+o3NaF3gp6s6bOR5P98L
iu+HAXlVW7a/BpCkn3y5Cg8xz2T8LK7PoYljSurm8CXQWPjqGzC8EPHIsGNfRcB29XbDKD/QeDm0
zNM9lgx++7FbmW92nWH0BX4RXF6vLhdvm4y4qaP24pXQfWjIIXVNyJhZuCE/7EYIFaEU2VP7dtCr
HNEgaNG0j92X3OVYL2VeEYTVtR5m/C8hGHzZx13c+ubiaL25f/IKYSO2E8yfRSHTtG/ymM515MZP
MoOX1l/wHfIXijd+zZbvtRLUuWoU7JRKNnMemGpqj2D3shEKpkHDO4BQi034RJ3C2Iib1dMyIEG9
biSiDx4BGpmp4wD4kZ/JaFvkD0m0jXdE8E2ZNoxXT7nalJo+4LnZUiz9E1q6yYHXZ7ky8ryQy2p7
qVAzQlFFeG7DPl8uLCiqC8Oy73JWn/WD3enLrJbgL3vE0UCGvkGWYG7IZV5aiOK7jpX4ud/o6ial
57z0jRfa64KvSWDSoZiTet3ZqV+3tyKMzn2SCysjWM+q9KTMJ0UDhz1XEEEjpipVAxVA7k4E/R8h
gO0G//kjJ7aYGa8U7sYPpzmnXJostfvlsfuIYJFeLRsKBpVyOuWP+mq7BWkkN22UEMerzx9GOTH6
SPfQKU7Gby+5HExImtwkL5XQ358j0oqvkqZP24SxA1oVsiaGlmlBg4D7XOCVfELqe8cwZ37l/wCs
9u+tv8I1ThYlapnMnJT0vOP2mJzpgl0Z2G3V1q0reqi48qwt0bkiGYTme2r0yyUZP0cmskcDNlpV
wGuje1lbeVP9apxF/pYTazXsleinOelQNoMfxrZfJMMbCON5zeYfBitLR5P2/go3CPagehTuS1yu
4BGu80KWZgNfd2mVEFDnZ258JTrkRKRIz7rSvBMTOPLHLEECu2kPaP/2rzQgC6YpqZ/3WyTdYHQt
7WxHtVH8YMZLfaf3UdbTI/vBvOezCa0YbPNPBsK+l+wfnMCs3MOFsXUmkQvrGwxDaeZpSPGMZdii
A8T+SZSH5pQhPnuQSPlvAPFKirYc7+HMmTduwu6RdXz/qOW1appl8qI2JvY0t5UxSJlchd1+5+CU
qvW3b9sh8VdGsqf1MRaDCb77oGM7Jo9xRHV7N69vBOyrn+Z0Ay7Fm76LGrs03h8YZBN0ZhglRhdS
IxWl/EPR15pBnIjpEme7dA7/9ihhvg1ugbYmZiADvmtfodga+PN2jww5I40tcBUs7GuAQdUWxPgr
pJ0Z3tDKnRSU94Orv5QYFfzSY/mMxXx3uV22fkW8lNrKPnh3/BzGRhAsHcQXAQ94YrQDdQhyy7xM
d/rSVYiuovPSFwVkVGuJfBi5gVMFW7zDatzsffTH7dgvalhhLHa0P0aQv6VGKGA2qJ1Z3TkEORNV
3K3t+aapH5vFxLHV+YzGIUjObLjXzCDEIjKNJyYBxhLmPvAKDsMk22AIic7SNd+Bgf4xsL9MWw5K
7rrZ29Zhtg+/PW/29z3urSL1y8emsvtW7eJdbMotXV6WmA+oyo6Lw1NR/yoQd+k+Enoa83nv+3/V
XkfriEROzjlXZFMcOtQljVnzv0K3DFBrEI/AStBdx4I4X07WtlBu0vzcRhH1u/Q5c8HNjfK6wnz0
J7V6kXa9cfTFt6ERE1Gm6O6r68sCjb7E6BNZa7HKWN/VyzTX/po2SJ6sHty6Yn0JrANTsRlOIdOZ
RBa8qQv0kCipL+DBoPC4M30Rwoy7LE8ciOp3ODUFeKLYTTF0xcWihGYUCdQ2CIEjH7E2agaxyQwZ
k4r5zeMFuy8h7d5oumm5PR3UVi8qG4pC8k5HrX8bYxT2AYvFRToclqzS26ngS70/Y9SL13OX98kQ
Gk1jIyEahQwVyJEJfpDpAh87RNs2ePQC0QNcb3w4rIwOImVpPI/tcG+8+l0fKh9qDDhS/NAvKC+z
BXMLTK2sSLpIlADp6M2oJUL0dHxFEMwiV0OB7dCZrwNiz3dDCR1XHThIbQWp7VxuQGk0QPYGaUZ1
7nplN2jptWXccgRu+8O8pPmikgIqz6C7aHcsJLyW7vpjIs6lk/9ZPmretAp3H6HfpU6duofHMgzC
Z/jF6KDKGYDhcBcS5Vjsc/TgB2kqoTdfFnnwI3ee4P7wlHDawRrWMbJfbAEtM16Egn0Gm6zyyhZZ
IZdYmgh9C4f3Lnr7k2GE1J+bCpOdfNDM8NUEpP2INkWmWzHzvEDnZU1AjJWlxryZdzqz+OcIpgXa
crZsKZ/Wyfudj7tbcYQTpKG7xDgUQJaLc+CGpuXFJVfhcXze3PNyzCA39CVE8bZ/8Aq+/KGf1ed0
sfqyhFt7U5F5Q3crBT0+uXyo9mvcqmSkAE3eLq4BkM7ZCXe2ZPUE5x9JJ2KO0YPrN+CohqnQXm7v
wq7skrA7RkKa7okxK82CQKuX6qtYf6VG+O19paJGkrehXW/9AgsfaJwcIewU2izhwUfALO7X26Lb
IXDqGzmxcKD+ky0ixBLu/cAvQUDEpDasA5Nw2nH+YVMVSzZiL1Z1afwx7v8VCIkh4UniyWcElh1v
PTCNSA6Ka4bGHBuqIgRyODgKzt5qlzuMkg4EC8VTlHWd718NmKK+UG0Kt7JCecqm6FW4BFJkKjEm
4qbVmbw45AesGILZVYXF4BjO0XAxllhlJ6+C34xfCKEyzkXs6DvcVhTkJ0ltDYvHYKAREXWKhhT/
Pax/ONbWoYO1ny8VeqcvcyZOAe0D/To3XcI3SYnyVL2zJkkKn4stqPb59nYoiAhxLs2Kvm31y2XY
vd9vXkdp7PRPT52EI4g0zWxJlfQm868vUNvm36/kwRU+FyuZ38nIp/fe29VHO6c/APSiLrc4z/VL
vsomKtZ36vjmYz5HhZqIFvsgvC/1E1LPViPHBCfYIEOwnAS3VCO14PiTh8ARLUAp1BiOO4XBOhW6
ZtzRUXC9BIOczRAyrIYWakFcZ+IE8tX5sR59rYJ8Fdht+G4ji/3efXdjF+fhkNIdM5KxaaaWgyky
4fCH0rS0KrKBrPW7/ay4sQHO2vndQpFAmej9vtNzzo6F/J0JQgw/iTOF6XQi3ws2FeVFXLx6i3JN
tauatu1pOeqy5EszjSHVnc7qNAOOtLANT/ozkiV53VrUo37Q+DLBaXpI2uJ8aWD3UlwXX7LsSJzk
9YTNBjSMxY4jjm9dMyhJvK6UvMXrF4vfbHl0L1Ak9PzAASwqYKB9/IqpdVwaywIgC5SrPr5ZirBL
l5mt033JHtwMh/D4F1oObi+WdYsATjRfyCNgpiUKCfm7MZpvxWQ2Op3tf2d+nBQss3sp9wz2ex4W
2i4m/vs6Z2+Nb2bGJ9BkEhAMM1KBTlgpnCOwcaBgmUXNFSvoEMDQWzlog08LP2qh0jHAz3fvHbCX
/jTUtI3mOQlJBZPDdFb3T2UAp7jR+yIlPYEAu2h2o/Y84Si1QXAopMOsDtXRH51cQlDx2wOnseO6
N4p6R916sjcO6ycfyGselyObsuHI8uTmS/VxmKACiQRwUZ2II9WNcNA9FXANRAxTTNA/UcvM65nC
GXYUD+pNurAMt/y+SofS0brNWWT5VqDxT+I33JWDR/d9eFrzuOSgU3klSEeOQY5kFkedPijLhJkm
SdgUFpRX/cw3IXZuNYtS9o2FbFViPHx4PJKRWmmNRh2Iv3ZegmYGDQ4lKh5NAvrqYITsSMmUovtp
+lo+naAO6To+o5DpFVvfMhGCQNORen70KSpqmgwFrI03UQM+G3dgDmPb/Sfr+iO3LlQ0a0TCOofo
/3X5eQBTxWNelrW9nkUVpXdDpsKGMkSAvdqrjH7mbPeOdewE2qCvu0zw9PSUg/M3odPgVF+pQpx0
izvlkjWcE/KlT05KfGXnC/+WWeXQ9HwLnKvkwyG66XuhC8SnAg1l8zCHCuimRSsdUxsSPLZ6O1Kx
GLlR/F2qNUQUz2hXn+Gx+9gvxG3yNeFaRYmqFrRoUfP8xiO2VfwhT11zPHeiau8EKp4PBBKEjbJb
OlSvu/vc3+7x91v23BQWbSfVfmXp8tpLXPpPmCg3Nxu6GkRkclVTias4ICBx/7vOiZQNaeoYDKQc
BzB6RjfEmroeR80xSzmbrL+SlaiOsXEIS+gggLCCjLx3FV3kQsrTcEa1RYLHpINvNqEAHvusA5lh
7FCji1Ut6o5xb2lQ+9ULGaaOBu29KrxkEVLy+gOJyjnWdx6d1th6bMno52qFbKcQ+GmSB6qxA1tY
x1uTIAtvYdNgw81+WZ0i6GlX/Fmn2KUqGSgC1hoFqnw0is2PdSnRBtcu0vjgXTQXijOA+OQ27Yuv
os4mgALiYiCOvBLJE5wSB5GGvuu1VD1cpQFpeR/P8t1+25/oknRb79/GdkgXS+GTmXhpZqVRvB6R
Tzi5kpmJq2w/ZHia9U+ur26OR2BeZYQIRRLMk5QC30si059IsD0XucaZcrZiwoaN7cmhGFZBoPYo
pfNdyO72H7KAe7EraV4yF1ncWs83QBZMG4KdgorB0mda0xt+mH7JGAd+DAgNHge1d7bz6JUhVE5W
YnyZUmSRqjhNu2dSvh9KK3bwnVmVrVjewGwPShfl9r4Wxu9TCNBcempH6L7ciJ+BFVm21L4d+WfM
kZqEPmUv0uNxmeggQU/oHOZ7jbKKFpPGDnDuSnHVq7t0oQAyWzU7YmaCAmAEF9NgJXI14E4M56HL
0yxpSOk15/obx6HPtdPQGojR7rm8LYS03uk6A0coRZYwmd/1RDl0kjNI5p5+VR2POJOpfTKNQNdS
VAUGaYSak1y/hFEWVtcqgT3ZMXhWgYG1Xvmgp+r8WjHQab1V2oG5q07YAUI68aCuX1WcxYFVm5RY
d+/zqh9qv68LfSwrC/JJIgqdWCBnuDH99o74bhMVwMsDIx7D4oOBJ7dDuIFStjO/Te0phVwrfLEr
YVxCgS6GGPWym5by7ajiqj5XjjWPr4XvsUbPpF07WAn1baDWA+B1LM3UDVtjlNclmR+arN3zf2+i
z/uF8FoNcWKbEC+PM8QEMBDTuO+WAqgyyrM82o0tlmRlDa+WEguAoaSGsT1ULxyQp79pcqN4SdtA
oBl8VnVkF/iEM6xqQrVLbBd8Elsk3+1wcsrAHgpUS7/QAGD5CHSTnXnxQoTfyY5vWF9wVMEpHpaP
KtFLEfQ6nUXen2mMc2NZ5w8NoC15NOCxbAEJgR/eQfO3+DMti3qsAYYlypV5Ceot0Nn22v0B0fd1
W/iwxKQ4w/jZerGo9u7sn36zNKgkKSFEt2DyGpPJ7JD1WauLYY+HkVtmmIAWrtvSVgfSzEj7TJa9
fClw6C4cE2IJ+0FEYgDBnmUIgm4vyxfdIT0lZQXlz22ZBJp5ljfm0SabBalT14I+HyT9z1piXyi9
Sdx0KQpe1IEzKZtNvtrtQsMMTMK2ba9Wz9HUzt+S+Ax5XaqDOtfWH4C+fQcyeBIKP/uODt81oLtu
dtkHmUhlkxlgLmbxQYnLmXchn06yw25nE+7Y+c5gV2Bbl+rkww6KcMl2NvsOWQ4WmxheqrVKutI6
AGFjb3jCILcqp6HkPUnLXTR1XwbUDbgRpCmly+yHd2Bygoo8Pl1AueiVFweLFWBcNndKkOszNggd
wFp5MiYXDJbeVw+2ig45sgBRY9lp26n9TxP8+N6MB8zDtEK2d/g4tpOrwPkDqZEqUFk4lV9FGb1Y
sLZOltdyfOw2D9Z+2Jqvw30fBHc1ytUg2mdY4VsH+guMsP5EEvVmAOoRa2dlTyhUvjeKZ/PGM7rS
mvru3Al1Foc/KqDfS870UPzVKtxRN0EkL+GqsY+RyE77InCVVjzKh3LatO5s2Uo1TP9QRsKWX6dF
f0h0oVmPRz9WunK5NYfyLr38s/kt1u4vci+ia/HAwFuXm+5EnGoerFTB6uKBBJGKSCjVqO7zbbSM
mCRelPmZzVAT8KgdK1BihQN2XP4yHA8y6z5yWvPmcqHaPsvIWaTcLwuowGedrVZ73oowb2m+A0qv
ddC7YrDWwCqMnLTRk6QJr9V8MYC+NKjFVn1B5FCABNc+sOA6pfYpQRHzLVmsrfp5eeJhtritcd8Y
T+4IxkVwiIp9MWLSw9gplIR0hCdkR6BqlDDAjd23Ig5QNL6ikGPHhe3jbNvLR53RYab2qj7Wirze
StXEyBvBuev/0eYKUQdOVVYzOVEGlzC2zCiD6XRwakJKet6DUctzgF6tjwbppDZDlCtXMKUGvzqQ
d1eWNrt8gu5lHw7rBvUY2fdSDKDSYS+E73o/1pd17yyKcDGZRzVX7PYSwLvR5umRdyA9KUe4C3y0
fSwG8TX0mLAT/iKCbJmuaeYmgeoe0hhZiYGJlMjFGKOJ0tgOpqCJ59KK3ndDfjjc5YLxc4oKO1nA
LouJLvInq41u8aDPo5j9Rx2fNrJKaGeDCY9XKNi3ikhnJDtbGcAWjYjsr1J7hHkxRurDqviPZpbY
62o/Lj/3lrFBroVMt21uC+keuw9KwrwIZGwoOsChWCxkkO1thzeLveAGrYdMpsXU0K5l+hmucLxP
WMXu+JnTPYnYD83F5hPzmLTkoS6wxOvfpTXx+6k4fkG0Mv2UzeY1Oj3qD43b8+aYy3kjeVxyrjl9
YDm02IiRe963/9wTB8l9gK1OpTetB3p+wr2ReORmmIPtK3bk6kFXAO2oWjYE1vx+kyuICrJEHpzY
slYDI1e5/0YEG0PjXP3wFzo1CdpDBbIit9FaXKeMzQWzUzkfCkG+brmo+oB7t/NsHAJz6q41yT/J
kdg+CjHlOU/x3po/bXs7QV5yq5sXYsiONqoLXUU/28fhrARzlsQ14nTK/kaJ47oA43bVlFcmlf8f
QbzwYaxHfYcy9Cuw/Y3qTFAqVCIYgzbGNSbQtalRZOy5DQGaXx3EPEC/h5Ts5U96mlxF5wzXatHQ
Qe/91V7M3DMthNOjHB+SOiCmHeXLR2e+a2HJM0AfoYyRKSoUvgJituRH6BCPgu4u47WQ9p10zRVx
HDEYNAo1vuZxyUJDAUpONK70CYHQu0vpp9DvfFw+5U75ZA18xoveZIWkSNykYzAu+E3/waoRczvR
oGUw9y+rEcBU2kHgwAF3EL64ya9UmouYL8R7+PwT6bGmE4QOq8M61cIBiasvgJj8qNK5ybHsM/6k
L0kXvFmlLs8uTyJmOclmS99oB0aWDIX0rExk6zJwpJ6950qxeC+JKepKmBQonWPv0ZNZHBgg9xuy
qQYfXqsRZ/E799Z7las0ySd9XbZ/KQy4rYX9WNJpGgKxgyeGQteq0KYtQ5NVFcCUe+nbdhosaTEl
4XaYAkSRuRAOmaa4gVHowsVBwQWQhbi5B1h9sUh6NQOZZjYp+IZbZnUEIzZNOwukV0VTD3SwOGyG
5kAWDHZ1OhUe+JWmYSLqg2mhPi9T4iKn4qvFBpbINcCUoqBsrROCe1wNa4ERbGs0i5MgovgnsX1e
Z8DZh9APvNlMz2U9XcpTTcngRbi3Y2XzRalx243G7h6i7J2QZpy97EgUEKiCW9B+cZIoiNYs1jA2
hhdE7PDPAnCb09ojcsuAL5jn9euSfhxz0fLQviKG9DaLfo/akEL1INfPWgOCy5W9LaKTAh/pZCv7
zvCM2O9zxGH3l70QKW2Ko7stUvaML9cKVh2gCw3E7Scnh5SlbGNrgMRsMP/KQD7EkoyWuCgnvbgl
1dxFkFeswULa8cQyq21ybYDW0z5In1rZ/ZDyGTkJJD9Ft0kByGWAKOUR+0l2uuEnupLYoiJIkrDi
gxaQMITIznRVHqHTFlZSXQ7SxIQkC1hl3O4SxxFIKTxx1c+3RLadLOqglSzEaDqHe314i0pNoQ5v
bpZKDLsk1kdDHqiUrq6qCQSh7xais0eAnJhZjcfrS2AtZznQ9PRm+wEaZtVe0MvgQ6/EOxA3+bda
Hy6e7JwvL7O0xL0ylVunJzVtG8uiHVSocqpZQzcvGH9/OxSpNFkeNNW7ngXqOpSmD92Q35kRzUvK
bIWM9xoDHcWQJUgFEpaBHF7aoFJzGs5TU5HxAtE/S23+gEjMI2iqW5Lt+R+NebTc43yydLyi7owU
zMkBCfoLk1TmZkQhcGT3P2bBV8DPRegWWL8Da15a3yqiVomqaCJZq/9wq2V3pPZBJJ3+aBZ4AksU
3Nslc/RmCS7XqhlCT9uxhAJjxkDtAWi2SPVu2CvFfwUZsEAlAco7Pag7i3Cr6x4ZImvxI+u/Wkrs
a6VNvdV98BllFH33Djt7ItzDm90fvCCXaFpcFElctpvHnpJnRhVZ2LYrZSFB2/+4pKByRnwAi+ss
FwCzqTGhyMkiIdUOK/k8lU2VsDeXkT6rQIYO47i4JQywXOPIbAkyZ5d/YqPV2XByvFJTyIWy0XIw
5qK/o4+M0YVjxyYbiIieM81zYxSvfY880Uc3AHjDL20iPTkAcKwG10dHUe95AAdKcCc+/YC5yr6q
+ZXPePO3+pZGaZrrOCSQoMxsiHvGbFXN9sQIUFQ0PfEpFimLiS2UQJ9aCrZT6rlTF4HuWd7wZ++A
PvcKhb7k9WmQ113+ZRVq8EQpMK1HdtxAz/9IV4Zu2CUbVrFUT/dRpnumwQFKt7kEbx/wdmfRlzeg
79hSJ0u2hZshxUGMgPMGpDkRe5EoUwKtgFHpRnLtFLgXoIUoTHH5kYx1lWaRh2oKP7zjTdwdAaO9
w0mnTI219BnWkduOTeqYq2+tkIxEKv8Bwfb4EmkbNLRw3Sxam244UvdF49iuUTmAaT5s3rI8+2ya
/cVRSQoYBtIKwJpLU8GXWSNNrqr/TYRmQLadPJRuKXJumNxadsTzBbyNdzrw4+YqyufD/p49rWXB
SwGxwlioW8krvDp6BraFqtiNCt/PrAcxB6JAY2apr2OfGzuaxm00IBuhflhj3qx2zuwhNRspWWMc
WvFY2lWq43U1vxx0iptSGS8L46nP0Z+RUpK2taWcnKxfT3jBtrQ6fp4rKVSQx2rthS6gpCkRFtZh
9jjciznx6ajpVoHp6NcTp/7Qcwa1/ZBAIzvMlKMCwHw8kAqPRVqBSO2E6+H0NgzIRW9Q8jIxUGk4
at+3q6H/KJnoOfG8y/JZOYT8pJTBMhN2VT+Ogkb6QA17YWcKJH3ejk5FRFXMOsE+vIYLFi0DQfWj
GSu+YQQcznp4AcsgvJ/ERFzTGsp8sGChm1cT0htYsgMSnbBTXG6+zDkOcXDf2JXBcKf31nTiXGQ5
cTH4gTIvKRvPj2AYdD42IBnlRFDlB1sb8G7RcCZNHe2Ye7rJP4WK4F/Stxzk7nBgpJHVuxyQavL9
TjES/YrfWnjVSB5h+cdJgPEjzvEmzloc5DfjqSwhPfrNwP1GYasJf7whikKFL9fDjE3JrGA5/1DK
0X6+rl85Iz8UPElU4OR7FcuXJEV0mmbnYBP+DFnOmkD83FOZIh0IBMGAXVOE3ww0rkqXqWhGxGbh
lufOPCnGzbVUVRr5v2Z/X3IFzmF+x6lnk+0K77uzXxAdIy8i8f+zZTNAuiR0/hzHvKGpGxIuJBzC
zWqkaQBssHZ9IRJ11bvpgMhKpUfiJy7rvgvl9r4D/3Rpnf+6Jd/XodXyC4//bgw8QxfOlYCR5U8H
snG5NF99L9dEyMF0MjjltkGDYOuyrnH/ZIgjgdyVeeWsOAjt4sozytyMwqPtiAu3GSL7K37wNwcs
DtfU43f+dbAjIga8t4poccVSiC2PglkQ738jJERy5NloPMR/UUmThLHv3Jumv+fW5uNNyzgLizyx
5T2qLBF+XQFT/LCTWtSIrIFnFH4xdig/0DYXeeOlHMbbJdbhpFYJsS/W1s+bTMGSL6YLCfzldSD2
/JiICS8T4fYv5WbKJMrrfFIr6ou8kyPOxkCqJlQukAAt4ESbAPMyP4NENEQTk7KD251Dyv4u9roL
7U63sr06phWSuqjBkoRcCizAZ0NEWGMl1PRf6jirC0eu+IiZfb/kR5m4kXbv1zVXmAxmz9BC5h5U
Ra+8YIL1XOHjgJsrjZ11RTNihuxH4lRub49a6xIcT7WnZTdPyhZUN/ZPNvlrLHIqci+lyz9/EhR2
pfI8SQVJ4XxSNLK632ce4Z3FyZsSEZu81mgsXbvN7AYBSXRzzAmuf7GSutoNDXWg+EDxGHN0+yXw
t1EMOhjODQ5oQGkbjHPW8HqanYaB7psHu1qP3Ok7JAgi6ktYzmu+A2qiHaaolRj31Yew/bCB5EE7
L9T0xn8wLikuHulFzY9lNqFsfnPXiXcK4LGfa/RpP5G1SQWohNmdJpMxQRodrQXQq9/e2ZktcDNx
rmszGt4kE86kcbzrnrKJsw9yKILqYjMSSmuhQoWVVMWwt64nQdw6vAlaM7UXfvVZbuEAZ11ONEtw
wSsQHXUKL1pKI+2F0xkJ9XHSY3BNIxjmzqcgL11QBr4rqQ2IAgNXmB+X9H7sfFCsVfCJ1EPLLBjc
8X17//zNopGYd1MohXFDpg2wsIKPrqhImoabgvCsvHejpSEWFHwZgA31kyXuChtMsNngUna0LOlJ
WJOUQOtSeVW0/xjJIzL55QQewcM0t3WTcPJyThHO4/pGmR71Acagveh/e3UnGhpXkVL2/FtnlCdQ
xHJViBiXH2KnnVDVZGxcIzioXoa6eTqTaF1O0m7MZEhx99oyNZlAzN89zeqXo1YeYmTCmuCuTnPq
YIWRsVSq4Cfub9xArjAORiGjw7KQ3G1xCFjAlH4aiL7sg7+DwWv+NvO/xYRMILXaSL2Ij2p8QK7l
9TpKqcemcEKAzjYP8cJSOIbP+Ifq27oTfCssLBIK76fVZlVHAR3qfeWaGFdmAX6q9BtGpXizgsB+
5tZRCFgiYSCKRUShLbcigld4ox42Y4ixnJIR6aNvw502h/SF6zIo7ysEeYQKNXq+TflN+ZIig07t
QZ+KjxgRmYnyQpJRv/+OosvdU3wG0Q96uSrcKMtVtJcKun7c1TX3JfJPwwUzeghpmC8O1b76+N4A
TLCZZY16dueYpoxr3rqe++a+zPqEUSOycAGMI/mjQFMwX36Oi8QUo+yR6Kca908DVHHsbOoIpjMz
aO8Mm5eEj3XAJ5BqTLfsTC3Sv/Kb5cLEvLAoY2Is9QDhnalhdRXwv9v/jmJpriqPX6yAq36/paei
vlrBIFkHbk+Wt7VQGnNMHFLG3bm1FFdL0rnTmkTKwtBtJtTkg7GXeynHj3gxgtQJrJhF/F4hHTLG
w7l9q/E56kyvpQDtiEMIhcM1OJq82Eey6bqpgSYrPj3z0hhvEVJ79oUDt5rxb5gjuytGGd4hl5ju
kdkZ6Zxm4G7qLbumQL0/qJhV/MsWtksKMuybpDS6VqD5JTQNUvRAZZGtcHt96Fa2bWOJKJ2r5Gfl
SH5FJfvMYZTRAyCepsI8j/7JawN/7aa9+mJlwIDsBAMrT3hyNE3bPocZfJrZ9Im+OcF25k1ZIdwD
a0j8jAz8OqJdDs8SY4ULYVI+1Sw2dyYJ/g7RnvjGVynYdSNKDYYe0+p26Q+dR6/e8dwDCEdHsBgF
FJDyn/C2gk158afsIfNrH782p0oqR6trmcZPPhIo4GgFqEfZzd8pSzMJ/LdzH/wJ0GqrDVWODBnc
057KpVTKvNoBsfCTHr9GqnOu2bvho+v8+EAIlms1O+6X6/CzZVwfTxUqqrcEQ0A+QfttR+YmfCVR
M13ooVQfFyka+f+FOy4kLxkO/W4L8kewUqvDcz8htZDF+Zuy+qWbL6byIjBCONWL5M5L805Za9Wr
4VH+rRysG2X7y5SEkLkHJw0CwCWYNH76ilC3xcU67RGdR9VXFvzotVSPjlkIdX+KZeQ4fBRihps2
FWTzO4fVdg3DmlfSoEYhnlL8+d7CRS70Ni3LB3OUjP5Lp0xIZMhNPSsnu2ZDfN1jQjC3lqaeFscZ
o5FtFtH+P3gLSsVS3L5niOA4gUdEucdAH4FCj5mzok7C9JYGtPcgTNM1Y5P/aVrAhFa1EwtAcyjd
Jz9n/LCYLcY+wcZGNduGx9duH8pfw8qcClwodRkC0iHk6idHR47xlMXuT+1QNN39nEd1JFQ7fTEe
JU0/v9/Oe2NHnQvDklR90DMRp6DVFkm7spSjpcgZFWLHvUFrCE4ucy8XUz5Z/GarxVdxktw7nI12
nmDPeRacDoPYkIOPMc2vg54Oua4qW5UpUvmXouuAFCdCdgae6mx0UJXRefW6kLl4VOTPx6ce/yve
6WC5e3tf+xyY8JYPeAwUgh2Nl/zdi3E2B9ZnsVhpmwwuzziIdXkXSQNkwt1N0lLy+N02hBHhpOkM
CnjLc3AIAwvTYPbb7e4WqmwoXAQme7nxfgFstQLd0ktlxIPpPbY8WtjBGsjofUTHkuMWU5Y4vV6x
sbx2Ijlip0Y+2HLsZgJ8YEauRvQdYVdSksqBEXoCLiM9IuJYNMb3JN5XBAdnpYDHx0REkzrS00Fn
+WtM3v/I4G0huQgNVqc4P5ylIgMTfisiI7OI6SjoRKP/o7RvSaMgwdNxNESm/9WDkc46ozVIzp/B
enJ/kopmNwd3y4xbalPtBFf0NarFc8rNxZeHUgee9jGgNf4jPCmMlAGhFIQzC4ry/wtWD+bsA4U7
NQS+P4uZpaMJgwq9WvnGD7sC98hbYpcomX/eWg8xwOXukJYpPbpjktZnJNeNXusxHppcPkRp7i5t
L3sR+B1k2FDVcXck7r/d5ZgBMpjYdqtZCiGyr/ziGvtkd1gO4xNr+adDX1+OZYqp2mCnKDTtm2tn
MIPjM7DqsYGufIAJJUxRjJI772aG5c1mat+2FeO+rJgAwIPrcowdbTlBX79cxQ5Q2PQhL266kKwy
WGcq6bCAWRbecFVyeCkm52VIcWKMfGIBVtN/ElgsIJ6Xbm3+0RutsvKnNQm4npDdbn47dtwLBd7G
NgzWuLXmblmPal4kWWs1Dxzu0YsHlzpBXVGLZ7VjxI+vbgre4jMiFD3warslRTy/mBPk2T3UBdgF
p8sgxEbCaptswe0WcvlgMD6wMP8v+8FqggFCSJuk2Y5Geyo8kuBOhzdvtpsHpsp7eoptoxozFZzD
Wb08wwhm4K9u9x1xscTq4gi38tuNKY96CN7A6QkGyie01MKwxUtvVT9eyh4vuHyNTAdlKiCakf4G
BWFN8oXSB/Ycsn9Az+e/Ph0iNUkH8GcvUvwwLtKClclI9HrwdmIwf8Vu7tMvQ73FELc2iJOdGVGK
U0JFe7Fnefiuoo1rjqxo3My0wdpvoM8gpqQw6OqRfr5Eqr0B/dYXemXjjHVgGU9w5bn0AZ+Uoxlc
jR4VIMRUCh35G4GP4FKXOknuZgkxdoW+4/qLbAzeSZ2Tr80rs94PF45e9X47bqLf1GQiAGb9UWvc
u6lkjrzR9TkqTYbOCadBZ94ZJVwlNyypyV6aqwWFt7E/d6UeILWUkuNzh5bX81ErfiyY82t4hmVN
+uMu41fut+Isq6iQHscfBrfKFrw+Ro257e4rQ+/6TNu9rkqwtQxYx6KhhoHKaXXeFygF5jUmMyQ9
xOZUm8N2t5YDiP1lD3Iih37YfhjVpPwxam+WIfLvKmIUPxWrKAgjSO90DrDqCLRfrxAa9hkr/3H2
C/5ZKtNwuW2owXlYZa+G+/zsLb3uMH78JmTmtEIxg7TWXc4kAxGP6abmdq9y+YpaxWisK14lJe2q
F8htEDDShZMPe1jR86O/nEpbvI2+vqIvoTzThUALmhH3dz6uk8+X34MJSeNLHmZddzSxy5VqwWD2
YnOXRdyENCJV0p6FfYOIv1Sjhv9IBz13jojQ0BoDJLRjMQiLGrUQcCOKldKUNgb1EP2JbgQnUOlf
71NvlrGs5DHIqmK0UnpTbz1sxWrcfmPQ1c/HUTO9H/qE8GYcwlLu62Ic0g2hAgVwgSmPqlrhxrvI
+iBlswIBXFJ5F8UseBS57nEnH1Pev2WpyohVO3Aw0Czghl6H34ZI3jO7U1G63ZLBDad3siOeL+zZ
OF0T76F67MXFZrbdgDEOAKFkxDF1b2J2rbVw56j8tJea7A9GgeGuziH7RH+5O7HsyspKoknuZ3ni
OgeR8+YHbCXkOm10dMXWCXXBmaOKfflyfXh7IETZgcQ9ugOgQW4hmeyqXU7oE9RYyLin8g3n0No9
SmPEZWiztlwxvzBb2qm1Nklb817mTwJ8KNJT2LTvoLqO9TAtXciLGmjxa7ghZKrMx3S+nXJdRFJ4
CQTK/FqBum1nT0l50umrKtRcI2pmjmB1noTTm5FXDnohrtgkxEmvPr42Vz9PVZptn5YBx2NDoVdR
RkxqlUO2qi/sGmQmH6caB+AUw0l7Lh8I6TA4hExCf2Sem3Dbi2UUAbC0xL3eq4KidPTPn29VJjXC
ycKbMJsmQJ9hqWiPgZHzI+qnmRyJZceQ4Hv9J+oVIXesIyrzvouhowEz+ZcsOp6+e871EMD0Yxha
vIQRYP7K4ao0t+htv0MjCT/0vJUERbzwv3R+JJ4Wt3kxTMXk3zMNNvccAsWvY8+A+RH4kRO8sRkz
xN120wHvL+QqPzwUa9AcLFp8CoF6SLQPwMoVIVi8Av3Ed94+zlAfIG64QtaQFAE/KVND5F34dn5Q
ah3yVx0y01+Vuhfr/ytHSvyrja+eIlU0eh3sOXdULfDDVr4AkPDVovfXBjtci/cC/D8cJQIDl6AJ
j6kIZIk/lMBhXLF1OGYKU6+vHNqg6xn8+G3v/8kq0SOLgcEdpN1gEQBfAOpf56y2CV5ofghThrAm
iP31vvj/eBy6WRzlo+IKVwv2Z9ly0MF6B2UA6iWiHFojQslzQVT0DHYrO5JcNeAiTHcLqTLTAW6V
s2IVPGNBqS/otuQhqJPRraa+GiXzApq4N2uSch5FWv0lLINU4uLNSJ/Hnzy9S3tmKfHHcD6c0XSS
fckGyPEOmex448hOh9ksptKiREDyh8+y5LXKj51AhJLBNRmBD9wNuNoeljKxoepZb2TgVSEhQfp2
mIrU9d/z6HpSCYY80vhBMQaUQuD7IxKh6+/hnR94me0bmr2VnVW1atbcz7sSlVdKf39K9zn9zBb6
8c8do0wFS8ZqWYE9J+MdCmNQs6UISHq74H2uDlRVSyach0UuojgVIs8KVteeccL7myc/HHiiouis
Isq/nmtttZ/4/AmeLNSl2M4Z5VRsOCX7TWkwwb5MMcJQ4htXvNV/RVVgELhwlXLrCB0DRxNa+rc8
UZFbOfyGdb5YCnLvGz1o0wNaVSFS1gy0x0LNDezMAd8dHXFQG3E8ykzkN9jo51zj3CnMOqdiNuET
bU7QUcVY65UXeUuhJ3vbmkSApI7lUhcLAM/AbcVofCqoWdcYiqMTizh0iYjYj+20bizxnh1zV/FF
sDcVspWdP1XN6LCvSLv16kiyR/SqyIeio6Rn4llDqx57sYCPC8HOGpry7Oveub+Gc5RwuObffhQw
+RxKQC84ofeqXl7Bh96Ca0vwfXdChCHq32yxD05WStUM6NeJrFVbZ0xLbhx1dOLZEeRWdDTTNATb
uj4lj/JFdJzZrwWUKu6yOwQcTJuvVKNiUqzJRC4lDXe3Cf0unK3wBEG5TnN5YvsFcs6Unz5+GwnH
dHWsDSwS0txXapTClzApHBwW/DP3311WlQyLGCtpzcW3S+nCSxkg8aJxMjF85Dw7NOsCkDH/qDNX
eZTjsWeSKGKrsNWKmKDqC/jwjw2UkkROSytSn+b1QlDeKMm2ywPaNVaEiVqkfcEBqHcu2Vb+DgrO
yGjMilV/7ObzVV/dKsOEvK9q4dsgA/xceoyYWLeVey2Pg9h2zZiQ2sN87cjKNSpenVLayIB2Io9J
4VQ4hRc0n56ayZPgEfuVA6CKjB5rYx/w1SepojOruCsZ7qqJrco/b5W/xrB5lpXCKHN6HfNnkTKC
Xori3tG8USMCO8pRTP6vYqSXHwI16RMG3BQZY2bUq895HiH+RG45oqJTGZFse4Be2RGvop9BYQ+Y
YCTY3YOM3ad2qSbDUYcuotGuaLL4rGME4jpHJS3sXu5skaF5QAl8KnR2YkZqMW59edmhG6os3GKE
DL9zLluDbV7hWqxTNtlFmcGEADxbWtBi7paEH4pFn0b0JF+noVhmZ5zr6b984cOYLLOdh3mTm0Ln
h08GWWJ3ie4zblsdilNkAk40PQ808eJSPcHPPGsyqFpMYkQzCL/UWQRbvHkVaMuUCKTk7bj3YkWV
HgRMMNujsfLWzPLD1nEKJvkWrg/BeYZghHMHglvm7WgHIYhEbUd208Woq+O2K/rQxg18qw9ezwTn
D/HJhG5tl1BSeYxv+7bSEigl1d7G4aCo6EVBXopUrF9HlZr2qYLb23NtpfIJAJn0Hr6H0tAivqpX
qYxhBvgoXDgqh8DxCozRRqTOOgTOQU2ekAFHnRrNwfq/6tEB5s7ELPdGfkEIH9QXm/i0U7oav5Ho
d1jUmS5cX5q8nolS/OGB/cYpT93nT8yaI7qdAHr/wxr6uFiUTptbxdZtgjxuENnm9m7ZQrwVnA+y
BXj1le9AefiPODYZJT/vFSTuvYfixLbeJAUNkrxzYGDg+5SEHY8dejRu/At+A609v9V61/8m1FTe
Pnc8Bz66pLp4DdUNOgZWA0Teqn9zCwlFO33TFnecdNvah9gXGeJ/Rs2wrV8oVKk5Jnr9GtEYyZaJ
S+eZwEqqPcrCblSRiLe2dKglaDaC/ALkIo9D0yb/rb3LGGNqVTh8ndMCmsviHAqSsB1IamF2mRDR
Lm9XbahtARpGEg03eWOn9YKLMcOfO0U7bosldblM28l+4CrB9pk+9Ph4mm70CHa4phkgzWqSy1wz
rjMb3WHtCN0uen+mdpT0s5t1SvaxFVBkqpUqJntxXNRKtV+45iVIksuttNw9Ge3OiIeHqb63tOoG
2vOYvyPHoEevgY7dOwnUQ+hWdnjjhnivCeIHeVkoQBKeGKLtmmaXKTvX45UulS+bzJuaKZxI5Azo
Q6OaB4y+5T5vw47RIr12QJrgc5Xpw72LrEmyF1a96NDCL3vk79fjVO3ZAE47j2LFfiMmw8J+iBAx
xdsvxyA7MZK9ZiKQ+wIvKiTqnrbFra5fZFsHjFZJNut4rBwOEEmN7wl+hxHzGzRGARvOakNtPscr
vlOldPi+yPbVBsK5hTO7X4ywVedoLwo16Rrc+g0tYz1B1QCy1eqsmxS0/wl4zzy3slqD+97SNjoO
jCa2NDhdiYlxkMlRRPbdJ5HRl53MijneS2pSkxKfjxrdpnAVXrxZPEF4PKu9HPRVCrgGOhxko8MT
Z9SH7bTjp1LY0K3gDLHj+5aoKO5BWlzSu5GPz8seUr0AZiGM69PFjTWuQ28ixlyS7s3x15MVOP3A
DQzV8KrmuPI8R06ESxhV6J8P5aT6h5kRJygPz/pBwdW01n8gun0nD/Y7KUtt54sBWviD6ZnQCKml
aNyN9p5dPeL6LofO6MpPanxpIsfgrdsB3d28LEs0dOdqJbJndtVdyvA4jmDZEfl5SdVTyUnzzrVR
Xh8IYA5Ms4GXebcXoqisdeJRDs0DwlaQWQPXpLrz8LZ/0JoR+xnAAQjR0qi8AESND4Ndd3Nqf8Bd
6jfw8Oz2kbga28qMTtXx0+4T48RCQL4mEIENxsaHm/99x2p41D+0TxFpkNdps7J5tn3iUcV6jHPC
uAggqOGqt3uuRPca0+j5Ql9yfhaQMnASylFcGfGleHWp2tIyhJDtlrQYaW32zMtfdWUOMUcaSzBU
NTFRAmyY6OHITSoqfbHOPHErlFI4wHpDKwTYqsaUc+uXSVvymQ58/APcFiMKB+HNUNF2t2DZSCZF
DTUSEdQqo1OQWk+/4fffJkmVJsPNmOdySodHQloNzcQ+Al4lxES14V4CFC1DDDfn0/rP4soTK3aH
WZUPdLEGGJcwRIf1dEnV/Fzu7IYQcZh5VHJjAjmW0GcNjON6SUd7xnXvwleiYjTRaPE9N0D5Apwb
ZE+HgrYkb/JwO+CisVK+MADHGumspik3DUso4PdPkHutuc0bD26nJ8SJ7V6GsP0jha64GZI8re8T
CgXnH/Y4p/2/wH5wz0qD36bfIlsM+BHODU5PY+XZcO5l9pM3s/ZcPtYS2e4cynZV41wur/toCXs9
FvfVi9t9iEBj7tUrvqtHmBSUT1N+olxOWHcINHOgzRHH5Yyoeu7kL9T2yQZtjnNSiCagY9ErsjYy
W9U3uSAYafpx3YruyJeT929Ofk+ixiGvIqubiwGnnjh80yLdO5gdUR4EXq/jm8KC6DQeSeQkGPJm
2Qr3/QSPYintjnZw5/B0GXqz/L6kWdhmJ6v+nLPbT/SxUbYNhRLo4TBauHj1nkp7cui/nf3zAvOT
+G1ULHrMJGOncSiPGbbabWbUn89z/RZ3BozVu0RGQeDl3ZThRQU9QOtIqYnBEgjQQwOrey0PFkMf
bpi6USRIXkEPu8V1tEi7K5V/fte3f8jOPI2qe8o3aKc6EEdoXTxIe1FQhpmvm6epXJbLfqpeEuJV
JOAoc+X/VjIuyFWh+NgPda4ZE5BoRnObE1D/nARRgzBlfHSTm/C3JJA/S3F0xcPOaQIlN3jvpmV9
krwEJPjPBqOpVHbMOK2fUFPROh51FWMksYktKr4p+3tojpUQbDsg6Z3WknefcsQvIKVBUhfxELCJ
kJ6ZX/NDfpoGNHdg4O0UJ+hLIaFrXrWNsl6PgCZ+cWK7n7Ix4MgVVQqRd9+pRY5Qb52QrpxzcTTC
tZV5k5WnVnK5n/slvIEQSg2EuG5pegt7oe9QaPJvx8tQEKevh9OdK1Y1l19+5b8Vtr/aT+ACawYZ
DkofFiH8Y0+Kg4xe/cbNtwgwqLknfofYRjwWBa3YJdsHY0FRN+pIQmBBFWzRPFFKeKF22W/TaesL
QiRT3sj2QtXrBUNlrRW5T0Vmp1ZAWwqe6Phlp2zjRXR2mIzmrNd+zOZiMwNLwq46XTZvubejdhn2
NSnai0Ex6NYjrwkTiLsTCjtiwd7OuZo34Vfdxs7pp5DpP7Flcb/TDGsuZcpWa3doO6BBQ34sJQQQ
cTQINIlTjeWFi394W4XALvh8zR07tTbNRmVJ1+RMyFI8SVx6Di+OFyjf7vwS4MqWmWKNeKI2a7sr
aXXeAkKstKuFnP3rugg1pKGWrFkNV/OF4Boiov817tEcMKUNuoUg7cpXFJibLiPw4VEGf6Di4Ydp
tfW9mYru1IPtRw2Qx6S/42etP3Sx4qXCQWxiX531pO9BRmrujVDyz2rd04FnO5KApuD0dvcS/H2I
JW5AhcJYU2TB+7C6u8G3o5B9qB1pVAwznjbQLWL2pW4PB+YUuZKN2YW2m16IwrDYG3InH6zjGFpn
Zyuqgjp39XkLIr2ACacb6QoHCPSS917+SMc+yAnL4lHK5zhZgQcnrsXPZn8wap90CPINhYFMNVcF
7SXqjV73CzYT7/0ZuxhgYnws4OOfovNcVAli1o4oAKpBw81RfI6u0ZC6dRuZUtB9jMJEW7DnBs1D
+PWMLtmyRhnMhBwqOIt0acUUCpwaPsp4c20eA09x7dywZabWeDGHRYBUdzw8tHFRPnsvmn8H4ZYv
j6uzaKXd0eoB2oB/DQE5YElgyAbvI1mkgqnfNy2DuA7ObRjm217PN5Sr4fukK1ID1SNbGDrdx+SK
Dq4YEATSawPLfcCgC9auazHWxYtwGqDTPhxfJ1mmXbPpby6X4mB4DVoVEXpGRFzO7pj25cCToyJH
GqQl07e+HbscXrX52Eguxr+sSasMPsWWJVaKTxwt7J/dIu5a+x2o/sKABSrcp7tJlC7lHDQRgnl5
1cs9pu4Plx4i63j3s1oZ4XvHb7ity/UIDUhPjqIFft93MyxqFkofIQeGwSGVUolRYjz+MRrFEwFx
ITLGS2TPhZ7xUkX9E2fyh97jd84dW/qsPB+O+p6w2lbE+3lWOxBkeXvMRxMhZRXQ34DbRNRE8WiP
2bxjsgq52e9sGDq0pEfBjNDH3P2hvdPxFSiLamyTMwYBar1F6+4DeRfNM17CLiIFqAuV6klNz5qF
iAbl2z7Jz9WpbCUozrqFmB2oYTAAm47g863jd8m2jmj0ZB/OUUPXCzHB2XeOMqWqX2qCPmtuqaYU
JJyLySzFeulIx5P/Hj397vw+QWOUtouuyoXlkdqmzMNwAgFvPs4hpUEOTS7rzBD82yE6eDnsmDZr
rzdhohZSEAbkl9zc9AGNTxTsI+vVPdCNV04mEvEHypl/maGzavsGal5BUeHTSlCg2P11MPQXLnmF
oVxLS6Zwsh2TAJNAHzF1ckZ13P8ItEoiEGEjgO/TbwQRPOnStoHsAn9zXtRkf+A+m1vKlTUX6V5W
YsSkdtz0iaaK8lTFiG7h31jOjhabJ5aDdV0XgaAA9TIvIWckEszwOvReYkLu8ZLSITZvZcRQzHhd
fHoUO5XubLSP6CDvXs2sIXobovyyaRCB5dnROy7IaUc2g7dPf9yid+dRljoCKdcYyG6WBYUiKGE/
/JZXJbiK2xVyWfwqCYfvFCypzkt0w1jjSP0s3hXh04EORs2HN2UwSmXiRr9B8gPtFi5VDOEiRH5q
FfX2BIU5qjfONEKAtP/wLCoT7yFVugOPMEpLmawinbRC8g1W08I6FUJSUJamGIZl+gxxv0WS34KE
5hCVFazsabqvlVeaPw8aZVD4r6AJO32pd5T4c7crzpIZOmGIkiOU36x+w5AMge254mWqNey//x1v
smIi16li5ml5aZirw3SGLF2qfnxU5gKYqdgw84jQwqguY0nI3lbMoXZ0R+htMLtg72B5ApgbI+zd
eHacApx0GjC8gEA/KQ5TpOZjP7zbKy6ZcYW5luSe68R3uhtNAZD6yoifDG9YjlPXfhUEzSC4K+d4
OZGtVuC5MaSYZM/XSDv7ZmwiGYKcUe6/rxJ6jy1dE3w7iSA7XBfpjbf9aR9Xqjq/vfEbbDuXrIlv
IR+RQFKhWLeRWoVhH4HH7GyHtdtfi1K4mjroMHEhcrb9Hy9FJFBZ+1uNG14mp8/1lmvIwyB6yUZv
wSaRoNlZRl74dAHOjIYXU+Re6Br5TIJTEVI4IikNyqj0DIIjr+X0g5sNestlMZSyQ0z310c6YaJf
S47sL2/ahMMR1/jro17QcqCcFtClr9Mc4ON09v+RKPbhh9gvPV57Kocsa1RVxFeqZPwoqb8laMgc
4XFrAQ0lDnrWgyo2qpWYj0YuYLBrwpC/5A88m3kgetqJQ7+38FGQbTlZSYtMz7UYyKSdZzSeu4Ue
nfqJ+nGBkByVE5nXfhQLo0odR/JaUepDd6/4O2+4ksDEq4bpHzwLtafeB+x38zJntiuU/SkzQkJ3
Z6kDu98PI2Cipj2MTI8Q7KVGteedlPzXIdV40exqAPmPiILavWLF9RA2zFwVnpUfWm8SlR7e6BUI
N5TzzaHeVo7pqLudXnz7Q5OaRc2CoUaZaHPro1udZ8dwbbXKl0oe44rn73vhsYXp1TqIEmZpiIS+
cBzIR00ZVA07cklH9vPPcgEDO7p26UG6MSX7Zui1dgJUjo5q7DYaFnZi3c4ENHi7sGSI24fdmVll
R5X6GnQbvbc8yBGYxHFR3LSw34GncaZQIgyB+YHYJxUmACC0Hiy4Qjit6beVa4gMgRArIZWo48TD
NBS3B3pv/Up8+k8evi3Y+6E9kHtVLhZ6Q64RUsV4JRM8KXfBgl8N557ovcYS/ljNj5A1/To1KEyw
hMno97z+t9m2e30rpsZkOHiXoouq+MdOS3G0/KhGQzwyn5SZ5tBWfcD6hTUo3s2p+DmUe1s8Oekt
QuCYDtquJY6AXCVHlZWc5cbRbWrB1xExooGvz/Ss2eeNryzJuCbOrm2dvhfPRYhPL61KLTI8kds/
B8EUGFAVvOkd8+8/rF+EGS5srVtuEWAe87Ly40tk7svds0JgsLPIZ/IjAGciMjljmLY2ONj+U4oC
3ktbytSTVDdFH51YIbjGLycoiE7swHIuN4/7Lyl7mqRKQ+Ds+3z6DqQvGEuGzU0RQkALmmEJdEU1
9DiWem0ZuqZWfrcEI4YHdYlhl8w0CM7j58dbbhE2M9m/1/v/upS4c9G7yuajYlBpOEjkOwvLnil1
L0MgzxpBaY0zcK97boPGsLFhOnhxfD5s+aWwbF9eKEfab4bBXwhUBezbLreiAjW21O9mIT1jz1SJ
3eAGaKAU1uC9s7J9bYk4kRDWPWyJszvQAvVhCvHBKewHLeKV1sN0wH6zShJHJfS4vCbACVmhETQB
KYRBjF60SUCobkqVyk20JirvIsePBlBj61HYkGE0dokcvsJSEkC8KPKP0O3LAThbxKS/uiFKJVE2
UlCPhiTsB+ySfwrZSYQtdkt9hDsylRKd8cy1yO5xkH2xe7ZfeEpTXpYNdA4HEOOYE4Y1Sp46CIVL
HOolm8kRbjKEe6X2TCqtM69S/5cCuqBRa5UPD2UHnzLYfbf2Ab/qC2czb5956zXFcCKjPbyNMAaW
mSRqNCWh3Dkn7Vve+CNcIXTAmG4noqov3hPEb/tqgoXTezTWbSeQgOE0a3V2CDO508Ah+5bKl1yx
kKV7KWHsTWKxTCXBsEVErPmdj4yKNCRvG8DEkunIMQieMu++c2m+OkpwcK7MaSsJLZQJdA4Cawgc
fYFP4NvCrO+V7T+OcExisHl1egvoF4ng0h9rcqR2UPtFLD9VHPj/zqXsIc6+27T0QaSqhJgJk6RY
6kR0oMg6tQiVWJqBbAr5EN/6CBOo2hBZKwgiKVOWzDc9r3SMW6ESVEw45Ubto0/FRgb1kLr9rqgA
8T9PWVQ00VaZCrfULouoU60fgqyzs9oGMcgMbU3UjnZP4Jt7VVaiMdiYhH7Wm/9DLXBDGud2Fbmb
HB5ZOm5FfN2frrcSU7B/zDY2ZJEiH1VQp65vXmhmF8RWA7iyemCOzxSgA8Km1u7GSJ5g0892dcDA
Nc8JaFxA96R58p80V45ZW7LJDApTh1IImJqVu+T0Yb5ntatX0Lpr+7kpzkeb3nPYthzDRCYehWVE
d2XLQyYTK/++sEWhBNZ+6D2RuKSoX0Z7wpvjv1Q1H+C5zPd1+KnJPc0exQDCqRPPRiWjMuROKqP2
WfC/RdaPFnORYawvztE9MIruARAb89KtjWmBv0NSisnQBa3OK7Nhf7TS+RFEIsOjutyXwDAC6hGJ
yAJgpMcNKPEnCgbhWasFSZKBgaGnw+RkoCRyBQAna7fuN0zGBBKgGHfG2diLDiDqZ+WDmU+nGi1R
hPRc+vrLFXGejNpv5EfLCi679NZ+ivkGP3NXqhp0U1a8Vsi/8Bwr0B4yJsGxFqTv+5Ejo29gItls
r4ZS/mRGvo+6ZtOSm/i6hJZ4rQzZKxWirewqedLZTzvGJXKlrr/9V7xAriFuKcOexLOUOrcslsMD
liXDQX/yjCLcObWzdDhkg3UbK7eXKpUjZ0jvtz3+bmJJRSj0mVSkiI0Fwx+xQ+oTVHL91APPTamS
LbTJajAnyA8rng8Q/bch70JdwXC+wMnVUlOnRmLLWV+5b9HkSfdqrFbktDufDORz9YuX+reqCnvA
qBOp/5eTFnX09Wuw6C0PhWRuYFT6HR4feZ4ic5PeCv9ZPORI3rfMSPzOYmy1EZWr+59dz6Sy/pfy
1SB5bw7W6ZD2kNgKBImZJdKRWnSybR4pUvYwOCjvwRzWUbf7WhH+4LOLyCb7v7s/+bw/M7Y/CV90
gJj/Ro+adBZxNIsKyCWYrF7PaUNuJpHlh2Y/HtlRKgfXpu7ElWShqb1QIQNTibrvXWGAiB3C5BRo
Y7yZc9i/kKykT2gYMUCssAQcBJxspgNg/5Gw7chY1yf+dIFVgUCcCtft5pzUwqjl4/h/1dLemZDN
sk9dUxXNRdy0DKPi1rJg08pynD9vY7gd3Ag3LVj4GzoQ3k8g1V+jHTz3Gh/La8sCFef6drQ0pSiI
wO5s3fteGcP46pD6fQW3Htil/ytCpkYwTMFR8U5mEIW0T8U2+ciP5S6GrJd5J0UNKSBUxkGO2qzM
BZp2kJK3fr3L9osFioGLkNbUejXebkbNcQeYbZsRSPWTUBsoHu/PYeLJZijY9SCLgUGccUr3DAxw
+NHLM5KaIjI5QO/q0pfk+U3K0zxsv5yoHheHCId4KSPd0yqv2W7qGlMsXayScIJDYBb7qKTq+me6
xWpN0m3khnq3GzsXf9PTiwqBhfH8vBtNCzo1hvwhynQAXVnYUivjvb3YLcX6Z77gYzOHEesSXcIC
/sbH2s9VrmohJi4pvSgD72JLANsE9Ntrad6l3wZ62ca2EeX1lc04UOyvay/8Hzw3OZ7jF817lSW7
GHxUhYCUfB1wdqvUIe1jlLO4nrzEQDrozekfwWUHcsVI15mbmZhgDOcPhpLQbIewAHZcZprfAZty
wiWmB86j4MYGoLFvOCIrGEEZCVLZwbBQZf2RQp1cblEHN0qgZDM85dhIgDUb7z3W38BWMSRC0Rw8
PruSbp+wCC8GDK61YOmdvU2g+8AiQci7T1f1Fjg+T4E8ZFjnVyHO+9KntCrlAwOWV8Py92z8+nNN
PNcvL2Z1fkT7Zu3Ja/nSEJw8lW8dubNqPUCGKEdjRQ0AJpTbcoxecp3IBX55ddB586P80Z9Iqkmt
6KDoEPob6MsJtfYL1qIMSVZBF8x2Bxs9rAwQmAzmNG6sa+LT6thWWh/NtzlRrDQGh6dmKXW/k45b
/gYMs9BVuJUtuxylGmrDp6Gc5dyxJhmsk/9p7FXxetFQgk22xsJTN53u7NmxOsHDU5tqrWlHozGZ
MiRhwoaVuWaVOQgxYq/kbrvnxxG3ScNjDE6WBxp+ctZ1jdxnF5gcuNd7M6KWFrKCfFHVRKZVWqju
6sXEGLU7qJiHRRUx32zoxP5hztbSx0hcLsXkrc/mrfkT6vkr8iGrgVgJDRhI1sjc7OLktY9GLvUY
zT9QSXFW1t5tvtk6sXDGbRi1qfL2WAGxJDch0ncQsZ4uKjhWvEZy1Fdh404QoW0ZhBBddjp6JmJQ
hQ0SqifFEY/P4XF4SKhRNS1MCfOTOhOuicx8vZe+ePly0L99PPkqCuOa/aTatBFakU0JiQWSwQS1
fawVKDleDN6m2hKkCsl6BFvMaFQw1cwkXE5W8jzlgduZdoJCszYK4M9+K7fdcJFpN1K6HwKtvDqP
2i6BluKpsz7FkUJwDfpQLiXz0RJ/GqVBWkHYjJ/n3QIIuXOV7wpdRab3iUPTuxFLTb5uWF4VR5gq
ZFVBT72F8uFOFEenGWPp/D++gSsC7Q4FJbkZhneujzBEaEj5ea9WzSgEo2qRKH+ZJ5HTpUQ8gZ1N
Lz3HHUxGXF0riYOMaf2fj/p3Zc08fRABo41Ke5fq7tn0wktFT5OQB2pWsVIuwO2dbRSclVKknn1T
tBrkFLWfJ6qJWyUDTO6PRFw6aW9uFl8m8MWbx3VXUrUAjilPluFUGpAB2zZjSbBGEXu+WN4UTqRt
MLq31YyFkHUPqPW8qSx0+r/0dzlxewypvkjnCpUdYvHyk4Pxefq2v3okGDNmXkzrLSY+b8IGTKME
Zp56iz+D2XTcFWQJG9YXrQjXYAEXTWG78BMDb27V1693GxogASHm75QfD4SULI+JY01hYiBGEdXe
sV4gbWZ9vxug999ozZyPK3WylKWIKl4A7Trh9BJt5x2nWN7QXO15oSUFsC/t5isg/VbxthvF5QOI
kG2AzQNMHQOzGwMQxJVx2GnAo6//1tkvvDc5VmVD6OEaLMFt3uByToCnw9dAVBHOaNslpEBndG4+
f9sNEHoGOOZvFl9/CoO9Pe+w32CRiujRmF14F9GcFK7qpzobmEZNiJ5lYP4Ym26YYKxSHorjbBSe
klfnK9jg2SVDjQgbVY7OZvsfJibOH1YlPnOlxMfExTK0slURPbvxx6ow7escX5QM2YHHYGWE+5zT
Ae0uAsB9a+facX3l4SzwRRtbi+D6Le8//cAqArEliUB1U+bdBeHqjcQwgvlwee9sROiKagtNxj5b
gshA3Ri6QHRjhllzWBMMwlQLWcRh2vyTkSGCJ38pYs9XjQS2CpryAdqwoRg8Cqrub8Yk3RfRwQat
Tf1GJpm6dK2iBv/JNd40SXz05gfE/Fr37K+TjbCZ4EtaZKTeqy5jB5zaw/pD1lr6R7Mf7bXB4SeQ
Av8oAXu0yH6oJBnhVSECZH6g5dxCjTumXM+ZcI0qEfS6HKZPIl0GRipw8J5bIQoVXLWs1tyeAbUx
akl5B7JMmNj0kF9CWDu6nZl3DeBZSDg0eFS5FacnJyvm+XhTs4RjxZpudxlFzMsI81q+nkegzw3U
o41apTFEhf9S5iHuK4WMUsWYBW29bsGdvwUqut2pNp5JQzsAb+kQA1TCV+dfzBH5qR4A2Up+Cecm
TKDXB4CEzCUs1FFyKIGe4oow0qAPiCJF7wWIp8GZINVCZgFPuWTW5Dq+wcj9H2XCfsciZbuuSX/U
+eZESpEB3Ob/jOWb5gaN8aJFZVwXVMqsdW27XeeIIP65I8mwLnhc0Hx5wGq+CoNF6B0daOmluXfR
3nFGelUYSsg6OZujV29mx6REB4gDJYkH/3FGhpKcOGnHFxrXMqFv41nb93I4rTBUNDeMG9u8Fjpm
rvXz4konesub/1KHC5HfMO29JDUC18FvXLf3Zr5jcOWlSHJk+kdLaczWj9MRZz2oKWEexr94QuHX
ZI/OQK6k9e+fXA92HtAbAkZbXGysTn6wnrxUTOZKw9isHUwqEBNruOdcVp3WprPysgV29QldN2rG
BTR7U5hl2mbRtA2xHvvvVhI4QTfP9u28YGuW0Mt489/BEkFDNKffo8bsAOMRLi/hfLWAFm2XvF/N
B4+KQt3Z17j82bb9RYuisQ0tdvUuvX3YY7ipLmcgnOYZpvnEpz0XkRDBzLhe+KlbKDc2T0bWwTwW
ZLBHK9QgMlSqwsUx6mfi7G8ySuAXH1xpilJGeHDeRkjEremExfnx4yQVb2n0db1Bwtzn+fXeFUPO
E215/JBMUDxLowTNZYA/W9oyGXLVZGAKUGPhBqKxIFPaCZRnZGpjyzMUjKWB49IYbnfi74jV/0i+
t8krlLo2AD+JzFX4dVUkrq8D+5QpeQUWCWYgxW/Qn2T79SZglSKinVnqLeLzIZmVZRoS9srOiX+W
nvzMdECajJxAYbz+BSIIJtSkgD9ovNd1VyJy6MPet2JGLELSd/uBggqJ9rlTDX/Gvy3TBC8JokQk
YZX0/ypvnff6CSjBPqvk5O701I1MLRJEGu4ng0XawVN75pY0gl9MsL6AHlvwsqFEqdPPTqDVCtR5
kxHsYdDJDn/zTCNQfXM0A3ZDntTNPmAThWE0S6hTdCB1uxLZ0TwxSvxe41fmEUmhG+nhQRIIdD1j
neI+eU+kNOqupupXNSryTop+ryTMi+pbmaZop+L18p/j8UyyfGRSNztXP8A1lB9ygRxm9A7byVoP
sOOuQWz6Z+s3oRZ52f6vMdvSzxk4DkgXhAzuVTHlEF3HCMFsW3b2EHBAHfF9ZXec3YWfdacVA92y
lhJ0b76D6ua2NObeE8dtXnpwXK0WIpBhKqluXtphkuUkmz72p9nUh+P4fS+rcL7IM6hm1H36WYQw
W+1p4flYtFpDO2uDMTiaKmZgcc0a2Z1SPMPiRwGVO3+Al8Aoqkx3ldMdPf9mEGWb8kb96bupKKUe
eK7p/DRe9A1BSFzMAoUJqXkM1UP9G2uHX3OxCAypM0dnZpH+Qi6oiDYpmgJbH6OLrjM0F6pNTohE
IAFZZhPGhZTJocnG4UuOP5zx0s5kcgZfg3WO7m+NLrQx0uWUaMKUzVuIr/EgPuwaITPE+e4rhWwU
PG1/HJ3aQzL/8KX05OIaohnQiuf8BC+uQ+5ur12YhRqSHLFR8+WZqasNC/u1YUwgAI8MSQ4RxOSj
n0xIPe4fRVKViygJ4ul8I5N9SikHlUWgDUic8Bmf86pk56m2KJwG//L4t9bqS56P6ZqdZmjjrP9L
xaz8i7TQ2falnOLpqguOxWno1pqa2/JX3j8WcjlUMm+a2xGTXuD4xugh1+DE3KmBPby2x/Lkm8dO
zcdbiINoNiOo4+74mM3qAHY0Hr4QyPDOYDMAn61BQ6g+RRRktyGlyO1mkLwAy16qTthhdzYKlIyz
Sgl1UOaChvNMIJWLxVsp4sVXpL3vEvBQ6ZQRS0/jfhnyyCtmOppATbbBGAhImc+yZQSRbjUGQbXj
zWSmVg/KAVppI90EC8rjoRMSYWgTqBtY4hkzolPPNGmGtVvlh+t88oJ+3bcsfBeZrPiGBh4mZE22
JTfITfSYRTxWfpWhpN9Ukj1r4LrZisT4WlI1BRjQzja6kx2Qf7jQXbRNoa6U//ylDWnauNxH3g96
bYpIMCb7seUetDBkGwDDOPZjgjufjy+Oa+n0RA0UCTdPj0Fu/tOKu99MR9///J03vPm+vmtaapLA
wzj3g/bCKm/jUhyrGsjPzhDdMPP+LgT1daCZ/r5AZ0xFP96g25sFU00jWQRfKHvUONpOxN2A3tTu
gv2a78qja6h8rj1O7sf2vQYABQmUW/DkcFVGF/ugcnXky72pQp+meMwGsKbrMR7nxGcYJ+m+oDIL
Ben6g/mfFt9/SuunD/jmC4lX7HLxtI5M3GPKNAJO4ozAPQNaaCPSIvn4LJcTi4dg878HkAK/SKXL
8ulstKzIWeOih9+9CR9ia/vKEyFDCCmfRgxaFLrlC/eDzK0pytA0qJOAXB5z8fqOvWJvGK74Pr4l
DDzgfTVGh4XwC54bYJpt9P0Oqd2X0InNWeqMKw/aqtLCOx/vD5G7aevfLuxYJlg+xXnXZ+XE3wm2
ZQ5/08V4LNQ37jixg/dEFrbY0AueMc3N4Ytn8Vs50WonzoBnqujP+XqbHgy//DtXv6m9+YLxoTHh
7zQD8Wi+7pT+7uBa2wSFuGOcbBpnJUMh3bBgqCdaxHbCFtwC+AplFJrULWUt7nTROcR4KcbU/5Q6
tjwBIiGRZo5H3Yg6UmN1ravumRxvUcP6I+vQb2l6GL8xT03/dkDtbFeSZ+MENEQLwc5EbBXS0CPU
on/0+6jHqv7jF9+Dm4g1bgYbWrflZ8S6cd0Ad4axYKoyF9dVPdYwcB5mQkMMK9p8xhctOO0d/UFY
zry4s9xMJ5xaVHFjLLtJ9XkJ3bS18Ooobrt2gkNQRl3G24BDrms6pMnGKNqrXvhxWMRH2qy7zbyO
tNDi3flOwJSU1QNg1sPdpsKwx6n9ZKsz5wmjVQQihDEWL9HyzvGzEfJ7hrRKg0KYy13+3KrSua/t
YQaqXC5n0nQph6+ERpt2LH/ivm51TgOwBfyJLqnlJN5m4VpJ8Q7/20WOJzNGnaMVEBgezmMDy06e
zBJeNcEgDB4RqsxjnmKPq+hHDroTCNI17KK8lfD2lnxMGLGihUe0HrQcdCR3/d2hyCE6dhEuxF/D
Qp8JNmpdSN/W4Y6AHanLfYAoG9MGri6kkgAw6ihIHaxNxC1N+8AwYST9DnBYHqnw2meGptnPj7P4
k9nGPlaxRbOOiIVfi9/QEWplUAqSOMK/GADjL694ffyGIRPga8nJ8GNDkt33Naoj2L8Gxe9plRXU
HV5RJp750JzjlikFTjhQsxnHdmGPCoyHDC7QACZ3djTCxoLJJnGDUmyevcl6gU2qIOrBEV35a1NQ
Yrvj1jR35bEn8mf7quQ2R9oJ1pyCMe2ddRrF416jlfDbLvwf3Y3xFUwd0mPpMvbsewXWjyeJbiGh
hZu+ELiL+xMcOr7v/sFaAY9FelE0QkPPOri4cSJe/m3zb5zNY6fzZ5z5IZx4zPeSo93uDzK49z82
ArM0pzdq3TP6KKPx1e7l3UoqJrwUFMgJdcwFOuL81KQNG9/5PG0AnYswBaL0vXVUkAkqlg0NPyjI
uSkMMB731NFjhjr5V5a7jsR/W58swfoB402kPrhZDYShyUFhYxW6wzzuNgqToDFUFr+czg/QnpQp
dyKcc33R3W8OVbCFDHUK/FCkfNt95TEaOm3rftj6G3TOfUqeoUvjgbhNuc5s7qM6+OO3zLs506PN
qY+IbbEFe0AzcKdx/1l6AJg2jj6Qy1VQ53aHtJrxevyvjjyIxjDhS5bvPkKiA/DxfeUjuHd5ZTUi
z+TJC6A03URnoyZhWqNn8nuSIKY77UhEPBsDq+BSFYY7Q3cBxngIPlaxJIl00/txB2xrrA21whIH
cSt68Qa8RqJzdFfzTWWtVhru/4s/5rgBlJYgQKCcwUoJEX4nN6yi0yoJiOHXJhBckFBh+UL/FVSU
7ITTzXWsvzXsaYpn6rS3gJOSUVa32iKK+AsBV8Le34lY/zF3oXlWeJGIE4pe4ekpSYWx3rqTss9T
7LoCQQgXOGN2LkRMvLhi/eZGZMW+ZIjR/TkPQnn4GeAfg5z9akzqqxeKgjnpOzoP60ogNhFxmbCu
J5Un31cQL1SX4lWR3gSk/hdWl/yt76Ca677NPbpdSYLZeARFg2BW1waq9EoOaN7LxeP5I3jYBchv
c7swvt6L7WNYtz8qEKJZI6wGnw1kUvgO5dEcOFlCyiQyVQO8HA0HZNvQLAwAFMw8Rz38BdIyo7J9
lSHAcGisDV7fXR3YhCd2psQAWNhwILfY0Dp0uEl1IBkTkz2Vt4Kt4p6jXq4H9jKudJhMZ1Qz1DV7
hSkEsFKxIwE5KQa5+T9M5l5xgA+bU0TvQe+Tm+27N9fARKLwAIrJzxzAOEkziND+icv2qJC9hKQZ
9jnDR43ZWav+gqwqNCYyI6k+cl/4zm2YWEtMyUmGTbHOFCIhisUpx500RveJ4drA91TPCO74I+Fj
QdxiksyVUeOOJYKFBJ0osGmsh9T0AtQW2NABUuqhoqgEQXtBehRMaf40AS/EvfCzufSyYt/SsrPj
IKdfbqCBKIWQQPJXBNsdXHurqi2BEOXpruyjyBDfeZDBSt6wQAldA3ueQ2oDwXh+YGK4TcQVkqcA
NyM8DS5UrFNZOA+S8+rOcagezkYe0Emf2zKMzCPbMt7ntt5Zc21C8GQgp3OF4+ej435nESU6E0hR
5e1DqmkSeTQQTl58jWHwQUmfFpLGKU7UTK30ycKd7xpLtY7NxkFMkej99RYA+AIiHVp2WbnfJDCf
wTd5xLyQHfeGSgNQj3GFJWzZBrXBrBN7fWsCN74OCRI1HaRK47ShfTHqecPo5OprupXIdTq1ECJb
KgdHQDzy3ZnigCOaai2fjLVBY7WfZ51NBohiywvmWbRLnCqNGqtWDoRlWC0Q3MDOZv0OAgwYX0Co
RHCKW4Ut3Zog4BsMHM+CWCj7U9srIMpcRgy2RKmqlRU5L87mpPeJRF4SHgn6D9UZy8kzeaRnm+kv
IwhJCWYZVWweE7TdEGQrzbe7aRCxTW0Ylw1YyvfGtDtj/YKbc//HM16aSEXPGYgmjqw7Jx+1x9CD
MYUDt/VpNb5mhc/vG/gw+9KAbdiTip1sFgi5xfn5QjjdEq4NLyYJpYda50QF1VzDRqcV5RkNfcRT
5Dn/wl73SyB8Uu2Cu4RZ42FDqFzKYq0s6crW7N1uHuA4KimXUl3SPPkpWVw4hMayQf8ce9kQKa05
Oe0/7PNS//AR9RCA4wpLAKfVM9Hh40oFEWkJifjDapBcL1jhbAFCGYWK209IhIv6lr9dTxeLGWcv
2ragL2Eu1YB+pAsd5N7CMAGleLAD6TdPUj9aupn14FLx7aPiBv0/ppbzqMka8Znx9laOdTc0KCbS
aXPfc9Fuzhh1ODPRcrsKeT44qj2b4MNj8+Eeveia8sVEX66MsT8qtqHMPPwkzDUMHjMyY6G8T9Ay
oqUh4ig6ORU6hSe/QPsiPVQv9S+Z0DYhWKczzqoQ8QGmOBmcwbNazDkeVBdnxttqiImPNGI4n/gU
j1JW88MFrxjgqYFTy+7g29mNr4EncmDDyF3CkEjhmJPJjZgv/2jiHtOGU0Fq+CGWGGJrAyERihcm
uzVzGAkWx83d2OgwrzoqoFUOlgSoppNdXHdrYmZ5yvxRDbMULfCIsejWit9jLa3tW+yFq3rJbFuR
OcUWi2aN8oQi4F/zxNKHdmcJXdYZMc9tHTa1QIKPwD2YpyfskoK9fLNeQaaGtpQKhyeFahVVMtU9
k79cYqPYS0unXbYxU3oxiSl37520lBEPDGY31N7GqJr9KphlibzC6niiaujtRztCqGMBsDc/Fr6o
SHUtFjn3TdBxi1vL/0XE4rVfdo9LK1dwC+zJBHBQxGX6ipv50DokdixKmkAELzam1gCQZyA1oVUN
L5LdHpTkEX2wbLUIJyz/SvbiMpIvqOuiPo2XymC1fKvAWmKUt7xLnf+tavv1oKIH+GKXUTdfirD1
CX1/Il6J9RxYNVOFP0P8BJrgO2DIMIX6ckNgw02TEIFAjd7zpZ1citrJEdPmXBSFj+DaVc9UNREX
LZZPD2cg9UGYMgSfGYT4N0JrskM6A+x92CyDCzcdC+yEfEJVX8banz0FeHwy3/22LHOprmH2grsF
RGccoVJnv9MG2+JM+qQY6Ca/4WJs+cbyw05ZY8yJth03zhv9geCB/JjiU/44FwXnZ1GebGluWgdQ
MU+bFIn8auenFQr3mk568JBMdNw4zBy7eQ/pPFcB05pzRD2O4jKiF7c/TjcvI/WTXl4nIhojQFyy
mbRqDTeq5PcP6wKHM2tQLI6HQ5JJw+H6DwbIujeDwsvnWgw09c6in1RaU6IKpt1LllAWkq6/Pwaj
rAtKEBq1nA1jBEjDUBLnI46HZ6kCg+9/WY0gdzfETSV8RN+oOKxGotwjS6cgcahIjQ3dS3n5T+xq
FbI/DBgmgLfrL2J7rxLCZUW2nm5/lPYaHKIttp61/r1uJbvUWMAJomKEo6nOvtoJ4wMwj4u9RXit
R5Iwyu9qkGwwvEsw8pWbHS9BlRmKRTgtFFi7rDMlaPB60S2JmgPr/FMMSg5jzDmA/r4q4DorkyoS
xr0yxSW7ZiAoCF32rr05ikhhB6j0Z/9oEAMygNKTp1ZX1FkECVIT5RPuPYWwp0T0FIXtfVlg13p8
IEgS+pO/gzy/VCJM3R6J2JomyCG6Ol4cNvE5oWynf4k3Z9MN1jAIFed0Sx5+ORyw/SK3ZLaAeATL
V+lDK4dGaYOPquEe4vhcw+x9ibFiDk9vhEUys/fnUYXGljX2mNL7vTCGeEAzQYTy7FGH/M1lOYoE
MTn9P8KJpIJSd7bOCs8XCeR+D8Bz/dh7mXNZ4ojg27Q3OZlAK3thX8oMM8wMFfIfvNpINWwvqH85
GYskCTYUNT79B+LF2Xt43Ql9sAJKsROybyFFWtUrt8W3zhMwJ4D2zS/t7zd8/h/kcBhA12ShDpuO
1WM4pn1eDKbwsUQocI22qx/+cGXS75o5c3/Gyy4vIfUdTvRiZiznUQ+jbDUoM7YycAvOVGmPCAv+
8zu8/6s2TLZVvjQ+On7IYlsIJVaH/8TEFMpx6gy0NyVa9gkGLhBLN8FjwDq2XJfTmGBuuQz03ss3
54SKfF4ACPDik5p3oMmmNqzr8odFBp20z6sT7loQVyxNBeRV+8CXXAOYSnTr4ItW0RDBwf0sbMlt
Lj12cUbkaNNt2emYwzSu0hWlonKYTS2Pgt3YfuYCTqquNiNaS8ARyMRgFNGbNTY/JpVFw+I/aTkW
uxGcuLxeAZg3TrWBng+MCwRPTKOVbOrPlwt9Zpg39iuuD6tYCYDDvaFoH5vfSYfHcg5/etsAMiuk
qAzxr4/QslfLIPlZ22rvFmJyY0Mhlhbl6suNBVFfsC1wQPZArV+8pynH/gATAaLiDWfTOKk95iuc
P0H9YdLYpJAJlH3mrmikYEZnix3NGXLXscOYp4PcRCU+KagZQucxr6Vj3qPqw4mfkxOUIRAQgM+h
1aqWYG4gAYYNToxorDmTSf/FaZycP1JBDf8jTwpFB0LIP1eIGJ7rAEcXraz5e9GQfKNi1Nzfvv0x
Ut5qtzE/c3mDjJgwZ2lc98M8TI+9MPX9odwkqGUkda7ZQUz0gOz86G5Ph9b5tmZIK2xOMKTc/8ge
F+k7651kePZrJaY8JJr7CyVaPJ9IRB1/GKlXgq6orGi9cG/jb1zJ9jDna5bWiH0LEqFMS7+WguHo
9GEoc7iKBkz/aG95PjIBGPV8jG1dUbFEn3uhWHzfqMFrz7DxBMEmk2b8lT/yTs+xqW3qyUPlyQb3
5Vw7czfOtS7aXyyEo7HXdjsZq0mqTNz1XuwFLdz5BM2ZYa/eyj6a4j7BVB3D6HT1Q4fjPkjgMcDY
WZROKxGH0r0uo1irZx6z7ia8kHCYMNuqZf1Tp7bcMX5iCG0W0vpaufbmXOBkJCmw9TrBr8AzO1FQ
PJXn/rOog6jfhYap5cUHd9M3jVy2E0maOCh8YGGQLCxn8CMn/XEgPpZKL/J5nXvJCGNP9Flrdv5j
hXAa7ahkLzQLQAJaPR8bsXf9M5YVBDKzOTLhHhhXAO97JSrZVh1ENYeQOz1FxXbyelbB4wxM3gYK
hQTFjKd2Ov34O1HVYrSlc2Y7g7WOQ8Olk00Lmqt7NIAXUUTxs/S++NtjN0/XvKVEZiuFUsRxgeQQ
W2pQRSJzvgUKH2HdT9Hon0MNIFOEimsa7mbdwXDOkLgkeaWBqtvJV7hFul9NJ1/lSUWPvy950NrC
zLF5Fk10+DS4lMwJHKq34ASAw4fFVE8XuzAc44AvwK0DvjuC9R3haL3kkcFHmMgdoJD+q5386/Nr
b1ojSFu8jTB/fdGM2Ic4a8I0xGeT3JuqbIV6ZuxFREmypMo6YVYxWEf7PgnIVLd4/aVylowvsT9O
0x08aDcj1Y8XhkxxwCzz47tIaZXqDMa4/uV1bDEoQkYIyIx9MuYNpej4L2ZPyiNtLmuWE5KgoFdT
a2paWEDMQX+/AoxF/pzd0oogSGZjVlAH1+XZ4+DfrprfqCu8syn14k4lSacK0GrOrQaqbHd3y4b5
xab9N1Drwfx+lkVWzIKAgvRydRcy/TAM4N+sIw70R+eJVH13Wva/vlmWoD0iw6nqQ9KY8zA2Zgqm
kv5TeSQeteWV1cC8Eqt2OHuj8td1w2P5jrRs0hUIf/qH0b4ibt1Spe2qatvCpChMYvVm7oAGO71k
JpiccnvC5BHhCsy33yJD+uqeQny15XIU1EsiqfZtFOSYQsraoyIlWGbfj/YmCgakolm9aMpnDbA0
owPJxU/vFKtxC3Q0H23UABdcgdgRGZHLm4piG1Z2IQ7YvMKjro0dtb3P0hxUjbmkT3CnYzpMUi95
wggVixaeVNEIsCAD6gsa+2GODwQbpvyOq6+8LFysYvScePUhByfMrXI9imClCzaxqFgz1RqT5Ahz
E+KtnIJsiThQ0wBrcMD25NpITVB55A/5geEtXeR+H5k3pnwaBtJCFsrkIuyepi6xVlRKLAW654u2
HBDLNKaS1EmKJFZamlNeqmAMjY0tPG8HbInp0bXnXRyZ0uW5OncSIf3qJ3e/v9mGEkN7gqzupYCh
IEy3g+/2T/AjwyQHKAPJ1SIw/wKrfRrl8SfHwuf+1KlyBaoyzfLzT4rAfmP7KJIdhQ5xGXJx7jy+
v4yK7UkTh9434wOq24PFmYfrQEGBjID1uSMQA9s5+ynPT+XWci71NVHgHXBQ7xLByqY5DCNuzor5
13eNLUxv71XYs60c89yWITou6FEI/Aql4I/X1ZBJy6UQPNN7STv/DGcJetnFLyO/xFI44z9ux8gU
8lOC1fQXF5E6VbEiJeR6E81WgFo/fCRCEasAeejTpgq+gpKHpv27QwerR0c/cygonimCpjFLf6IR
Gucscpz1PoxW6HpvlJ/fkz6TZ362gdr2oh/jJcmc+EIQ6hDKS5xPsib0gGA938GKGiCeh6ScZiDu
2c/f98mGUc2lxOYQE8rc9Yh2Qab7ah+3uvFlCoAaVEbc8uC8FrZnHL5vG2LG+sQ39SkBjaNltdSk
tMlvfm6HdWAu/F9lyVdD3Rc+i7+1snRmbBuXIHC2qaxs3+U9LYvyoXlfh34Nl/B2CWgeZsf8s6Zc
a/Wsse8IFzVfAS35ptXwQW29Wo80kF8zQ4x2baUE8pQ4eHCrqN3Mc7GpID9tY/xNa/UraSD7MpkU
htZrIhCS1ZGMa2UfD5dD6da2ry6zLXdW9tFx91jvGXTpZWVqkK9RGCELM+AZRP7cHgpeootox03F
TcXpJhV9PbJViZFOk03yMF0Ogy4iCQJfB63f8RqI+kNpHCDhGrOobLvSK7nqOL3thV0pNEjazVIp
Fj78G7yGIftOUh+eLwloq2xq5O35YO0At3SsLijdW2fPE2dMRAiKWVySiFfneGwn8mVe20ryoqHO
Nf0MVZMXMy7LAGs256InFU9AYZ+JaLTBo6Kw4Ib+flMoaFZj4ATjy1WJ6NnTH6BeULYIOWeBtJmr
Io8D2Xo7XdxH3ELd2SKs3BSiOK+CCdpyPW6UWe+YE1acqzETA9hcwMvlfTKCWcYZbhb+V/uMZ413
3LjgL07hKxFfa5Y2g2xSFT2w0GW96yrvqnnHljOCLp4Vuox2I08KJ/DhoQcCmzjkG5YtBzxnq+0J
SmHJ8gEv4wEN3ZKIN/op43v8RmsdlHF/hNPtiNQ6DyjTvXK6v0lPfuVmCB+52bM4znUIv89eBJGc
FWuAhz9Laq0BVlByOp5xZCg+v0vbk2rmtrv+CNkQZoAOyhlDkvGou/SNvBqvn+AQHZgC/pBoijlk
2yTlIRnSwcoSCZG1mepSVyAYy7rzVGFCeVBt43bSMyH1elIXIL/O8qw9TWxAcsFZEQfHVpX3KQOT
36TzDqY5Efk+lJORdfbb0fWncq+cpJqVPNpGWprttqP8Z17wmEsV9PtqCI8I5TjL5U/05RBZAa2y
NHZxqPpOpIwLJ7i5LLFNd7TpaGmnzL5G9Wk+ETEMosR4RLDnVQHLPbJ/knINoubvuoFtkJGuMDFb
tuzVLFGagaqumMwnWY1YF78L0f5/tO0WtgBFWkx9juc67lAluxDJji+rosZ2zMzjzWGOXcVI7C6T
GAaPP3RiAqlr7IhndQHs5rkVVrKljnxln9+ecMSeUuJ3i+qMH8o0S14r36guSmrX3cFd7ik//GU/
9T/6rl6+9+oBr5zG47Pxt1P8mj7Cj9Tox93fuQ/ELwkujWuM7cFK+0Plv5JqY2AyisvajjlFSDoo
l4RoCsRHdRw2W0k+Y4RQc4Mjam6mCModTLPoz147AxrYkd3hoTYf8D6QvTj9MPMyDMo2b3LIW+25
Bh9tcD5FcdaSEW1iHFXWbC/YxeXhgacw6cevPiJJNEdBA4S+JeTF1qmsRVeKr6nLFGsbjul4fZBd
jLMAL/xBZzC2rKpsCPLZDVA3i1ca/fd2MTUjkwgnNHQLwSbhb9TSUg/LzaWGfpacDnsL0zFZkWDm
YBJP2o+uM2n8kyMBMMrM39kZJ5/tdXNiT6Drj68v/i3V3CZDJ+rTbwyN+vL5qh20VAalw2XwMJyD
59b/6olPKPg94TE1oZLdFcrK5JylOlIdoIttK3q8ZNxCz1pEJQKdDpeIpe1iHixPzF22noPhxPys
DCQiA3l+WNwHSiKX2zRYccQ9ZY1dUnDrV7d16SlP5DtZhaBbh0ZpNZBnmGvEC1iidGqHEYdnt9xl
x2xOgg9qNERQMQxeiKiNqwLY4MKxNqayAhZ2r9jh7hHrXXRqlpmVrk8hVg5zuoQsRXl+BMFjHsrP
IdmIpnHTWwxbECQ7Iafk4NiaOQhTKI1i541k35IfMBAfGw5hTPT5xgbZu7zX98kr9MWVkQ4qmgP0
1fjyGYL2Tw6NxIWSZq/Wpq54dhTzSTQRPuo4uPdEtghoOksuixzmtq4AQZPmOmfh0G/IHlSVsssM
Q+eJ3KSvKZPSuDYDoiLbz+YLYBC6E12iLhOxJ0q9sk7MwSC6IvAi9UZRpOb9naP5U1JOnJ9puqVn
wOzYkWnSNX8PHaaUaR4h1BHfXXeJEx2yADDVw8geMY4ubkdlPW5axKEfUr+EmNZCd1FKiPub+kg7
7v/fiAGmokfQHjSr1fxkeCIDLTvZZUMl+KGYWnEdnjpMM2freb+05LbIdguTcuwu3hpYThzg7W0Q
bsYUHuVVvwLDxZhUUBefSUVfC01QJNo3dmmstfFhKpQwSPPdmtN88sWraOqKOuWAAZSqlVjEUdcC
LumoFjnBEQFfe64egeD98VgXOTr8EhB++h9fDdv452WUn1w9Y0zi2ls6ZJWwOtFYe9bm769el+/V
zUd7iZqrlQt3WVVx2k+tJIAfCgoc4v2+MUs0sq+RsgaOGAW670Zuk3KJYLwsZHaIJQWh1R3pwcER
w8cUdsQGlkaK6dkxdYjIWtjiGfm1kChBK4KHAXISJzl+T57PvaZYGXLjENGkML6zf/VDMST++3O0
R+IxcnMET33zdWgoUoKovE3OOOld/eERFkHGgkaVQPEtnQ4bu2qEbi+/LRgbFSK1aGAGmpGHjKuv
tSWYJIDsAZMN2JgdcNB/qG+aPn7woEqEhLQ1JhOs93yIQ1dNRKbjn0uocxq7A/GhqI3kLHvhdJ0D
8FMUQ8ta1NipapWo8cNA19zyPn6UhwnfKSnC/kiUN7JMUWJnF6Xz3JOAQBlTncLsgoHtoVk5XDnj
bPb/TJO+IaKCwBsbHGSZBNy5Q67W3quRnR6XLs8WksSOSweQUpZ1naJrPNa/aSheafLCfPeN3B9q
zgfVXt6iTSiU0GconhT43FkWkRsrREJODtvGKOEqYwlZi5+vMT3SZ7freBBgXVSLQRn8St4W9o+p
wwJknD2dsE/N+DZGo0yLkgMxB3Ms7x83whtxC7cJuNy6NwS94jvs9VptMkgJb+5+fPS9L448RShq
ADJipi+fwi2ow/j3s9NYkuZA3J3ujLRgYtKszCfmaa3sI8K9tz/Odzf5ThhyKDX2gNOIFnaEy/Rm
rBaiGXRp0qOdnpHHaCw9gBHlCbKgjRk8Gir3ccJg3OvILeE6PxYaGcJXOP4Ioku2QZGf4ujeq33+
PVMKa325DaxyjbnrCjA02h3xv68hXg+uVKdaH4aY3jt8vT6YCqvHhgbblT7wHuGPxnbENRVJPTkM
HacWiSOISsXXkpXANu7RLIHX60IM38Fi30/VKhIPApz+6JGc1RDtHMgF+SQU24+2CcDMn1jk6bOK
OuHpJx/vlCoSIf00O5QmXs4fy1715Y2V7QfBfvK5YHi6WjqL2DZPDF1uB5lFnA9/0dM/qM9yHxmp
ADd30io6mOVjahaDrcIMGh+Q2D7EhQbO65oC7r1QDwQyHsXp8Dhsb0P0xmHpNagKu4nuvsyevXa/
VSWMFU1cE19foGYnsdspTmIZHT0xhDVeUyYTgPZi6hNQiCV+JBq2RkJdg3faA5bXDAO5IoujUnl+
iV3jUc1Fjg+DE5JDFwbWEnJHzc62u95wSCYPuu2rYQAy+ystC2lSdRiz5PJi2xfYfMLsgxaNKf4/
CnjJ3fG4kjkdmPW5DhxyByqtq1p3W5x1jqO68/XyuwfOyborW4M9hdHWRA982RRYYgzTeaGRmvrw
I4eqDyLdLrOerMUh1Cp/ujQd+J9tV3dhOU9Yyvgrq7M06k61XbeFiklrYJw4LJU8fnzfJShIyK1j
EVwgEuXMsXr3aZqwqZ/6Be7AZKvHif+deBktBRv6+3NNO/9Po2of3blgfBs9NHDUjgxOsMbfZqQp
gTBpUZWNw2oRTlSj7lN1zzPM0KNCWYXMMOMcM/zYhDox+4v115p3L7pNTJiLXLMvpQbt+WbJTCIv
LHjK27rRR45M/JApWwqjk5ZF425AEiCURr4J4jVCaL3ThA8fIBrWnvr6eF2QHP7T5+loSluD7Xle
/CY+J4dh2hcYsBXoGg2vtY5Qq2O1K9TkOvqg/hRLJIVdRNlgI09dodkKPTqT//CCTt+9+9MzGH04
PxUpghNYwX1ijm65AiJWnfSCU3yulO5NmDyVEomomDJXsrSTIPYenxa4RAzhp8EoqO/7bqvR7Mrk
cJCiA/EzpbmhtXrrbek8lrym2wl/tQSDpyNeWdNJZ2QsCsDmAb+EFoG58K6i1ptl162ZNBuXhfWK
RZp4er/Nb+f0WpwaRCdiLwJ5C5xTxcTpG4yYZa65tyvY84UKorEUzT7s7iARHZ7vUYQbdNqoXIrZ
PCJ/UNmoYvbAJQQyJs/df/qMMpVy3bR0rq6TvdxsepNuwuQMd3z486PxGld/zrbyqkX5HEMgeHIb
mW/dvjHJFhoKZ74OADYekBuQfrPrlM+kZEJQQJBK5tCtvHnMEA6jyp+/ApC1X4TFOUhdIRuLgFty
l5D/okG046BK7vhLE7nMvJK+HF5KzF1otDqqnRrM0qnPW1AFVLxxzLzimb5TZPVzcYgUA22aQ8S4
LThDif8chzB+qscGpAkUiGvnpBkaeBgzE9JgbTZxek4Q5czWwCgWoBW1N239HbZHIxwegvYhTsH7
r7HeoKamVv1L+c9JdC7bM3XdMIkF7dcFZiwzzE4RIM6YOCiL/Xn2KMMaM5GCSwwt6m+wb643OBdD
eNXzVEHoMOgCz2JYIQP9ZEqadSGxzSw2cU7zC+Ljc+IcJTOA+RKKdaac83qkBmbcUiL9dUnpNz/Y
j/u4rpG+R+DA8G34fDxASvK+0IVv/7tMOlCX9SrGImm1AlbeoTXVaMn1Z70xizEvj3/01mz9zHU7
DeoMBZiMmUp1QTdCh0b8bXQg7Bkj+HWiMtcbgA0CQpnRN7YAMOf9fDg1f1/r859AJKAK71H1XgYH
q+TJpgw1r9M1ecQWQEpkJwe23IFdjNyZNXCCX63zi4GCgvy53tbMARm8CLkCB008nZUEJdveweCW
jkryXMRIR55uBKzCUhwz3c0KF1xSbjv8mhuGG3WUngxwOV+lDp76sMyhYC72pbgObpNB9DvA1bVy
NC2qsMDVIfMah4AYlPSJ6yRpzKfxAt7nZ0pJ1hzIRl4N8WUDkVRGBDtWiNXWJllT0qfsbmE3OfAH
DuJZo1vYKaqia+2j+lmhgznCm87SWEEHEs6Pwv10lesWwQR8qEH90qy88WalGhaKOBu+U6crhK6l
EfI7ylp3IwFTDbpDCEPU4QcHk/BY07AImKkbjVM+TK8VAvQ8b6sMt7Y7BxPhXUjsG3HGGvJPU/1o
XEvY6lxjZQ2P3UvfAvbSyWBdYYePb8xHj4k6vyLJ9pgwRiqLYomWfNTDedSkne03+1VenK/ayS6u
nbtC0NZpaB30lemPeXq9/jXCb2aHP6n7VWgisi97mvZZGQDyswObwHxICYGa9ZTt4nwf+OBVD5w2
cj1er8Qf4nuokBmKoD2p/q5PWER8r4sAjxYE00ny4ZGnQQWclmokSSDgKQ8+jvryHgM8IrsNhA6z
fYmZbJJ8HI4GMQ9LeA8P2Fcg5c145/WePRol90G8YrKMAyRfu677Ca6Rkmc655BwupW6L2HucbQn
Y/3ME7S8Bmh4a8NEyDPd0NeOF6Sx6F3ETyTktrz09lNzsj7w+9aMUpLkwYO6tMSeCgBfUDVqB86Y
m+n/Rbqgg11soTbJ2ZI8SpL3WHUxTd7tcKcYumyLHtAaLqhHS7ldctHZiV/SGUfY3aOhOlTVgC+s
mO7Qto4O3sFQwptcJPwYrGylp+SmwPRdf1TuBKopt1dOlO5YIYcW3BOHOTWOH+pnlkj9lSw3oOFi
qCs2VTBKpBNJhik2KNn+9DbM8SApuEMqApJlN2CvRWWUzkNsGGXejznGIBV0aGquxISxGGdts3A1
ohdLFhwG8tgpkicZ4O6epy45iQfu5/J0IG0WdSY8ZslQSP/TtmfiaMkdtF32oyuLDqrwY/0fQegZ
pooS0mqnseUUhY/pX7QODYaHPY62D5BxD9Lxa/Dc4dweLLZJfI/Hwl56yIV9brjAPWBAlvVhfZ9R
qtWxCh8I+ixA+woAbaBV4AkJigyDotnB/U7imJBqdjpS/p95NR87V9cav0LKe1JiVbW6XkzhfYpy
Eeuq2nszmmb8r9vlgcvw1c0iQ4Ok1FAN3A0+rK6bOWUrB1AtBqDGIkCqB50ZiBOtb7EntyfCDm9F
z2uPZwE32oiI6x04naHEvdD2TdXPlQmG1JMvjzaJ+snZZVXOoCuh6sNALroC/Fe/Aae2fZJVQ7lR
piTBMIuiJm2muL4i9tl0WsyKr6V4rkb7Vl7tkA8Ye2LLCGaN7Ww1VB0dehfTpHLQan5gDRNP34IA
qvZVVBIz+mdeCx0oZzSnNg6VHXbH/d4nQFLLjojENdsIszPpthVFZulKoK+ps22nhndYmg2sjk9Z
JqTFVa75g362hZXlL+HWuWbMm/qDNqQoimNNA6ZBs43lwFxgZ+dhP7YdBXxz8dsnxlwk4d11eXg2
owHEsvsy3d2H40wEh8Z6JPSBQrlHAwHLseeC1Te/1NZ+mpHEzv3aH4zWrD9nZkdc8YVGT8vo1sx6
tYh7rya7GJDcrZnN81n7zzrk9S3du2ypqtLw9C1cDgoaGDBy4EP0hmLnweODn/H+E5mEZ32bdy4l
m3bzWbDPIbqQba3J6EVr9T6dVR8a0lBevYRNDzzlQVgncV6Lc1h0N7IJb2iS3yg3Xypz+YTz+bss
5Y4mS9r2cXoxjdeSL7VDThgVHWanJQjf9G+u/uoGNOa2wwAY46iXFPzxbPcU6R7+WoB11A+1KeX+
W04La05RyZV349LIxrSE8/cfe1Csf1QTk3g77c5T0/4n5JVYVFT8LcBl/tGBiavpE74RTOSeHnZy
+XaESVSwgVfIpU5kvd/A4WwX/GeAqacfHiEl6mDzrz7pIoY0iK/NH79bDdSFBqCkywkE10/Q4ZWu
ihlATOuLLm+GR1uing3xD8jL3teB0uNTE/PUA10kw0luv6WzEJhvPIJcYlVp5KbfavYCWjuvOdRz
LDXZqHNGLVppRzdnpu8ZztyQbJWuxypyxAVgg6UGNIAp13rGYLsNsWMXyZritnLkxV4TLqEQEyvz
+Io+lDjNujoK/DZyoGW3m0TTxY7Wm9SquZFX4b6eQ7vAGCZoGGEr4xg3V/E1alUeqy2edaFgmqHw
CWJ2k2gW/T47RY9U4nsod36SMRWCA1R6DgkYXO41ntZ2unBUlHKFNOxQbgFWOSZyI7AOUcp2c5DW
uQgS4SJ0EHTpgy0gpJiCRvceQOkV8/JKr2rSpawLZ7fdNgQWI0XvN/UynCG4HwHWUPf5jKY8Vudd
LJqbkOHxTWBcLxwn84YJfOKpg/eUMja7sRrPo13N8W2Hm638/nYMzcmKqy2WckXkg/p1RwoTQ8of
snuc8hcAXucUYIs+X/hNr2P8scXpfkRTaZQoPjM50LtVfaD1A6TP+AnIGZaOl/2Lpx5YDX1KZbB6
+8zBvz8LUBGYE9+Yw36nxloSSuGPqv6RkYJ2AgMbKvCoPyeW+dnJfvuuWpUWsBfKYdU8oR/wATCx
vE5RNAhxvqZsi4vV9bQm+3oUjxf2wF+ho/hg4cRHqDpam1YeV3vkPESye+b/tiPfXT5+8J57dPoK
iEpo3o67OVGrZmN7Jn1ozbvX64ElAwnHhS5kh0B8egsicZ7OQO5g42L9udP7Gokx8OHv00u6X/bW
fpklTdtb6gwMwH0v1epyA08BWeJIh0QPHqKGW52IyFCM+tEpW7Xi+eYmK3S6o4eHIeiPrlTsc2HM
8Hl5X6dMB8Y3q7pMctW5fypTwAmg+NxmieldXI3RlEweWZvrscIf/icNXmN4a1bfyOVipWf0VTAy
U0uIjaIw9bNOy6v3jVzGjMsCBe1ynwgONTbkI10RtaiJ77P6147GnN5bi686bTc2OgUL2cQmc8AM
64w/R/uNOcFhv+44RlGGxINVu4GKUiP4oGUTJ5Y5+tyC6mSki/nn+DbKzOZTZEL3e7Q+grxTpwPi
/4R+jvFH1dzQ7f5Zb8IPeyDxd/tb8PiKsH+/A9wjXHJC0BjBFYCFC4L79DPBd8ou9byn6w7tejvL
+7QB6w5G9YUSzyBi6vxd3qGJOeAcIrKgv7hL9z3lWS4IE/yiXXHW3lbp9sxrqE1rRviDCl8gkhMr
uj9MOLikuEBFAOQtriIXlYQ81oV6AsADXRaagI+RlzfZJqZrVDNpvjQjg8qvc8EJbO8FjfycMU9R
c2S77vw12Fp4/eu/FDkQaFQLmYrh+1XuvUfYLIVMtCs4fBGMWAUaHbz7Erq1LC1Bxn7Njxvd6T03
n1KatuXdHQdSnQIpvqYgYaZCNjy1LSKBv9Z16Y66zm532+EhAuUH6FpLQ/2w4tdWYQAP02DGMj4w
ykjlNMJZh38Z2Rr16XeNAQe45ICY8InSqskvWOaiIRdURKwuXZh1K06boFQA1Wsb9LGgRJSsRVEM
sMXkevQBDsGtC6vhFYX8CGuyPKVY0vdmNd8ock2aTkh41v7eCb0VUCFCnWN5MWLocpmRG3DMAU2m
fe0Px4BB0aLDTLz2PUIVXuwuWKCSz7IQXbu9WO+D6+ZSJjbalUhUV4e+cnuOlJLCbpgEHUBd26gy
aUh51uNFk+rLoPkaf12Zy+o9iRsT0j/tlBymFrHTazfCeEozEhFs141K5N7MZ3+Z1IcdKjKIdzU8
e1uDHwSoxb2PD2YzMD/6RQnOiuqkXI738dJ51n3vLs04cAgEBVBXSrnE5YfYP9YTN/SCxuE3XcHN
lT+7T88RPpYT+WvbX/t4v7ukHYZZ17W1VnTPlsg2TmPiWkBaDzZvLJZV5vrQosaNqlWsYadgCcqz
dEp+RELmfWHL1Anicav1uW/2tzQTyptANXvW7ShLy5CLdlcl771WaR0U4/q6Jhk3pb0gzA0RGZzX
4omI5wIxPspSurgIJI8Q17aZ3JtBpOItq2Ad+6iQN61/pUJjyM2D8i37kNK+ilcTatv17o7cH1sA
LuhB/miGhpieMELDhUvSvE4qieBNuBKMEmeRh1Of5XrAqhPt+5XqeiHSab/TFrTLt9g827YPAotH
8eKJDLxji6EhTMZS3/65amwRMgYb2BTT8aJW29uX9K40f3sZAEXc9ieP+inRKEObx+KkGEV70lVg
mjGqy5j6yk2/1+EFCjWWbSzCNjV3qMZ+DaLYV717ASEgpkRaqgrjoBJuPTsDjZbhcDmPWYApfK7g
7qMo0uKzDPDIPsxbxru2k7Xs5uhPNUc/TDPKpB7zBThQpI0rIuOGwOwcpoEi8u3mxj8vSUPNpUCo
dlPTCDjMYVAM/MGRT6Ba87ADbln1pEixklYRXe8qKOJdhuqLAPg1vG+GDhNKpAfzOlnYIdZas1Ix
owG8l88udV4XBJtyMCvkdRF8Kdl1cTowe0+qGpqJjEuj4ek3Pk8p5tjpNzZ94jlgCfyI41qo8FK3
8ry6qb+cAHZFSHms8y5iXXgD6z/M9FWiU4d5tOW49Q8f2gfvl5HkSuvM3R8yTe0k3x0t+xhbvoSn
KPOL4TfK1QYggbBiftsw3MVC3yvHUiwDKmmS5Tutm+hNzeTOAoBhhstkjNFoCh6HQKzUKiMivc3i
9tmF351HCQHDkIKRkblYhzj+CQX4w6bSVCSsLjr6TLxh9tf5kW8UYPZZhuu3gERSbEZta7JwO8GP
k8lkJhucN+J4RH6cXaA1AnXVK5vJu12imhfIT9F2CgfTzj5I/b8HoENoABtGKDktqWLzDLMTIMSg
gT/uZQp5OjWKWplmW5evt6HkUg95meTKL9Z2eLrDpYpLeEc/76XS2ZbKKUBsxo50e7D1H/uqYnu4
93As/wF2pDAR1Rp4gkGUJ0Zg5/5UmlKLnQ3OYiWYYCyBJTVGxtzkZtnQ8Yyu/QPR8z+p6NEtNFfw
TL1/ggrE9theWW8VM2pOsqKEijWsnJTm79nGVHdAbycaa8VFL1Yji8YEnKaNTBxzcphpuNYwx8Bx
GDEl1QQhGXMonjtGUKTN1NOp3jLN5NjXhu809ihQWGYyORmTC1UOjfabNT3TvW1GLWwTQyz8syRl
Z9is0aWBhOq3BOJ93K67tpol7FLbNwO5jCtKm859ZTKc2M9MR1c2gnIjDTwk4Z9k34A3iK07rmQ/
T/3XQhAWmygYNGnqfb4MOPt0U1olDBnyE0pnLpD6IMNjzJFmnX+4zclcE9aA/qrqP9Zodh7wfrDP
8MjrLUyvT4ZOhIbdnAifApQzjxLjbTlEvmTzAaYbxbtd8ycPlrXxYlJBLAjdkhe6AitQaiwsV0le
xXdcNQDn+tQdR+i+NGaxWTlg+pH7HRKvJTP5nIaIQrSAaapYKFoy7yg8r2ekeL7eUSKjkljIIZ/Y
po16mhu2NG1WCzICTXHUWCx24HRq9VePRj5yzRVbDDSjZ5X3PJFP4/CxMLQZXULmX/brepGh5zET
OQB3Mg+zes1o1uNi9akFT8MmXn+QdgZWnnTqEKDc4gXaNwM4+x+I5NguEI3XKy+M/DGNbT6Q7+oh
2Tv/b9n/ZPFP8e/SASuKfHKyWxeHV4ekLRQLYzUr0VeW3TQ78PV5CFx/L7fsdNhTlkfCDup5tt4s
7Jl98qbiYnDYzHtWoaAE7U90QrnxGX6p2ClZ//rrJ8xwaQmnUsTYlq6CNP1LLjgu4KU6RYTwBGco
qjq2wJTQ1766hc9QYhAXpLIVWBvEjh97A+S7eldRubwN0MGwhrwUQCiQ/9oGir9B/XICn/UTF2aM
D8JZByxqUDPMjLvtVNcH0tKh4HxjPs5dYJWcjdEScQvcvvLOXpz9szUIPtoPBZItMRNqj+S30X3Y
lNUYr+OUHbfrwvzfDaWVqarZokt+xgp6RY3ZAzz7vjMGeWLS8Pr5ZMU41o2yT9s/Ed2ACtyh1SzS
a0jsfZD8v/RkTWTrCPCYP5LK9pLUlAkurSlSucS4M4b9jcVjrn4KX4qUt+qpiHt47uoSHu88OXNx
16h5OrrQHsinpGgVITWFQoIC8b14finKRzPLMbsjuWmDREc/hi/9R/QwImuV5fJAHhdMqZDMKaw+
x/zTV/csotca9knbUR6WvA9pL7xb5tDm8zYBixUB9zbFV1n7atR28kQ7sLc35yyD4F19EtuT0NiY
c3vRM411URIx8b/Qo2lNU/xu0xfDxVq7MNQzuKVrWj7E5rB3icyjvx82oJQdMeQulV52TqcAyesT
55x/R3Etu6h+sTOAlQpd12ihlxJXfQOkU7DF35cP3+OMHamvK6PF+8y5X2Bb7RJysg5jIda6TzdH
V08DUUIOeQeA0y9NdZHFObjFMPC6dJrS2kioZLFRl0NQB/TaYuznF7Bfo9Tkq5vJJpFmLhC4endv
5o65mii8ym4FQjgO291JrJo3x3rkoKks0T1ixE5d0kH9ydAET4fSlQAU+LDeKwRT2DQX9cTnyu/p
2ZVNAOP/9UQLxUTrNDzfb8OUtmQcWPl/32W1MOBa2785SJboC3rDfBwPokP9trLqdlheOH5+N6Qg
V1ILdFHI8GoeFT+3LkUEgK5HxKS1HU0Jb1aZO1c3JvCdugGwx3xwlfgyUcqSDHHQGa3402DDjktg
0hAXAq7rHMvVZprKm+FjR/1dBYUIn+sZRgOmasnGj3Fw+kanuPp42CH52EeWAswFStHrqxc7hLs3
CdCNGhZazNH5lou5jlXqSbVaOQNKl4bk+9/h/5zzaQyXHJBgsixJi1vFKM7l3Wpp9n0w9pO8N2P/
enEnDpzRAjhg1qNrmeL6VtV8uFS8pJoPHq3UknTIWjj4o5Vrn3jgkHtr9QCWvl9fnd2RM7B11dvu
qreJzbsPMD32XUX9tiD+GbAr1Bs1N2Jq6JQlXEyrCo1xsRvOZHyML0Q2L5USsKP7Cds8MKeKWcIu
EbuDLzllspoe2iw5f+Q9QbCufTFHDkPoEo14panJnAsHVfaZx0wy4S75/sR8BWaiIjTjxll+eDS/
QsbzRix34rBpOoa8X/i3Ev11hWofK7QRy6HH0J5mApytxlOufc2CWPch8ydUEV2MRbyTjsXBVnxX
T3PF+bdEkNBdCyBpLSSYoEK0xJZ5T/UpffY0q2re5sCVyhoU5mDw88hu+3A2rSfH4yZpwQtWE1lX
a9MFPi+Qiox8glqzmayv0Yw2/aQZLcwhjrH2T8w4DlS4FCOANfTSPHJ8Zi5xIIe2u2CtYglC+XXh
2CO+GP3RI9jaOCVs7Hgy5SMm7ZWUmns9UOQIzfXy9/oCdYdbrWsGc1uwwd0PgXtUmWzsaxA4wQsk
VoHdLFAqBus9dtRA3RDRBKiBykUAPoXyGF49iGdphEU1JXDXDZGBisVMORoHZQGPiHAFViVmDtdz
HH6S9h7JeHKc9NQwsFbPA9x0peGBTErXPHfd1GH6YJhxkczzRWfzHpMrcXabc2OT2NrHl+Y19qMK
7Vd5tW69txIbmjf9+mOkitEcgBEVUL0vHa1bIUn3pZEri61GQUwQzgBj8x77dKKTEXYy0elBr0d4
67hRjJoaIosairVV0K9mN30fs9pCgxiKC8DjB7Cv6UXDH7nOEWB1zY7b1M83bM7uj4nJzE+0IW0B
/s5MSNjLCtjXxLicy0uyCQMOj9JUql1U9WGUKhl49vtQfj/GtJuhUQ8rONuwym5eytZWypJ2UKZD
8VUAConjrWGTHbVhbKZlrTvMp2kh8XEagWX+0ykiWpbOl2yKRIEtz5rCpapsFqyTdpDv7ZIRbyxb
30s+S1It8fmH3B3ynJHfq85MGNdp/j5ZNKvQY/jc0S2dH5qsUOJ2SD7bk2qpK8bNwACNl3Be7iyU
GAvkztUyaVpng2dQH53fPp/3HWUr2t8DIQkLJ3qqyluj7Q2qqTFItPVWfVGL7jYy05POlXxdXCnO
rdIJbjAQSDNU4WKFRw9wps5UjtKhTY1cuLx1F53x5P0yPJJbv76PK01JV/O0cpMwXdfxSM/q4AQ7
bH4vEZJET0RmBwVpXAZ/WT8rq5awLfdJ8tjw5ktioEOm387FzIqpCGfDwyex5aehD+T39KvMotAA
8J7VlnJDpNH4LOjNuWI9kRYjvgGa1bMn+UP3g42mkzvtZDJyVgYz2ZKfJ6niSf60vmFVUuXy3lg5
Y3wlT6axmGBDuYifvwXI9UoQxdUcnV6nWB+lk5wdoquJ+ZucymZDSaXzS3M+Fzw9dPi0kvm+OgGQ
KM5dFdu2e4P2sM4g9+BhcQ8W8lj3AuBKCOJ1hKTBLdj1FBbMDxjoj2sYmAZ8lhEvruVY0Nig9CDs
5W6/ixkLrQkeEHvWhPa6MbSx7w+AJHTvH4L7ja/DVgTrYq1az2QKCBHskY5fsX76k/ma8hxy0cy6
k6Ezp8NahbTPCGfuI7cjtfgKSkZ2kAjIXvRNNoDo2H9+OBCRqO43O4rzy1rEp9VkHl2Sm5cEYRPP
tJnb3HkApCNdFLSf4xmTFtFvWP+A9LyNw3RB+xxgJFXbMmYndR7vYSiNpo5Xn4wqbCVDDf4MclOL
1bNEma9cbMGMTkWu6vjV8jZS2p8Gli7EAJJgPautCTdfWQwA4y9SdwJKNdTWdmnvCqXKQCp8g3a5
N2nRBs7+EXrRJBz6Z6OoFNG5dVgKMmbqtHE58hGwefdGZybG03Rr5COQdOMqc0cYm0exKXof8lvD
LCrVA4dwy8HPou+AB8dJZepyJYYnMR7ercFLaQcntCda2CrrGRPyisiD8Fz/gQ5KEcjzNTVEQVYe
a+HkAcpJksQuB2+wwIdpS6blSXjzrekT+CVkbHkxKRiinHZNMAIFJKPa0jkjTAy/cMyWxE1CjE7D
tkpBce1BbBuFv5ASgF8WjDsLK+b9w/iwSF29IugeCIsDRgMWUbtv/5OGaK0rKHaKwHBhLgaVLa5t
mftP93tT1AKgPs/EzdXFEPKFAhe9XpPEx4AFgyPW+mbKgByjzCIX8xUXpXMWZTTeliKnJZaQdoCj
3lvLjQ+Etcpd1HioV9IGqGbNia0Y3TuMQZ/vGFMfxzbkmstDKd5iY1RffnrfWRAE8NlRumNs+dvA
3AhWBpjCQM1jw7mmzaSzRNLLn/Njd8gJ76VgwNdAzNCnFKE6dK3+ef4eLu47CbvxLqyUacPkExhN
PSh7S1VBv0fhAS4nxwk1BFB4PV6z0NDkKyOYrtNH7ZCF/wh+8L5WjC+/S3RA47DvWwcJ1g0PgbeK
9GUATyEHglwRBUK8u7Xh2BS68gT4YlM/ndtA6RMDfEMMpQ0C4Y6ZohrobWfozIgiceejrYxZJSmc
5RhohOQKNHHJvHPLfY9ldtCUsStIqlrC1aXAKu3tX/yGQ0JIB+ctICUbhtPYvCrjoRjV2/xDJfFL
YI0cD8/51wnO7i/m1LOri7yCRyLAJtglZE+dkFmDoUkxF7lt6HHDhZ+rgDT/+MtDSz6FGHArWCHH
9qkaMZHeqyV8XEjr0jWbfkLz/PvZUh0Ol5HxwGEdBvjL6nMhUyOQyBeH1qIfOte/86bhtCq6fMA5
q8PZma4ApbpMULuH11NuewBCT6E0BEIDlCniKzIjIZ4+TPNbHO0IaJwRFO7OKgEMJiTXrLM5z7B8
/jkAGVxS20Qr4S5GfvU1MmE2zKcsYEt2gBBmQ2XwClsjnLY0Iu2hTv0j4Xs7xb8OUgoG1+0L9Q4M
sYUpkeIndhMMCZ1NoIAoKWlTR2BgNGjcgOly5/XcVFfT5tPYE0RcKYzDuAEA8sOGk6FxjBwuARG5
1c1R1opOvboeQXX4+TQlH9Uj5R3tZD7Tu5ztTbEnKL+T52/4KmztcXdmTqbxT7Ot7gwpXfGbu7C4
LWTpljOJj20IdwXEsKpCEkcPs+wEMa3dg6BnxgGZA4Vm9Jany+ONeAXWu1v5V4Sy7eJ6IRPuBzLR
HumDwREqlZqHybvc2ENeNgHaYNzzxNufLoOEOev3GD3uy8RcyuxGr1fkWChdbZlu3Dy2uLtbPzsX
FTcqg549jFZZkDHZbB3LROEuqP13L0JAZE8BXeU4HVd6mnEUigmhokjiq0ineLyBwvpG6mv+iDGK
6JQqFwKruqvnnFAOSizhJ+vCGuUlXFgHfp4wP49xgUgOnVt1JuIMZZ1GcbKmXuV3J1i4Lk1yYh76
pXjP8zplirZXP/CWzRsyt01y5mxueV4ESwX2HIm3H6pr1wSeFr3OyG+j1CEO50KhiT9KebLmzbZS
iRnr4t5DpFfBu288YQenKXQuOGe6MNKWUwdSZpkMdzf3kTk+FmCNmKclBdkQQ9LbcbLN/EmG7ToW
4QBDUV1fr8e6VQlEskuU2kR2xn7xhfdSB3PBFhTgYE+Dhmv9cdGNagAZtYLqmFjLZDN0uEVii0kS
JPs9fcLjAdD9109Hfxy9chbUVdv5LOopDSkdW3jFq1wRbXdUd0l0BH5THBO8uPbHeA1AXwMDvanY
FEfMeyLfPMWE0e2m8j1e/kVaPJP4jkhmqsc3omHVxh+NJD11WQWattJjIgS4OjsVsMYJ3UGS43da
tDwvDUDn+xrDFL0DMvbLzWKoJdS4zabNncCCjzZaSNuZIsadFSKqvOollt1vKuhcddLWiptX3lP0
DC2EqskFIiUPXILTeoZOPK92odhOVsBBO/Zmisl8FY+RXxyOTDfJMzQ/Qqd6hAk46Yt83bFhaSGX
sceNCyfHwUu4wEZFG4xc0j8CEVgmjWgGmDPolUTYPU8tjkZ8UelNubRXiKp0rpzIvEYjM1EaGNFt
0Yw3N5Rs2/FyyK6L97r4+PfruCoh8SnNtVUEP2xvImPjmAiYr0teJNEiQfx+L6zQPjvw4hgQaZzA
+9NS7gWsw7vRpAexkiVW/RLmpvsEBQjovMvRadfF6sCjYmhnETLMni/iRHCWcdx55z9Zjquf7CLw
T/OL6G09eZwn/zcNsuPpWBrpjihh/AXl26lrRg4VxStxEwU0Y7KWItI9A7/+/CHvky/yh59X/zHA
w6F47XwvvK5zeqKyJgZu2W5BGaDfMise2bOdq528UcMio8Th0+V7IGsfm75DH9xJYOAPHlf3hSTe
cQkpIp/rO+ZGmzHwabspwt4Xz4knzpRiCRpP27IXZU19C4Wa8UeJfcdl9AL+jIUtdFwQ9xs3HPtw
JppPIrsY0LSHFYrQYv9eVL690L/o/BZsT9FTooidrbSv3tncRiOqSxb+zpiuVE3VndOz+ZVBELBd
cZq8DRqjN8Fs2wycGajYybkx0r6aDf18Tz/8jAjfwt5JAw8uc6e/tGA7iPIxo1HMm8dTE6/3VAON
zzci7+XeMIL0NSA+VsQPmK9rvmKaKpxWwQwHf19GKcbir3MM7S1iEnWPD0a5OBdeu6nrJdsjuceT
kE45VPIfU0ho7hdp4v4W4dZupjW0jib+8JVR3mVYeclUYyxvAytlgvoOaS+kvC/mrQgXLM+uBKxX
k5CkhTe82dLAhswbflGw+onFMWR6i+Eh6WnMeulQrs43MRbvyl1WrqmkjP5sTCh36ESuS/RS94ZJ
OY0QouLDwC/k3LwHLeZ1OdFTaqsVs3MD+N+fYCeyK9Drhk19HAY8nzX/RU4tsCzMbKQqAybN/R+F
sAuhlhXPYvfaXF9v995GNVE7/pyhb54q1U5hMASN1bVOCqEHK6yin7AMnjW9aMq1gqembthVBLX9
dly/mKKtp5+iekuTaOoIN4Lslcr8eguTVUBkh36a6BvKKVaY5WS3180C46R48A14KPknFWwPEnUf
TH92rav0QgEWCLFCBBn0n+/E/p8wnbYTOua23buZEe+xE+woGXt6pKfjf5etGrxPG5kbG20TMAW8
yWAkS/t/aWoN84rL19d03gEtdgy1j3pqnbHR0iFOWd9pBDrsx757Qork0MF3qkUDaRipO8g5wyOf
Rf81fC9H3vLlBodbMMUawkloMuo6msVKjopbUdN9uaBdczj6NU+58AazvWKVG6p/qZ7pJ0at6o1r
6GjvrnOyZfsDbpTEsLI357x6sP3D5K/9w733jxuYpOSj19n74fuUY2v20XPLb3OTO+DBo3aHQw56
iSAJEFAZAaQOME+wz/4/yHBil3DtB81MWxJ2EMRWcuSOCurKC0d469syfbExegdWrSFNyhh2n7k8
+uP56LfzlvTgMZZjZ5hZjaIq/r3Fmyyf0iV5u3zNZEddtqiAK3LvKdMpEHzUr3jXgXvu4KrbHqB4
kFpP1JuLX0zDOtoTBKCez/npWlaItMsy8igfbBbftsO/m1CG3wlUSgm3U0plQ0K4JQWaYf8XDE4J
UVXiGmhY1qKijv/e4ncl1++WyvECZtSJ8hr3LMF3BKqZBaovl2jQUgW4sCzYa7aexj//TVxWwTUG
Tn92SAHAqxM1DupqCR0LFOR7PzK4Szb75qMuI2f4EZXX6zt7CUPxK/JtVBHzvr39Z/CaDcBxUBXe
FgCDlBYJs0jxsYP2rm2bpAE9P02tkiR2JQjenulYb984q6Uo8G6QVIeoj2uUHq5dVmgJlPzCEJTZ
L26y5Wly0cm+mwW8hGOw8Dh4op2zWce/G7aWlwqzHTAco9ROAIWU1y25w2kVt4UwbBl99c8s4SOC
Opo0H71dOe9NUBvLZ+aJYIAXMskVN5pyTMIh5uu8/4av8siiy+mdw6UzEYKW/1d79zwSgdyj8QaX
g1htHTisYrChZdA2Uszb9XvvJa8z9B1jiTwjRD7HJd1+2IK03h0IGEhYpGiEnTQPv22mjPfgJhe+
mmZvfKqqHg5IxQeaS0dDqzG8enwePMV/uBD5EIXcvanCYI2wspUWl/oYyjJ40MpPGSQB6gDXoh3c
RS6KD7ps8I9N9H5HQsutCoOKfdnLAEbXABSmS8Y353g5PjvepgzSGD7dD0bnRrdLEpqZ53V3Zpn7
VWKkPK6RNcK4OqGNfOxUx83ir/dQMFSW/KvL7orQeyksFKUeSCwuP1tP9h0R2+nFim1fcqUPszVr
WIH03ywpJZSpl7p/g9Nf39/Ajrun4jhr2ktRKik2yZp0JAiF0Wr7JWN6fHX/Ch2R9f/qDuRvgOJP
/eKKymM0jduKJ33BCCPoy00uWvkPjWHjeB4uMoroCBvp/IE6Um4Iags3WNpkhTEpy4LOr+j7356b
0xcKDSe/0Y74mJ5BkREG16Ya8O/fg640Gw3XInNZ4PHaafC0IVKqAx6XGevXYVBKuYqxcDULCLoh
FjsCQ8rYN0gLfltcUPZn9TeNoAkI2KxhOLOfvaGH3A1hFT6+zwb3htK4ct/ifeZUMyLaNtvTrQOy
NjJU8q9FGJAsMU8dpTXIvWRm9SOGGNao9H+wRNvdEB9JWDHYXgPIQyKwELCtwtsFB7hEotKLDwAH
tuExLFwQElBrbfQikxqM3DPak/9MnPrwhqEBTZjR+Bhlyj2ib0ywkoUIF/0vco7x9fa/X7TFiFQu
d4c9rZuWXDKu6Wu3UPek78fhJlolTgeRST3x+T4PBpPuIszWh+KfHton27iF+BZypibQdHja/KyG
78DqjwARrXv/O5778XOHIvRPT4IQzd4WrPruBBbqo1LglgR7T5GCWjp3cmwcRB4Uxivtn6gVD4bX
TLWDuRLTiZw6jgDFquPHF81dKIAxESV6ZHIo1XD9ov8mLuMikYVlpNIoW0Da9FZ8kMblZb4/D4fP
REzRtD3ZVEIqM62eugaJgZOdIQjEuyWGdqlhn61LH7hcgM8f3WxJllcBZDgs4Hba861e84UpzowF
M+1OCDLqsp0M5fF7pJMu7xaT7hqyCiEn0pMHU5T8pGOpdiC7rMEvy0H+zl/r5vqZHElxW6XXKhn/
PZRFZGOAdGay/6YHl7LUsRWfdAspUQkP9Q6fjvJICau/7x5SWgpx/lPFWOKFfVqVLCmvM1GxJbs0
glN2GlrWXme9rE4fI3F+UUqHVkR+0aLsQ2RX4X7lNtHAww4RqmIf2RJ+BYFsMfRRSmZYKtwdCDht
P3r3FXswJj+4i1V38FI6ozVGI9hViZtF7rTdlBVMYodN9tLayVp4qiepVNKXfwPAqoaM1h6x1dLN
TbnGqtoTMPJLgYMJBbUi225W2cEPt2MkaJ5yPMYxANYv9YGPFttJFPNUs+Qzt9X21mhM76UxiMV+
WTbhwQ5a/Y50eTdyJNG4IxsuW6Pl5msNSA0KAnrNWZ7cZe61K4b/8zU7o8LC2GgSnoJrye0wDLIS
khzuNlJez0OPguitNeRSTB6o20zgrKc/M1q3NozA9AeAJyTeL/rPRUwT5ErKhy2pUgAkQndnB06B
4ud6HLBbqDKxNRF+MvoyqtytMTqoJnrcGXbopD7Iy8j/QNG54U1qcGY45dlzWVQymkZrMb8+iH8J
RTwg06szFpyhtANxc23w6y2Ls1htb/g4gV+CJHCmcdVGuaSBjjGowISYyV4tzd8aCpIDa4aBBufN
4e1/+L6dZZMAHM0Wu2vMCmv47c8BOTuqoVoMk2uAxYpd6RbgjT3m6Nwc5LyWW5IA9wbC43cSPxPy
msNTX0b8SDUApUj2BUA+RHO2u4t2Fa+jEGAilvb3d9BA/TxvytMSdxjoT15HPzipPUNPO9/OQjuz
IXaguPQyhvMX0xn/J9hVg6CKoo5ClMdKSI2N/7O7Wcay6fLmUxQ94MZzViD0LvRbp0Fdo4Qx/E2m
MA4Y7S62vUnXAJdNz9QGZ3+o5wgjBijWAs1xRzXlPPmCHDhpBKPdOMUhNQOjbXzfyKOf6qrnn+Vm
G0QxMlu2s7TUzKkxOTqP0jVlDrLo/00rck3JnMygL3ksKepfTmsRSzNQSn+GbU62KX3krRZXFERy
vXXMuaImwkgXem1eZT/dq0etk5zzx47cP5I4GjmJcuzo1RlH3gjxIKWFVEk6VKmjd5yFP83aj8Ot
HlIBBEAJ/EmPCdUWesrHxHBqrU4UqUna80h/fKBDROtV5NYpMXd5IGWvOjCUa748MC9glGJIXwMz
oE/YyT96xuknRQiNVCpqasvXJL0bgZoBcNTyDGxAO9d5J1yRioAQp5RUs20W/geRLLSR+Kk48Hwv
opBwLWVODdGNTepzdYfPvBFVf7SWTAWl6jfrn+ppaAnfZ7pGnrWbfbHjtlNQyNkzwzfK8jlO6iPx
n2XClSvLINMdqhILVnUor6yN9R80B1ESfdH/rr6pgF+4pupa/1wWzjxVmrq95CugTs8OxgpAPyPm
oZZ2HQu/u7hqq5qvBBeqiGHcc1pZN/MGJMVp2hEPfYCYIOfMEVo6lrEZoFCz2pqK6cOciWca0tVW
+Ze0Cq40X0Ms/Kzu62hEBtlB1yqZlw8bLA8FknvCUWmxEyfvoqxhK5xy2JrDuclj7rGWH5Fnw4v/
Owlu5+Wt452iEOrOSKKm01Yf8Xd9FJDoB3ZS1ZUWdk5D+sfguYRdwVoMidevVHx6yMnQkdbo75wb
oX546AYNUOF6Sc3xSlx+F4dUrlVTI2i4iqISQrpz3tSiVx/nwlm3QxIKBzuQqT42MkEtljGkvqrJ
XYBYagDTOJdxEyGA97lhlGccsuc7VR37TZV6upFyCXL2i65Yt1Vj0FdpXxLVLrCN+OvnxSJtu85e
ng5Etxj7brvzAIudhn2MZ8SCNZCXDXfxvX4W7Qq1wIFjcGzSBl8ACpDT/+UfWzjzgMS1AJpHHvNv
YDS9NzYyMlOJ3mB1O1TqB7laYXyNMugQsZO3OhgmVLTM/MwzkYXJOv72AiGw6fsl+EcPX44MTJLd
3xD6RZjGzX1Eub1cjd6s24bYQTyn0cFpkoN5S3W2js7pkg5J+I/YTirdIJwnKE3wmJdItvuRr0RS
xlk19669Hji8byBenA/8tgGXFl1kpal2X86pZz3S9sM1mGN5lzyA7eOHa4VLeH5TArQb9fsRZi1R
NIj0GNmQo9kba1aI/QAXyI+YUGHS3quk1Qu7ATr3ZfPdHMEZmZFhDneKWmddx644FeC7E3KaH6ig
5jZt9Hd7LhEDfZScI8bhRh/3tdc9TUvOoIU4uvfMtDjiGKCwAyzct9bZV4RFj5B+2F6FPxhs1ieE
L3kxQwrTqNwolp6CUbS8GtWH4y+hCl9TwzRVSFAHAO1EtzccRlP3TxXhqdQk8V33YVRlZrILjU6s
DzFukAm5ruwGHbk6XePsuXOd+4SQ1rwZP99wN5Ifk6HUidM/+lM6eC933OO3Z6gD9zQbBwmzhPTW
p8TNJgjxaAjKiepjZKub4XJ5teg8gXoRXIHDVVO0vN89CMUmr7MeDkbtCQFI7hDUtQsrwKU0FB5w
ro9wEuNsfsX7P+i4I0TKVWgKT9Lm58Q5+Zqp3EMbzjo8ujoq30tPeFYPzUvt2hYXlcDO85j9Qs0l
VPNKUJeBISTZeODqhhM1VOxOUgNGJGhQwJd0Ks0d600ZzlgMdlZMwxlLbvpSYqkz9+Qtk68MgP4F
qZUq9FVy17fu0YtxrL7hKqmx05UOC2cWfjbGuo/7+QwMjqnvmQmfqBZI1fxwDkgxnnH6i776fxdM
qT7XXyZRs76vLj9ExvFqGuHKpBcVSa/wzfYfOup3s0tQaFadJbBw4IgzYUbiXOkJmRpEToBLdgNV
tkOZ2Ah/vUWy+6Vl0OCXCHiLqt6obSFIrPkU7rR7zfEdLHtqhhUyL8FAPkrB/nrkH+lUlz+sxXN9
YoeKcRwxdNZ8ug0gOAOtI4ynP3p/4L65q327vbb8uaT7FD3ifIyZY5DunhCwQ1rCWce6W1SUWot7
f1hJJrKRPNz2y9nockOqCWPobl6tBXjHVmSZXWWlsVTVwnkx7BOcGDM8FFjhEykjQ7xm3AM4QeWI
QtLwlpHHArMayxEl7vRziG+pCLCc/k0qcQZk7io8zTOEWjZ42LmVxezNHrmdlLU5a8jKL1TFwkH8
CXEk3rYStDtNRAq5BQ8cWIrYWkFyCHlJ5OE1iLfyjeVrxgnTDcQSF/ueY7kZPsSMSQlOC+Ho05I9
7sbfXZR0PIGloaWW4tEmeLkjjfYlFiq65SC4iIdS1RpUXA9vXS6zHg2HwZ2CnSC1tPHmfV7tFWrY
sFXlPt/A88+w1zGg6qtU06jJdj05HaSAPclueaw54EMHxq6B64PUBETe1ZA4scOvlgFVrT8vjXzM
pZe+gfwjgxbZ44bjVI4VEs0QENFhTG0wM4f3CuoGruqIKo+b7BVjkRiXSm8WWwy2aWe4HzpVSITb
5R55a4NM5roLM0neaUDdQzJAWmmAjMUXXOMl4RxRXbEoQNTn07QyIv/4z1eB/DoKZyXLg46iYOuy
4LkvFgARm/Ns7N0vqXntPXDo75Vp43kYjxtYxZZgKGIhiAfBMVH3DV25rHTofEYJSWTOfFNO20zT
qZIq6dqxA3U/2z0EN9hbsn9Xe0uWPx6aKU2SRcKxCMjgC7sQPeCbJTV2fKx/FF8ormGBPL5NSWYt
Ue3Nma2D0akO3sfOwwkhe/p1sYCVWAkWnN6e6m/E00aNw9/2zWNIqZvx7hYXJYgGSkLDjlOm96WL
Zlztj2pocPshIcu7RujKPkjB6XffsBG5wqGsXVg8gNfsCxFiaPeqnnYVIVqnebRF5Njg4QTfkCVM
4Mf54RddN00npLKfSsJpB20RfTNU5ZoziEJwuoOy/Ce3nZdlPKfZxhONx/GmRYZ0Ih24CG+Gk+25
tNBFM3uCKlwS3JzDdhju++EC2SN+JJkFZ5oTiYJBkv4BEfWd0QpHNIbzgKKh+Jb8dD7rk3uci5Ac
NSl/oOPQICn4TweuFZ9nyehszTDSuLNS5E5AWuP6QzzDqbbm+qbYhLH5bOvKZL62ACFXjUNqTPRt
vS283nMUAyeowkEQ877Jwz1frpH3vxDcYCjDz5nwJ48FCx3cxIvGaFpq1YJclTVZZqjzUnu43JBM
bS/iacVGA83y0w4VbCrfeISzJVV87mF9E0zEgDpl/ZpbcHMC+DPGOA3037zjcAtGHb1ak+FNzR2e
cNaSUwjRZX5sYYXqb8tOUg9GzFqKpMZHGLBxwRaVGPOZfk/KrcpWdrbmKIO+smPyqfLGraTi718l
T5jYgzx/RVBxkRwhXFZ7k1hSpiX2czIa12KqZ2b/a1OxDp6hgvoOoLXQ8OpDETGL3DENrmoh1RPA
9YbyZueWOV4WixqlqF7O+NwnQ50/8Caqdnkq7HoXvIZDdvVQIyYLW8Q/nokUKk8vjLU1B2Whawxo
aQYjPbOQlYInt1IhgiTFy/O09vPOQtyZCjif2yDjelp16cHM854b+9VoqCU62l0j/NXvKzmFdTUC
l3BN0c0AgTLpzeRXmiunIM9Ol3BnjZM/K/HHmyymmSekM+shg5fVZYVYYSstcAjRoMMF8DSHq19A
3d28C0Jk3Pq0zninKriC6FhylQVvU86xFo5odnBNDVKVT/LCMQPouH81csb42UrcgUrGkPxDQQAZ
X3RQzNpXXeYQBOJZ700vTPqdEu65bGvnK+6szg+nj+X9qIaLVABP1R9adquB3crMxn+xz6dR2TvG
h1MceqShMivKsqZU57qgzuha0ifw/XdemEpzCDZHiwzgZu+G2ZMd6WQweUMKk1GTmTjsK0SZ+B+j
ZAUlKicvxX/i5GfuwoblrXNFX0SXVhNjSgOyA+nIqn8lotb4DWosaxUANj4SJm3IFdUlyIoE7ajP
irD1O01ZCe9qjjJhdtxFZZOs/2bVa7hCyF+BDxpuebocENJTKUTB1yh0z3ZgKGrdYpHecs6MF815
mAytC8INIor04Km+pavUz7TA5495ZGL1nGKTA6VIQnxIyZbAbKhs8kxFdwRUxb8jKFMAGpUwUA35
GjNQ2hWiEzmC+9aUoDiFB227IKs0NxxsnLC990pKeghYAIMRPWmdL6o7sTXC92bPhRJWNjUwP1K5
IotFpJhT/r0TA/ez2iSnEx0+aqKNxadmheBLld06r1x+L39efqpd9CKbuTn5cuL6K2Db849ZF2ew
/4fgn+ZUO9hOwpzmoxgi6zxvbwke/Iyfe9+g9I9QDzqE7pHTNF60vw9BVEl1U2bNLk+VONC89ibW
eSxvcJ2g9u8VbfCPZqADX0kXZXk4y180t4LvsT3NLT7yPRD+O4SSYTbAhjNCKwEUnqdYM0/iLY82
mJ5e0pVzc7mI8ka2zjUNp31F06AszUUQntuWmf3oRa28s2L5KqL6g0tAX24IaRx3KuzvSncd1ypZ
ab7pUjsUL+V71RVACvlTqIxQHwulZe80AWI5j8EXzqhHevKpp/zYXuE+bDJHroJbtX4FMkfyg2mE
049moz4HH4yM5FvCbuaHhjqmN1U5nY7DHsNT56LulUyiDPq2wbibA1zophzmaeuoItsdJ/WiWKCV
jjBmA8EThZzkbEfoJLNeqCWpBgtSMOc/VC+LmDm3uckhk0Bdo2MpVkkcwdGFL0BKSwumLMH3M2Qh
ZAua2POXcnq5GnmKCkDXMmIfDgdKjY4J3RN0mCUDfFWYLiMe3GoQSGhrdbSOmFfbBN13CVYZggXS
G0TONYtdZWw1P9feC7vtURGlRwg1CLLBeP+mXT6/V4pv6mGsnnsa8mQaFaeB1WzqKwAeJJYeoyTk
+XhGpZetENC58Cw7nqZRHODD7At+cBAUucxJN6/qfnN8Ja2oNBFWoq31n3iaYhVBtDPY7jDo0aCX
hWMtTyKNA812G158wf1h3Y+P11rgTevKoQkanH2jJF2V2acCJ/dIMPa+ycS29gQwEpOXjHmI5Az3
NviVpoScqGE951eW+dPRs+jlzSsGETW/ykdxpoFArvp4sKocNXvKmzMF4BbKNfiLXO/vJdFyjQJl
jmovdfqRAfRYanFxCjZHp/7Hgnit/1OYv0UgsRti60gCqaK8DWaLxCVs4ILyNtUMBaE9VJKMFpK8
bWED4vhR8ddZ10SJApOn1lw+0V1o9LYnHI5im3eAZhQ2M8QO5q82n9B9B8KvsRnGdind4qYkNEgM
WD5AXZqtPcq3rxOuHJthIlMsu6b25NAGWdoRtroCdsL9va3hD2Erupl4iqL83WXhbpq28u/m+GzL
/HUGmayDidVbw6emILduzYqmtJiWlm/FKH11Yuk8zImo4tHbYNaPUpv53rD5SJiPgEAglN8r3As3
UEzL6vNFPHaWRLhAnGYU1u/cSBIYAQKCnr+0Sy7PzjGgUXuy0rNQKNChsrieI9c1gkAZfaIWzEBr
uyhMTxZD+NkyjOQk9+/wcLjgTEPgffs06TUt6QBeLTxr/FiYLEglD4miRuYwcC46oYIx2cI8rYAS
krjckkRSBeoftLX16gvuQ4xqEyUMLlAyFlYdWYv91ZVid5cdQdy4aA0JeJrpO4DpWk1lh7oDQuji
KDT6F9hJaDevodviqePVwUhl7W2antOumct4f5sYMLpqUg/+F6ez2GWtqs2sVcxWhmTUPSYNk8Ou
dr3z8CAeOmMr8uF8gpysxd8tirTYV1iy8q2y7doQFvLnZhy8qgkC2KhyLWK58eQfq3rh24vvKT9p
51FL5HHLGB+zBOuLMk3siy+tvNSYcRDsYkeSqmsspZ9BN9BRAmSw4bq7YY/PSwVjtGE6aFjRdv39
vmSZyWXTSfzrMI7gC17CSNtPU1vw6qaxP3x70X9hMHVYdyM7bMsOP2zD58/RSAM5wkaSa6JKs+Dn
z5GAarnnZhQ3ZLGF2Eg0oXvzrP95x8ikwkWAhAopMTNRCsgW9qwu66L1kZPJ+/3MCQLeceaPO7+2
HlCvUaoMkqnMnekkHY70NMQaQHZi5hCMUfjS/qKzG04/4vrBSVcj/MNhy5Coyjg5zf26NfAFAmOD
UUJt/WIdaPKHrUAK63+pGdCuVGh5+xvcamff3oMPjGQXHtzD9QnOZV6cZlOvBd0PthfJQSVxXqHA
IpGWA4VFtVUlahMif53olrkFIVAjIXmovSOQsaOT+gywtBYsJ+QXqPJ9hR/xVUlLgN+pyqqF1oWs
ofkQ3yAlQeesc3pS2NbWZ1QWhIUm1rKBgXsH8bpqWq3xkm+G0om8gp3hNEhDPvPXS31cytKetf2C
hvbF9CcMRuYRqe527pgW7L6DqBvC1FFfB8OIhpD9+7EBKJaks7QlACllrocrIPYuXxOGl1o4y2lO
b661SY4FbrPsTXY6xjxAL0+D+Sy1THRSYxZyaSMssah5TbRtGgPMK6lBlOegPe0rmLolofmZR5WX
gxwn8N7VmZNNvjN2naEUQBUY0ZJh3UYYRSIPhCUPrmKtaNNFSaXw7RV27vqlfj1N8CXHB0h/1xvc
l2RClJ2/mde1q4HmTzr429oTcBcuUAKk316+Xk7EcITTUSXzlELBLLzPegyBZjbS64yrtR+72WTR
+9TKguWjZM9jWxXfIozotfyxgHC5KQQ5V52CHHcgoCXsAd73o3fKUKRYDcZNlBFSGYVcA0nVeJtz
JyDK+4Oi6DqW9S/md9RmT8+AH5UysOui2EZCliVG+H7VXLEXB/yw8xbD/g9/tvNEDVbHCEoOUsOF
sngMbmw8r0/3Cj4mK4A7f/Nl9fyJNuFzpaRuaqk4IDuzIfHuX9B5Qh/l2Vz6FCchLIEfko69mfiC
lCUTZewa8bbn5HPOHCjo4HvZwQEh25ozIuIktNPZJnsBHV25AeZPm4eYH01w1/IaGEyV6Opqp7m5
uuvbMxdREOmVcWtw3/urcQOJyqCZLECIwNGF/9IKbkL0M59URfV0wU4iL/LjKuwnVyZp0+KAzDRI
t7i8lgc+oXouTpfyFIM8pjsk0XzzdIYbqneP4njSkhgAzA+cvPrMJ+AS9qsOfDMOvXXBQ2Hl2XVS
EjnMzHdyYGCbdq+FPCd6KesSUqN2BldZCXTzfp2ZfU4PgpLhtst5w7yN18zOleTjsjjmPr+83v0q
0P3ZuCn4FxKkOWnIInHwBZvk7namclXPr5TUlQ05FEGy6ceRJK/e1Fb395qYCXXKyTwG8mbSzmTp
Jnzhp4J4jvwbMeUPpp7wpUNrjVcBSyUXvqaXrgfXKVoilwzVT3nRNOQkdvmo9T7J64ocS6DOnhkw
uSlf8Al5genumH+E70C3Aw5ZNDPpor/vKygdA8xu+X18IxnFfFqd7gEETCdmXU0BhxHLYTVaoMpY
nztTuuDxFxUt5VHugbLFmNnQIhJBDqCplGAIaclFSr3HeXYN/VJdo4AZu5CjncHkBY8uM1X8SW2q
9zmc7IGa+SipuTbBGonUyRlFEVhJirol64/unkk7CXt/9ZKtP18yBENESNFhpEfV44dSkZ8Gh5FS
jcbpGodsadqivrHppos0VHv7h4LDrJjpu35yj0fTyqf6Bfc4QurUgN1N7Ut/Xj8V/TDqh9Qx/IqG
4vFFd2gPtbGTHQUOmT5BjJZ/qEX6VmfvDUKnIvngEwnI+rc6zgAdaXb3hrmgJnT38+5dLFl3xgKe
iASAsDbd2rtxTN+ZZxCgA7PGPKnDypAHWph2n/kUgjiEG4x9J/doLwo73+kujsCxwpy/G7zV+KNq
O+IipjEgzh0zbPYbNrOSlYLugX4t8qqWaOtLApiGoaax7aW/4a5KrtLFr4nAT8r35ARgLU2+mq6V
1JzAZtpga1xTrNxTpjjltkl0gXRtHDU3btza4S6JN0KgX+uzauBPD6dvSfSUVNrxmTp/zTj/CRpj
6vXSifW2BFVzclfzebP8IxG2YlyUuTtv1UNyKGNoCTPrsYryfzdtyiJAqvmvUcISOagxEdR6Pvkp
qqqeGtmVYBn1FrgXSgDDgMIjfjgrp8aMCTYTnMw29+ryENJW05gRE1hJjxs4aI+p+qDau9801DEb
enaXQIkN+qPtp+WzslwHnypBx9GFNs3GxWQB9Y48nCGncH+/M0I5D4ApWPicRW/2Wj6SsjN0SPap
Y/FiQjQBZ3RE69hgxWEI/+v05lNM9yUcOKghEEnZSMhYx5ohskzDy95jRY3MhBoGGsyFAsOSWQcz
RDEbG2YD52gr5bF1JU5qZtQD2Td6YWtxq2W4F9omgJB3aysux78/pCBCYVHzdoG+FESsTxGUF+gf
n2/vswVZJGsfCiCyrDMUbsWea/1VU8ftAxP4aYZIhXgMvqfqrs1GFDacarG8l9qkBvWBMX7VaTN4
1giB9AUcCWOZHH4oOKebG7I19OxTYVL3lBwlRzY+K8g3uzK09nu0VCcpWr2VP0BiRlGZmY0JCjC3
lAQT8YKRt3zJmb/qVgwQ5kJ2xGKPo7uKJJqZpMmYd3I/jdNm0uim+TdRMJLsG6BU9U71USDIkUcd
dJRvv7/bDRPHShDGOuddAJ7dO4QZ8zd4V96N3rxhP8yONPQ0xCNIREdHphtDrLLQ982af+Jlb/mk
pM3+uHAQnXZyt/xOLpkGzKsNDN+nGiHkyIodRi68H04eAX9vhv3tmyNBwoRgv0BejjpITtJdyium
GvLu+GuiOk5ZsuY5GLpQWq7taujY4kmh2MZHw3MQZ4mb9prgyf+y8L6JcJ9pQT9ybaIbGogaM+GF
w1QiZ0XUOZwMSqh7JG9E0qqx1pLqL5EMPgB0kJzni5dwUZ/P0tJZWFnZKhqP5X+IC4dPF8L5l531
dcCDgiICqBiY6aZ7Pz2FuIrnXx4rmSYj3Auro9daGw7SBoF+Gza208JaPEA/cF4us7hE7SKI1PJn
i2ANn8maYHW2lPwOJOt5/SfXMfacp5QImCRsMRHUD8yoZNf5Fx9X85G5BLlf7cp6WefiLGYmFbgA
lQ6aG9q7dVBoRWWW7ioSmWQRbIo72A6JOLd5tEpGKQQNKPruZwuu1+PFsfZLSmAhs0jTE4DT0LxH
cigLCevPO9Yyggy9iWr5KeHGAw0dV2kVWju9SpOgabY5jXkMpneAwmgclT8mAlQvicR3CAwaLTOS
jPwiquqa3HNL/DqBDSmlwF34xscSRU44+kX5e/eyoJmH1oMy1ydQibSa3HFBkpp+Lmc7fvQZXH4/
SzyzM7WVG15+91J2KQRBk8Bpx4HhSg4uLyULRhOJW25ckSq1XYXG7o3xfNnvNjhGPPwW3ofBhQGO
p3c5XemhHvN/q5oOMsUBLfQHHRfH5Z80+3SHxKecxxPdTKFdG0RllWyZiwJfV39IqgW7oZQuFz+D
F4AKipU8k+RkgF/sqY4PadHrw3VwFfj3DR0FubbW7aKx6Wb1MBAm9sinsE6mOzkZitTYUi79S5EO
Inn42wWS7AC/OeQ3Gegg8pXLIb8c1cbkYZq8aaLVtAbfpr4LrTeIAmixxQ02U/3HJmbNP8b1DkbI
P5AblNy00a1DzIpkApoWshU6eibI2QSoW5sVDd1ZHX84pLNkts3VQDeGyGdXdwYEaXqNMTU8qTJJ
n6vowgPa32F10rSjdNVmD/gj0ZUjlN/OtnjrtHSyRsSggSTXaYhyrj4V87sXHbC6NuYarspN1xxE
7qzpkTJxI/9RJTmDRyHLujxL6sPqbkmmONt2ZasyKBzFwChh7BmhkZCmDDEKIJM2mzyVBocPvGjB
9EGKW9TMZvZoQeL8Xb5b0eya/BLjFb+aFIQpxXMzXZsQ564L3iH1LSE8CJGR9lt02CcHdC2BIZFi
dU24j89yIARXcpelloC954i1kyyUg8OIS6YS0OBgn5K72hnsP3tKYIcClp3bCUUC+mKR9u+3mApj
wBe+74kQsfiDZap6MuOXYKjjSEtU7GiM0YJ1QaHws0CdFrP32459vkRkr6n0uxOK6VoIbjEDmBH8
0fJE8He2CwiRRJ0F8p6G/euQPltfbGIlFQagUwhGeGE5PPG5pXWdiHovKeIfHt66n2T+XTDcow7g
HhHP5XX0imyRLGMPLviex9I/U+DD8oVIk5GfS7HC5S+VpTvAGve7Z2bciQ+x27OsJ24BaZGdfioN
tcHRmqpZLT186f1oyaJ0I/BkeOWKAg4yn2LMP3hsyWtKGzM1BbOzhZSwGg+24kAjabTfDOJu/9/z
xbzFwVSaGAFHuILfIDwZD7u4CODRbUxB++OaFSw2Bxw7Qgt1GEc1B37lz3pt18+YqJg5nt5CIDIa
MHRiesSvwcpPgiXnXY4+edC3VoJBH1u6/nUWVt8vlUF+SVoR2CtJAMAsuOy3UzixeFbweeyxt8V7
lI6/pFQ+3I3bITe3efpUUqgX2U4vk9SGD7PV53xVoe+TZ0U7kDQhfEqRwSIQPRvS4VNDMnjqTvAp
BMXFJwMUQwGvABHTo9cYxgfqGWPd6LXUJzdHMwKVqNpLY5IjQPoz9BbBFeX2IfuNZ8Fp+TC2L0n4
K5fyqlcnP/qkywD7XqwVrVngybVHNk/v1mGiS+9xfU787WG64qL8V0qJ9tLpLwPVQz8vng0J1HCH
WPiyu2hJ3Z893zNQwtW5cH6NLq9cp0Ladhh8MnLAfi6Du/zM0PU2mT9pCshhHcUWvhbEXoRxeF0L
qYbdQ1WpRItzsshKrFviWQA4+XdKjVeueT4n1mEW9VIH7L8i5rraN3MUI3ZGRDqa/h48DyKNXANy
cWzeL2QrOxwrz58waKzwbuf6sGavcwz7iiWi6ze0sOk2lSYUgXzhvZ8WNoC+faSJ4NLwBuDRLNQx
AvBP8p2Q7OmvzJuSyou3MZmfordxXY5lw2wW85HKCVdjRcpc7MBS4gA5+SWSFCl0oUbtfKi9ii7r
nnNPcEmYxi9qsYJVcMAx/x/qqhAzDVNPzez8dP9ejJ0CxtD8k0TgS6/s1AdBR+TGJLrOsF7UYPVw
PLfvC4UaCU8zdeaXRfvkT40Ll2ji1taez7cWSWgJS/DJPpXzuB9j6G92IYaDfDJJSxdCekk3bykc
aGOdOCnGlDMS0Rx7QK+4rp0GPzcZzrFLZfbFqJqBNBPxzcG/DaYAtP1hMaqlzaTS0rRJK3UW+/lv
kgRPqv952+W/6qXCvsK91qzZQg3AM9PMJyJlm5j0cp0+fSaqqXMg67LIPHKHj7ccEKp//rOobx9a
ozaNZmyL86oj5gRqwJ7lnA9F7CgfCquE3CRsZmlUPLpdH+aZz0EyDuJnzycsrdgd1kzjUzAMV470
JZSj6OVa6OCq2oDC7wiPojFvGYlbUOajbT8pVmbeL8Ab5XtnmMWvlNAk0JqMtuuQPtQLhZJoQYMf
4AjWKf2UZ/qk9XRaCPuWvYDH4TQilWfGwHWBf0sbdAUCHBnGaaew3XwIcvB8xsiadaHwunTUy/Xd
MaVOQnhj0LmMZGBBMGUWkEyT4LcW4qHHOYlOuKQDzKkYAg5s5xYZxLF0Ygrs2+dVS7HY2leYuSr/
Vw6C5SCT6inb3kQ3BYaPqicUKo0gAvuFgiQWQZVmEoh/VD0ST3UBe8vpKAlF6/FTVdh+q3byzdfc
NbJmFF4mw57t08BTgv4ES2h184F5bk0VJZjulHCgI0uk+11uzt99Hj+H9y4hAlgF223fV7iS8Pgn
ShZ/YJhlIGcuQ+TSrksQNardSq8d2QuUshNSG2ImtM0Pr/YO377Vlgy0q1o+CcLdR5DhV6uzgpgQ
x/1yHw4uBDsVTYCim2ab90uyPW5UjDrcdsLb1K4RFmmZ9Qm530zsSBMgn0xq7H9gwpgJBgqbdQ14
aYdospqeTB/NDnc0fhe6uddeWh5IhL0LpmAb3l8QTFHLxaQWCCN3EVBL3DGn9AH9w0g7U6bOcko3
OsNT49ZFdcB9cGKSY1Dt+rJ9foWaV0WS++qVwJXo5KFwkmGPtSUfk/13Hk+KCfKjhONKhIR8etFj
LVE/5fJwxsqbUD/NwMVcdSMHrZk/wk5aI9pk7aPZnHvNMPB3U1ikvW9P7a6Y3jj1I13fn7IoO220
ReDhjZXmJ+RQOmjFDUjtTX4eE/Y1jMWNbL5kX48X6pOMMQd3gxceR2k5JjSsAkDV5JNQULHXN/0d
SIsyOA+ERNxxgwrnoxzh8Z3wIBFlZs2ritW4flufB3pNyaFQQn2R07nMRqwew0maTk5bZT6GihxS
bNLUKBxCBiqikYMi/M2VUqbfmRUC7yEMGzgHAjUGXcA/MfwFYgwFNwTCLRwnRTfo546GhMoNYbp+
xHJXB+llx/SqyOmr0XYzL3ZnFskzgWxt8DykqQGZMEwA6jN5p43xUIAHQTSH7OTKPM7IuyGT7RFu
id/i8Z1B0GbQ24nViVoXbQmqQWlh0OxwljGNGq7aulo/rl85PontOWwc4ajoV8r9wfakecAsbSzi
GGrLH9NDk4ZWNuGNMTeBkxy3wZu0dM8oINvUcUk1oVMPT8HqstaLqgn1XiU9mIFhHxyzB9q0+RKF
qTtjCqywjoWqaIJk3ggZre5pFZCX5aCi1KQTqxBGdQI7vXxAGifXtRvzVAiiZZzlmbLqr598MOvH
u5BZ1+YWIfTBPmB54nxRFSXDejU1m11U864Ii7pdRDOtv+oAv6NLHDeInsCiSU7ANKyKrVBqlgtH
3IbXMgkB9KucKLBRRhpJ1uotuSQohEvZpUIA7pO4P+NT8Le9wpiU0EtE1XZPSbNZ6S3sxjnCnb2M
1mvroXE3rWC+u4yOdZruzUigBi90JY3TiRrYpAW9/LVCM/QzA/mFpwZDdmfPWUvyYnmCNsRMi4SV
vcltiSXDD8K9wVnJYWcOdlHm0WLKud37NryoGbm2R4kp3kNNsSbiTRTtpsmyaJTx3SV2OhzsVbba
tmqEpQuy1uFELQ2kWkdFYtRAQ7e2KsNMlMpckxtq7vPBDvAg8kkGEmSiqk0c6g9Wp0DP85Y9JkjE
2VA6USxlBj1WONom9Y1rI28sv8RGHfsXHbV0hrBgZZAWJZb28Uwi68L7auVO9gpi//PyDQn8g+Uf
9XhQ6myz3qQaBWuLtbixM4ZI3H1gOubzrA8DRGCnMv4FVNdiLGZeF6EiQ7S3/KCE1695zQYVwDRr
Azl5llo+IHvPkPnqZr7q/x9y23u9s4eDlWlmB29QC58QUj0xUXlDMYPt3o53mClnA3ir4N+ppe3h
qcSbm8usCuPky7ahl/XzO0gjeTXAw1fT2NFamIDBB4R976N21sxNLjYNJyqBWewp3RTdqpWjMFQv
/euY4Q+kuCowINZtgl0db85enKXmRBbY0x8hWNaShhm12UF5QoCZuUDdOrbVHczdHfUKaeA8lCpw
3TM25fD4exF9r5ipjduCBykE0r0CcqeQEVY28krHiVDUbTyfGwWmVxk5EAh6XZMB3DwEOpzIkcR7
5tQUMTsL4r61hoy4Tb/jmff5QeKElCAvUMppqMXRXVDCxNroYEZbqYIridwC6gXaFXaR07NLVOny
Nbjm1e1N97/wF1bC6q5KFULcmp/5ybgbUvLRfO4mdj6NTuJLC9CWh0+TgswAQbE2ojBsDgXQZM9U
JcYNPlGJLevCdunrVTrTvCf8F1NQU4ctBZLUoGETeAem0HQMW0sE7i6a2rTy4xh0H9ZVjCnxFnig
MqC3QF1zRYh3YL/WTwCNP/liubWqTMzOf4b/oSxRYoAB1RlVdrJSr60M/yN5aqEqOfLwFkhafPe9
xAFo7/VM+RCi8rkv/cP0LEJWJEiFI9dRehoSBy/AFL99yw/Zx4mkhfL1ZiK0rRYzPIk7CoD3cqQw
z50R4opInW84ynjh2E7Llyo/RQRKmQ7pf9cHAcvi5dJDxIW4VPKpDwCpu1b5JUU+aciKv7YRmiL3
l8cuv+Pp0iDBkowA1neV0fTNAoJ09VtgoSx6Eoh36yGrlPaMQu92suiw3GM3db7gOAv+qs7M/+cp
PVKzS4cKhqQmuIcjA3yRl4iJ2h96syCysZnYV4NWCoberLdj/QV1UBmNonsJSKhRD/jZrA45Z/fi
uSQbJcqVCOu1CcYPrMYlJBs/4M1Y4r+2ObWw4d4y4oV7rezgeIVUCIgnRnsTQzrikC+K1UVQ5QWo
APKZNW+Gw0ruOn2Urt8izvoaa/v9xUm8Nc7sE75WRe58/HpXY+nXozXHeqJJ9tRiA2oU+A427pg1
2jjOtJM8fEvk7OxLFjBj5jLAjLxrTS3NTTP51toqEKh1a6I41ljjDAMQ3mI/bUvCmko6xF8SR+b0
0FnXF53uxbrNCRudja4XAurOC9ZU6EAq3l8MQy3qZMNoNg0Zjnr347sWHfe5T/Vn6qAMm79lTJ9D
Wex+n5eb7MifqiEL/JBCQ2piP9/CxKTt6VkaB+gIhpdvrmodQh1O3H2Nnxhl9pizH1/q89IwyU20
lX0Iac4qocTkOhVenXFDVwoICoqoB51l5dopz5cS0/c01nrGTA23la07D47tIIWNoB+XRfOJ3uU5
0+mQ6+NbcbgzTeQrc67r7Kv5GRmO4ydMghVcq6YZjNEnJGwK363XR7dkB3kN3GG+fsr0rmRWNM5A
8KjYSAjj8Dhu7J3+eBBlQn2Ex/kLcoRHD/VVf5B5xv+kl05TdUGCa42ZbSjo0z8+Uw/t45EyE3PC
LmBfdDs/laC2Biiaoz1laaox5Ffed/tSp/bXBQssXF5xrjCVXxsrruTzhZTygmc63PFSn6hGnfoj
vbvelHuhusXiZFR63YW6vU2UVeM0nFJjCWxAnyUEthQUVB0nBUBwiYwg57Dgj+UevYxq/XMcMISA
DAhLTmYS2Y5d295v7gw+Z+aeuHrOmhKwD5Xjg1EuBE+g/xMHRjCRUrejMhfdR/ff5HthgAXtd/eU
Az2dfedXVNZ2ax01zySefZSw0r1yxf/p+rJvXdYfTQeV8Yqr8rQNTAJB1rFfQ23nDGiJUKqwvb/g
J0l00lHRxLd0p7/dHWk0a9A7nStXDqIENH/9PlAmWQoYflTQZe83g8y90GUuQGWJBzoaQ85EBsxf
j0yBEDjPJKACZ0XhMi+ygoWb/aQQqHtOMXzKSOk1/aRv22jCY8Yu7Urn6shf8T5dFYKj1JJerZxd
chzrP73ZfTrxtDwurov1tTEkb6JGmRxizyEa3qvvg8feDodtCEIICLztzdOYKLR2sz+klNEBNPy5
S+wMZdYWQSQ61sQmSJE9jlNO8QPj8cZRzCgh+rnLmhxGOkJ5xMIwM0gpEaD9Ty+qdTlbbUOLXy4F
tq1B4y7flVWtyAL1MLrPYsKCdXbP9dTip3PRDSy/h/yakOWj/zZjz0vQ+ZqYHguSpIa3s+9WmnBC
mJedKLEHnV3cq4c1HYXURjZf0HSgeohdcu9bRKdwuaaP1AnuOZPCzXvZ6Xq+T9GjzuwELJ6nhoke
WTmizP2KYPGiIJ1GpFuQ5Kbt5m2sq2wIWyLSXHc2Tq6JV7mIDIgNUSn88fHC3uuzwv3ntxPXONGW
+24bqTkVq2/Oz89J7/fDvvnOT6DaevGaWTG9vGUO0ZNzpeJCRrXSsFCJs+zv06iyemBXCNwlOQuj
El/5MjdFACNpmA+5C9Vmp7XtWaAucfpBcriszSgAB/4UVzWQISbUz/bt4CX+1FJX8O39dKZQ2WST
Axs1yf6CsY+uLwoF1HWASNddkB6yLkG1yiVz+mDlDxZW89Kh5NPVry+LVXCGTIM6ZOKgQOOMT0tF
88Y3d/ud5ZHHWll/zkYIF1sKyEOJuNehlfZeNS1JWughXm7mLFJ/bSCL7G0EgHlyLAvGqheajkjv
uhd6LLW0o+HAZ+fXZ2Utkugs+4fNrqKjFQ2Xqe8Grk3taedpoRRXOQH53e/adG9SwFLzSzHZp9Dy
4of9EuT7P4y+os2MCtHuIAPB66CXqkbW58tBveAhr44PETltuycTrPeoXCbAQ98OvwDrSA7zEybd
REs/sjBwwIAq5S3O07emJ5DL5BVCyP/d+rMhMLPPRVgbi9MJ6iDMd2YzDi2IQ3Rcmc5E6VusuOg5
ZkANtjN2BgQHzJt2X7E6FC/nO9D5Kw47f5rHQg1M9ppKRYa6TU/GF+x3LJQCQ9Pd1GQIyzUyC0MR
NVi6QR7osNWkHI3bsVtUDaJqhdJVQnEA9s077dHKKrAVvvr+6MOBH1EW46xkRbG/I/V1RnpLtNJj
kLX/uOd6Ksk97nI4ObSHWlGMrPIychFmEuJc53cCJydpegANkUb9u5gW8zHostLnjwCZZuVGq+Vn
U9JAHrKcNO7B3PNy+kEUBIFI/SsBWd+VZyUx2dvom0CcqzWVmRHYj66c1Fce6+e4bresDbHLhD0z
jgzmMdz1UQbycrjiq5FM025umWPlS6l9FTMwK8TVK8enOQ10XWDIfzACkIqFE2i1qEiBda1Tr8PE
bg9Gb/Bs2+emjUcjZlcEEHL8i2PjrbjiDF3x/H7TnefqA/a5U+EI73SvdaV2q6pK4QLuj4h0FVCU
ul2y+zEu9Ob0RSoN3mJtqzklpEBuycWnCxcE7SclzUkwObzae7VMw5HR0R+2lCDdIpP3u5lCPBvx
+T9N4048PSBk1OdPNiG8fUk36qmt+3uJHz7I1LQWg4272e8fQX/Vz4Hc/VBKbUpgt6DmX7ISKrwb
iGhbKMzPrM/SqfBE0nh8cMg03JVEyIf1XVYSUeUYRNtADD08CBj5d/Iqvqd4+WmlgIdHUlgXa4TY
GUYAdx037MQNaYJm6DznYOPuWCzH9vfgk924IFy///Ly6ivtOth5SAdVEJTPxpebVNLc/RrRCrBK
CeoUAA8+lOcQRudZ+l9P8TAYYQGZHHB8NBOAjRPo4k4UCTKh1ltiFr/QaDQ9N3qPlTuMgivBycA+
YYh1lwAb6+LMj/YeL/3ASnad1fLG5De7tWvUiOrlMfnyDTNQdz//QTTgD+t0zpseb1Vnc+zdkqbD
9YkWRsyXwIFLGChj9qPj2/pOa+XAUyIKyb99npwBscH+PSCg+4O+G3aX5MQPOGSzw24FeRbtFTIV
+7k+fhJ2tcp/n8JMEmt7TTyHX8mTsCi9t9Lf1LDRCbmjZewj6NDps+8aYcNNwdLzACQHVNGqt3UH
1P0csU6c9UaHETAHZyRP14AGq2EwQcmCCv7iYuFxp2Z992ogDvGIcLXY+IQTkp1AFpv79cPMUhr2
tWvi1S7FPBl4cNFp+IcRFN60xprBlmlQA7CiBx7a+aD1IQUGRhJ+CdHz0zQwkVcp1fj3nnJJFPI7
2QkSzNSYqJ80KxOT29UARm+WljiZ9EbB6h7Fbsuu9BcWC+i22RAJpFfi4SAIyd7RqqVVmcC46uOc
O1yFaY9TTu+bFtijwXwo79s/Tamt93YmZAuJpHjPTEtd8pC7zHY086cv4HzXTf4XSkAi0chhOTbX
x04fEhBK+T46+Vel9SYEuxcvkNFDstt1BLWAgiqxZsGHkhbe9Z4w7rK3r9TWwtXYhoKJaX0S9xDf
VHZ9N9c9czryXkvgq+qxcBWmA7EuqGkwRef5hbzkb/xuOAqcOwcI/zsyiRg4en56ZX6gXNu8Zy+I
VXOxGsnvPbakLEpySNLckt4Dz6+41iOXJR7WhOKqGUC7QVq1I/6ceXpFTzwAm4mxChqk9bUvEfFR
0Ab3GBpVZ+3LfnnGfHS8bWsdvzhg11BrFnityrdpfQCIB1QT00a7l63MfhLbBzApiVSF9gRstV7j
lKF07mQlHfVztwr3tlK6qqpnKlwA04MU0iIqsvf229QXASckMFn5ldVH3rFk//NdxZsWs/K/lK5O
MB0a4QIRC8yjwXzfC/FHQwNUzCpcbTYRc/ARFWhN9uTfH98+7v9MQlCC9fcECF1HQF/gJes5lnq1
0LbDc56JV6PylFGjV3pIZMRMFp7kRUc9FKTv2axAOpsABVbYDR0xqwDXewBmXMKqPqSHoRLo2dnK
1PViBnJojFa/Z8s6kV2LKEXZY7+en2g3RA6SFciEDbVsfAIzmVRHB3gXy5nuSkd2AXLpVq1fyKUS
k4nlKD8fv+oyx+JNX5YY3hapM7yY7ZngHR1mU2x6UoO79zP/pnTya2tg6SVpH5DKBS3Zuzz8Q9RB
fQxlqlYvX7MiARWXkBNKxpqAGSndFMS/A+V2VOMma9YFMcQm6luo8+AhPDNUUChKgS07kbZCQ51m
pZEOG8gtGGx4Ul2/nDBs2Ev6T6oUhd7Kd6DCzdgFX2Kjj0etOXmomSfo4xn9S9Eyji2Cycu+wDZZ
EPFF2IxRkPTdi4+qX/UnRb6AKIyhEc43okfcIlUx/br3CQwwHcXHfknFQvtT9wqT6JPWMgVigrWD
4NEV22D+kfO2z0wopcTxZ7dCwwAkf3bwlCjIbg1nhgVdXRWQ37XViL1s7rxbQ0j96dVrQhBu7Mjy
oiWzL0mK8QBTb/a+f6TahWRcml3wrJrui5ZYmlG/gcEk5cVOyvIz7xQbGVniLHqbCuYikhkTnjo3
EK6KZ3pMPXYWmUSyXcctsubOwd4q6OIs6vDxPC1FKj8wGhyXv2F2HbE/PiFZo8I609P4PwcpQNMZ
+E3NZSggwmixkeIstLqFMitwjG+2+m7gaeBxhDNTpO4gQ03Zj1iCmSbYxs3pRo78Qd/qWHCoqWLe
rzBZKxXaL2VEnWAaMUO3G/wEy0Zcd592kWH4pzIxVuvHc2oPw7OiPq64cj9pJAaV6ZbGg+n2vf0T
zoHvauBoJv78bupvZb8W8SIW2VkOyuyYPkr4fP6OEY2Rl0SnlH4B0DTNntmYHqwhc4pBl+FQ3JLS
6540897cXlTwtklZcghuFqM0PabWZ3H3PxskeV8nxaNh+jYZ9LOvegK/mKBjDscguNlomTYBc4Mq
gXLUjb7nNNQrAQ0AV77JA5VQZH9HmSacsSWNeWp2Q4iMOGQ0LU3Qluig2Yu4MH9Fv1YAcT8/50Gv
2yj2S/MADpXyvq6R0fIhGiq+xKEDF94Z5UckJPmdj2rlx5PNiUjg3D7rilf7DAFf1oxS4wuN1JxZ
khFL0fKTdNlzCOJmBQVW2syLLLvuAgK+iQiJ/6W7dM24iX31PcsPLdRPst4Tnh6VykX6UpMLfMBD
QChwch2n0wkPCk2CvwQ+jh0vHPU6DSTz1d/rnMKs1wnazzGmcklzRatTkUlGQPiIRM5chlyByizu
K0+q3Kd7Pj8xdeUvxA+WL+5O7tgBbgmjnR+7NisznTs6+AEULuDkE5sNtMpsCdzYpgHtKX7Ovf/l
suKAIj9jd5N9nwifmCRO1gI/lL4IFxxO2TmixjdYJMmnZqTSXXKKm5kbvlgRd76E2y2vFtYTfnBQ
btI5wP00I23/zd1U2/KiPZAqLH/l/o4bfFnBTrzWG0G3GyHAr7k92oC3vBpUkc3kbExADtYmbCUr
ccY0/XEolp86bGNLiMtWb8ZmWgXz6tcZabUNiDyclBINeuxH9Okpfx82XdoIDStMQGk5jq+rYySi
Ov0a2ryxsKhOnVMHVO0ksvJMp5N1l5CB9wYWfD32Is5F/N7JDqd+zQ30XXriOnD3VTaHuwqVU703
HCEXCLvxWg8BY2lIQb0IVzH0tHptm+MCU7HyAZ9GAoH10dahuI0h8KcEfKChJfRg8Y7m085GKqaf
Hwgu3gXD8JozM3kluNIef1AzbQAoWMJ7F7B9fFvgwWDRGQna3eJEUQWcHfC3N9hOZGJAW5Fl1mvW
YRjBHqzQJLozVdXFBeNBPmXK+QW4CH7M8mMPAaaAao0fLY/vfUz+pokmJpgrRCk8hM6RPvPH4Q8l
vPWPGRcj9SvDlonO3OJrD9MxL3M1yxzXwvGc4MczPyEMSMQkmqhVoTUsXAtXiuBmXfcPIa3rksMH
wA+SSfzdXep4yDJBVDVBd+Y6LiRCjeBTDjiDhEhCTSChiE2biAEHmdKlSnEzDmICDeLeXACwpehu
K5zIS+SYmY20jZsq1TavHgWGHYRwOoQyvFqfX27GKaULu6V9RlTTuUDnrCeQ9S2EsJlpf3ZSnO2+
dT5tvv2jx7YzIv1Jq3jHA7cvMuyWd9J9sG1jAJD5OikN9teAYsXbTq6Id6mfivuHg+qp+LIvc5DK
yBp2IfrLfpt/5rYRQEMBUfLXSbFfMBzUyO6NOknw1ewhhbDivrQEvEgzH4dXeOxKU8Bqkp7XuTED
foAmTkrLh0gz1SOUaxf3ODKE2PMcp5vJBXpmVxeMjQGMiizw2sUvke+NmMiTXNCFXGxGQexu9azC
pOGG9Of/AsIE5Rd/t6sqllG6c1eLDhYeQSs1dpg082EXIe6QKr27Hko5JdPSBzjlS6XJwqueevjb
GRYf4TW5uBWUhAXAonOUyDHW4NqUBZC27lQpLnxQwVt1vuDMXtNsNGCPBk9w4dJ4cAQaKp4V+Fpl
81o9zh5TqFmhUFlXge4DmMjQO3aq2mygDUb9VZ3DILiOVlCA0xTITRn3ndZZ1jFL/Fx211lhen1/
Qi/Sc7NnGYqKi4o8Qhp+L3xlP2PVW5G1xzqVe6qouS8zJfVZOWYJjWhnjEJsJo+1m/jYKLTrxUFP
TIDO2D+Ai3MNokVBjKaXDuyXrR52ZYaCZSo7XWF++dUnYsb1zDnvfQjyoL9LpVpO5gUMzpVk5UXa
eIDJd4Bu+/1eal/N27yI9Ej9Hiod20jQLrKXYiKuEj1cvUx9V9satoI1L1QgJBIvdir2X3qjEa56
Zix3LNPdKhNfz/WttE5S5OQhDrdgw9oABxhP26vy/22XvMQE4jWfwgVqpaUDycQy2/i6kLYsacJs
iXlAMnFE0OHIRWHJ6q3KDmCmPvWXhqqxtC2FrpTdUvrNG4/4hdyW8RZ3gADuO6M9nWJCDkc7NwXU
lLogyzM+7s8fgTwANQ0KYGSFTTCrOjthe2/mhEAOrRua0JAkdX2tDAG+KmAjI+MyylTUY31aARPN
0ZkwMadd38UpD/V5Zvdsy+mBzfbibjZl+DChHt2yyzmuELRd4dhuied/tbctCQUvBpABSiONHPI4
YAmuQZ3flfjbZGe73CLuyU0UDDQxEjES9I5n59hAGBIuEL9W5MahcnoEN0MJNfVgi8Ou0WwyNHls
4d23rwZelGAUxwDmY8hz8OFfx4heGQTKF6yVspr1cvH6AQ4SPUhYBotnBSGwUoSWp5fT18j/zKh6
sGRv8q+DtmbWrpXNpfgmZeIzkJhHhdWmjFNT/hkfw89x0K0v2M3elDbRJbN9HkzAFBg8QFr3aLg0
q1B47umERYCFKSnBnIL5oJ5876ekTPsS4CWkFwKx/yIK5WbN7/jX6ltEI/bLcqAHKqA1uE+rANtP
y4h1CpbcRc/nnkaXL3rNHKJKFQ1CVH9foaGNPLM35Curicn4r77NPIoYn82gkTu1Ie8IaeJf3tQw
Oa5g/LhFh5ddGsK7SnWh52h4eE/95hHH76aIAvgjm2B+yzD+aTbVm62kagmBuousK5A1FJ5Ratib
R9R3o/xP6J9V7VZLZ8O30mJryYYwAm0IsvIyHiWKu3El+REp2jL23Cy3ryEBZnivTqs7NnT/kUu5
+Fre3PwQTDwGw1ZR9eTIzquS1MDVU1gR5pfhmsh2L3vcihZv8nXai72xvkO1Z6RR3yUOHANjpIYv
B5qGnkiNsVe83DhHtnwjkJyy7fEvzMSHUHRwJGvLMBv1rt+kx5w9ZDSqO6cRS/ohnhojn8qDEIMB
S0+VGk3oVd9iQQ0Yc8WHyLZvZEPwkCLarTT8/+v1u0f8GFKtWuJyLX1yRFSeviV5r1nXjJM4pe/P
ID6bSM67DBwYPzITOqUf4ePVXBPV+Jd70qq7HNDdsbsnvoHfG2Hx9S/CsFm9kXtpjnsHp/3zPq5T
MA8BwJooojoaJJWxx/a2pH52NGwMaQwfnPSdnEBBkpX7rEtHGOsm6By7K6rqvHjx0kQYwSTZ06bL
O1a6umLOkhZokjQoD4ipJvkXLB22eP2KPRwZg99wqfUMxTbE7qU2RdIwOQAzhSraPfhF0fIxz5D5
bTAgqsf9YOQBbkZRuKSHA9PgNtdWPbbmyhyBebf6mXk5zfDgYglLqZDrk/iF8BjYdZODsr73R7fm
F44KN+0H2aDgcDUxQt4Szfxa90+3jK6etYsOgYPvPUrfEPemH/d6ngyGj1Ke5Dy9V4a8uVQDNdnG
Ow5dswVt2BAPNdHJTL5zA18IAguYrM9hhJch3ej5tdOCft62CdLj4mVEho23Hv43RbjJB/EXAcIr
8LpMMxUm4yVZCkVrfTqwg1cUD+NyAtUsNW96TbabotWOIX+n/7WRUtsArdbEF6gw6dt1HSLcHXtS
6Gw4fj/Mm6Rq2IH7fP78zd8QjtchLD/sBaMHjPSL3eAt7xY3DUtUJIkMaJJy2L2IEtgXpDijszk5
QiBWMRbJ9O03DyIqUfZS55BZEYXoDbqDb9YHlzbbTJdJz1aHO/jiMIl3pOuCgE3o5YlwnlJxli6q
tSU0/s7XiaN3s5VCCHqYA89VpArA5C7JHYO5Ds5dIiRUoU1eMJdiQZ6H52Vaf6t7OWPlIuwhFslm
cGDs1zNmtwSB8UrdKQEIiUQiBrKb8JzLUKocCIaGm8entGSqtbmba7maSW49UTC3Lxjw8C6idnRp
FOETfRTSmKRPmSaFKa37jHo6Wf+NaA9qykExS5LGTnfyBu/HVCts6CWXS4Rc5vUuEDGy34KEB/Gj
pAfM8nymtj76o12jeU5Film4kOf61oJiEpalaVznWTcOCZlUexiL+fmMWvbIu5HFeieWfsysQL9X
Oz9mnR9I9S886z6oV/KWqQlVWiu7za4SWTlKGCoq0QAEQZPvjvwvW1cZRpmA2iz6rf59igrsNq/q
7vqOX0K3yft4WCDBfC9aLxJ+MHYdVJZQwd+ubhSdf6WRZQWW78xJd69/WPcznzzqMYrKmIyP/fye
WKNon80DlihAof5hjgVDaW9nM8dwypxz63YhJC+iSFFns2/TyIENp8g6NQ5pDRYOxyOwJTXV7paA
U5CYkKpUu5vyX54SgOoyCAWMPqTGh9kD1jtECEWLl346La0CAWhAl56O3lSrY0PHH60evr1fE4hI
yHNF3bNc3ApnA9KSnlBl9EXEhXWcJdCAEx5Wb65r8rTsF2U0euv80a1KXlaGmPsVBAgC5h2z6GB5
54dVFmzwoiEHIQAILigySE+C7S/+XXxjP2jF8tDhxZxvwNnDPll7bT3I2U+eN/qBk1aIbSj8CEGU
xWCkS4MTjnMH7tqxIA9jw17RoLIM3XMbicJ15M+0nWQoHwKy5OaMUrqyLtgzCJtcZ3t+y7Dv6+Rt
t87WYHL/qNpdyxg6xm1v9LPYdoOKkRfZ32FfypIIvt3OzwxIQDjs88RVnxURO1ymUqwlCQvvA/GL
/jdpVm4yoYCdWL7UpZO1SWW5BCClPWbeZnKNc6f5nioD/1KI6qxsSe+wIZ9NFI8LwGsJ2CprIqPO
s4b5T54cii1IqOIswTUx01S2mmO6qLrq/W5jNRtKbM2TzeNu+oakOb9opur7jm9hqleejxX3U5+c
a7MYheP1N/TeM9lginebIkb91tv3G++Qwfyjt8Y1Qcb/zlneZzNvMAdQe49likH4BSym6Hyq0fpp
L4SoxfBKEzGLlHOUnndmYyzN2Ia/qqsqE1Hlau72xH5p80IHv33lS7DIvZu7ErXMBJSB7GyuQg8G
9cH0fdtPTmbRfm3ADUY3QPSm7xoYjJqBrzx4b5qsMPjzsltSv2oZE1tyteUhfVy2F7ze2bXyjqhV
64SKc6R+nvB1S0ogLjOkUERfN9SV1WTvzwuZSbO2U2cHRVYINTE7jeWQiBPcZgE1Fz0Qt2PJ82Vv
IbZAADXT6kGbV+CnE6mEdbeAAsQzpUwkvQsWF74oYE3VvH9HE77PlLecZvqoZDqaU2+fqlr2u3eG
hPYf3biBH2lkrrPkzHRGNzn+wDKWLIS4yxy72P5wwTYmU9b1EcgTIh7+jC3ctnGVk7fA2pb976Y0
236cFc/ASpLNJ5CBDUgr74jO8C8XV3XGKM9t7L/89I7kxyb7gu6Poaluezirri8QyTcMzaqdtX9q
pMxxDS9KJvwOtv5dLn8qPkdBe87VnujftQ3NJI08gOS6QAi/7YPhdAAPgxTBc03w48I0ynOrJNrs
ikJi+au6xv3S5ureGyLQiPWqa7VYc5Ja2SXEU8P6WrweI73WhTIfzt8ewiFxhFhf6XtKW+radSpl
Idc9Cwxq+4Qj4r4L95seWeP8GwthcYCDmef2e7pakqRu8T2kBvFqEnU91eVVoyAkZ7gWuubMdXrW
0H9T/0CzjRsG5MZnYFzoDX204MBTab8v9Lz08G46RWNAEEpr5JeuqojUGlpFf4fN4W6JLnfRaeEi
ltOlQJHjV6UiGdNAlhDyi83QWnAhCh1Ash9HcVJspxvO+cgLLhHHKoTXH74L6MoE8xWfhdqTUDdL
dSuJiZ2pZJ9foAFBsz1FIBYBJyBOJS3wZXSbp4wRc0hyvxKaWDWaO/ao7LxYgFQ65l2UgaKrGhiT
FPeRRdtLWhucPEHlrhRf5RM4/SdDF8hljKuxIrCL8h7BGP4vZJ0oiTskvre0d/XVUYKUBz0oAI3U
3ueytxQal1kXh+bgMs+dMH5q1x0sXx0PumxqcQxS0wJxJ381Q0r3RhdWcfpbyewRxtLVfFZak1s3
1cFnKLH+N6D/cGZp8VYZI/lMAMtdmSpFE8e8mY0rPEQss+OcGlcih6MJkQzmoV3n92Jtp4nSOZK9
aWjYZqfQ+A2zNElB7AY0j1705b6HCDy8H+nEuhbxKXAPTJE2a29Va///gHcx9iPtDIx8OYugvR0N
wKhEo+2FVs0IY0r+tkFEnwGUbYp8+jWPgdGMf3+kqqlA4RI528gbGUpH2dz7abmsGSzgVTetuINl
Qa8Vln1zoZDPSs0LxHzufpNm6I22ifElhUGPYURIwCSDRHfmBxUG38+bzLx/02GL4mEaWh1O+DuD
2zzflcie4sf7vxZwzGcLf/ZqPa1vRtQaAHKh9vOm4mF7qcwbqwBETypGPfN+TRyXT8KEkJ5es6JK
Mx85iUEjdTEuJ0C4JnVQZXHqIA69XzEiMcuui2JCM3pGFA0RdKt3s3vQ9/ZPsxNigEJkHKwMIj+q
CYq8OosoD+v96UKLr5Dxgyh69uQdX7JC5iOGh0v4455p+HVahA2/4W2LxoEHJjqnJaGmw0aEc0K2
Gh/U1GVpXF6KnHqVU/rptQ5WmvwJ+SM1gdpP7F9fXpnxqo+pcHc4TX3at51vIvkusdwfr2IUAs0S
M7l9yiypMmDQ620tAvmav/vjaTxO8byswFx0cnnmBnqEojM2yIuSEbz8Frfg01X1LzMjd1CKSOSO
8VF7t8I+b2do1wcQnBAOonzpygGw4nkxq0gofjJjg/QYhnNYVz63LtD1SW1rs7vncsU07XqQnTRG
bUMMkRt0NF/cFcNc97BD/7DfXRs/aUcWd13Ido3nZbt3y+bP6MsJzYi8DxzMNPPuD6cuoNVECUSM
zOmyIRys8kfv75BXsl/DtbWaBJOMfkXew6xwmHwb33sNCd72FxcKUUmOiHXNqnDrVzsJLRssm0Ms
DKhUwH20mzIwX53oHDc1D74dthZRlUUmW2RdLh/PY1wso4/CaTIRXvapGw+0aPYF5be6JrrzgnM5
/eREaQvZiMi9kmKvoAqG8SQIsLkrqnY+EB/26fVYUVa/ztqK2Ae7VidbUOAPWXyBM8sSWB/FXuso
e+zTiX4yYboVpyW7ugQIQGmW4M3V5pRgZPWKa10EJNeVzPh+dVIoQqB34G9MNAMzT91oCpybn2Oh
mLZLvMPfBPVVgS+Lz38/r0Dh5xcyp+lOqYFM+uzGvvilm2EWxmtr9dO6vJoZH2FuA9ncp9wlYEFB
ZFPJIcAkNkFFpHNEMYKM+F0odKRBX/g1OBiD8skaOFRhvj0D0hhmuaxCB1zIT+7d+D5mYatL8E06
zg8RaQcozJYH48HAXPaoJXiR3h9Gghz9niGshyYkexnXu/NXXqLHko0tQX/1bpbglgKOtWNMxDxW
5XHzXFWjULDdLjP569i0xpoPQfMGefIdtRRwmi+AOmRmHGUVuoBff9Ew1j941aQvyexNIexKREEU
BE8/8QECRHb6PS3nC26zgccIYvBN2Yf1r+OVbXg4bpfuM7nYAA9UyNKfdYt8fYpSZ6c8WmjfPBas
paTdF18r63fBN66zq42N+tohc0qYp5c4qlnUe2FNM6GuaKutxDUPbiaOKvWgwm2OlHRsMbejGQiz
1HIWp5ZGDE7J6M32nkIzA6vqEJzVjW5oyVXgScNwQR14KdePy0s7NEUl0lCImakv5CNKDmTgym5t
m3ne5ywdXGQaVSbm9f8OGyrb2qq3MQqwwqA+1iAvtxH7zACPppjL8eKRwHiwJ4wrodV2Nsm/VeJR
/dslNvdImtYYzJ64qPTQnnrSm0OXcY0h8jmMQUU7NbLZ44aOJG/4mV3OceE8AzQS0dmQLEdURLoC
vhrw31VcqMQppzzqEeMCUCVfkhhlnUIT9cG6m/zHp2THY65Mn7CDnXazdmNoBh/oDS1LM9e2+opF
Hw+7wQwt4SmcXNVZdA6tuK5BSRIubn8sE6ALalH65+Ohfk49H3v2cFI+953LlkAGRMhXsnRS05nH
mSMVfcPsAcxAX536Y2E7owcbPMylpLqzTt+7EydyXnNid0jdUFhWdKIzbYtowgkTkNYYui7gUK79
qi3EmEphwA2V7T+GzjXddOIFNKLEomvQeBD9sM1jUAJcwqO1e2NWBN7XuGkjM9IKpbtbU/OvCTKa
cQKsUt7vuUhGr3AbV9YNMIi+BZ6Gqwxez3nHfxU8ZWi6/DliL/y8nyOpuk8V/AShwB9Xm9kK44oA
xsIOnybzHusP2D0KJG0KcHwenI6QRFt3+d5Hj5hR4OfAFSgIUEwwWq23YJrDH9zIq4oKwSner6CV
zYEXJtinmgfDAqMnHqt3bHtexGPPTjdr2Vho3BTatewqf8hVg+ru1QDWUi04HlwKeE1SgH+nXiLw
Dj3zQfoiflMZSEzxvDdGQRFg52UwWxoeBNYPsXH0Cij88rtqxUX54Nx56oijGtl3jaq6zUj6DJG0
DA/UvjOAtYyghOeo/dXpakNloRqin0dXmUidGj0lA9iZ1SeHM0+cr3/d+8ddW0uPEJNz9OoYhowH
9fU4no9cg7pfBDjS/DQX9gcrpMYNY8oxZx5P5JEudFwTkMQZCkeQuG6XUuO1/WZZXQ+DiuLJcS+e
D2G0TGWFeQONgpUYArpt+KeM/skx+YwVVHEuQCJvBrWEByoVTvH4Gin6dFD/q+q+YbEdpRVhNyNS
TsQaedvrUMnRcJFu/5Bl3Rm4lB2GL7tUmxztOje7vsvAADY7q8HfTP8EyNGNrq0xL9iQDh6dxpqm
SI3Z26xb58UTyiyt/QcIu7P9QN+E5Boxo9Hak+S3w+f34lAhkcj/xvi8NATD5iUd8kQdlSKzFBnA
CTygHZ63XP3v4fo9s5Igo+h9vs7PqncGbGDm0M9Xko7ClIn4fPBiJV4JIrbVQ3MBbk/dj4wo5X8T
oLpIIejYlzmPZmmxtuVmHQx2Gpo4TuFC8VlAAMv6k9gas6Vw37IlOkrVz6lSJVZtfFvpUp1Yphb7
L+HpWorHYJs7yxGWt30UBE/r5hc3pvona8+6vhQOqa+yarrW46ISkvFlC2oGAmi8xxkVfTtsXlGe
N3jvr2A4GcSr5g90HOARfcqko/H7xSDli3GWiKjjTehOKh/WzogFwTsUSjSMzFe7lyDaXJCbDBjP
P/e+guzO3FKRv13IkIKC8WgUpKLz+Kiz4BWwl6Y7d8Zd2dVd+ZMIv0l/ZWO/9KWkUkjWd5UJqlT5
cwre6c3vgJydaiEKIp0IpANkYi2YVI7dbg4ScGmu0Jis+I9VQZpZ23EQme2E+RAKUIw/LQ+pZMep
BOralF5yFycgQoyyIg3uRmLKolnbOVHdAnpdfAyBpMhbhIdC6wIcLyWszuSzM7tJLHTobiGNyPAx
UUOFtaspTqTKybk/8l8vsy+2TrP7oeRSnUgeHfDO/rzDPwiQac+D/l7PKKzk4zgMAXqchL7A4Z5b
0hFndXqF/wJ+hlRi8vgWcJXA4tcW7KJUbr0JlJz+OIN7OTIt7KFNyY/9vMiN+FY6WSsUO3/s/3tP
1kGGq/QbxRSFfY6vLy49WLp22dPocXMf+bwSP9Fi70pJ8AdNb60pYkOyieC//laGWkv134Upn6yr
EgZ8J8k9QGjib2jWZ60huts2GRbcu18nkMLqMG0nql0TPrkoE2LwlDFkZgIdxF7ALFByXATecC23
b4ZeL+Ckshj748EV2h0TDK41ZwW3htd8ysAaLro5DQjl3SgKNIan/r2b1L8cJcaifMb8q/1Kj0/h
Z/zn4EeEToj2s79etp8BytBCwnVaWc6sUgb85rjoRXGgYlH+ZmRIuHV7DkFM9cBDk9++87xrIfeT
Bz3B/9gyblblAj3o3fGrGnPWumSbk9Vao/iwWlRebpORDWIPtyO94NayW2/i1qVFxqketP6V3YGg
7p8IEboe50Q7SI0n6e12H3ywW0WYjik/ukiUAEaQmVp7yxGBu8kbz9keqi+0o0+mIkezQ42GSGCZ
IadluptkwipPgNNYKBoj6FNv5Bcwzh84sftzijPONbHpJbKbP+sGgO8CNRK3s+nM1dIpqTokHLGh
wm8HsvSz5Z9WQ7JdZaA0mv9Uui24lOFp7mxENeLyTr+EUVtEK8Za1dUE7hayUa3s8Yo5eS3hdSuL
Sh8w8TCOAfPWmbNFirnhxuPNUZrXlS3EDth6nPaSe3Xak1OrSxafu0/IdM2Ym5XIOvTjMSenrOQo
35IM27iRFC/NeyrYB162rQ8KWZN/DFHH0r3mKj/qztkLKjvAGXgVNljVW76R80AnaY81lI3EnoCl
LvckT+DBi6aoOAmQMeailT7xPKmt2fN1FT88EM7Vp5YEB3wVkytBD7D/QorqfaQzLR8j0iVjTidF
u/3r4AegXLbw0n+Kzft+2qoiSCxhLwHieZa0Ofmlqy8t+juMVgNjPMeQhqL3ckgZ9qfXU5jnS1BR
E1Z8OeZ9RHWidpVuWeQPhUsi1toL02qfJLmedCUS02CYgW5wQcSKez6XMz+gnoDO7ea0RQvpHayJ
ryREoaMleyzQoeCmKrSvHoVg/VayI548YxtsdVY6BizdEYusprJXMbSO/WtyER50FaRI9UClvEZS
Q5NSywjVDUQOHVYZRGTQDe2YrJMczgE9kbvfQ+JwxDAB1iWdRCrOFNthrRQe8Tvn09xudFPh3CzN
eWFO/iAYwKbNG2TFuTDEaS6KrRZ0b12JBw3iYAXoSobqQGJAvrV0MMSZhUU6Hl093at60KJg7bta
tx46eEqIyvmK0o7fH0e7UhIFBtyriOS2A2iN0JXR3KJLHyjLDZybtB72mrHNProZaekvqbayPySm
L7x2zg1Cf6aJjx38gpPrVOcqvbSXKE+/oY6OuaH+p/vtkf++sCH1gIkJnSrdcbBjepwwmv7scm71
N/IW9V6R6ZvBVEcGlp0Ir/uOLM845SSgOWCGgZi1sAxeviKzFSeFdujR55HIfNh9EZq+KuT+HhCQ
LaDE8r2RYjkhFqPsuM0PTxFKoqSbEGPoKjwL2vpT6p250hIlCuJAn9ybr8MqjwM92I+Tx0DnHBmQ
IDBPD8yXqYWSU2Y1GI9uxoyF+5ek7/SZ+bI329BC8z/AZqQJhVzEXRMOZBLuRwicYY82MtvFHqT1
QmgDL5wbntRHaQcxuWWTTMlc3kMd9FzvGx76+7Z/SeWXSPdxtxYkwuftGyFmKKbu+amr/02wTee8
fW4uNP5heyi3YKCuV6AHqCF7eo1QCdr5zxXIYFnfU2326wVYo82Ah5VlZnNcRTL5Sj7udvuiEXf9
6scYOORF9s8ezovomNRUEtcag1eXUKkCgpg+dvedIkkmpPS5O6XAyPcCfCfm3/c9prkwioGF5ZeG
3oTwipRGWieBeG351vh/zyr5obOUqZ0xX+iaZSunCmLzVkE5mafYWRsKv6uqweioQQPsybrVtA5a
ziLccxIw4UCPvD48H3uqdoEoAEEBcGMwqnxKJf8GQo6whEt2TgCh99kR8i60H6tIaf0la6piuH4Y
XaxLFeKWZtPayHl+DjWVdn6OuXrjEGRqZwUuWzgJP3Pq2/SF7slK0UlONiULCMoBtj6Gnng4F5QQ
+gEWIyGyOMUSTs70+HmPJBFwSX0MzcKNeBtEZBSeLNTDDmC3hIVYak8+CHCU56sfdI2fA6g9EXg0
x9AeTpYMC9FJpqNQl6f4K7fUxqHb577XPJBnH3NkMs5doqjXOGDv4qGRclerjGgoaHU5d4CyULDE
bIhuKsaPE5JGRWpM0G96MxH9o0nuteW0AVbfh4Q0p/Bb1bqlDIP1KQ19JcYIdrqpdWjoP9jCMWkb
4GRj5qGWq/44Q0SHTpAffR5NMgqG5GdgGB+th9idgTTO2msu86Jey0HHRtOEzY6H3g1GHm0iOmU1
kU4Zzzmj5/dcbRdBrdp3tGGacbNDdmN0zt1QTVhqdpPQffO+/onb8VCNjWdXsznN7L0SY+gdeoQv
palaTBI8ub3DCeYMGghFpaMDlsv65tWPKRsfRsk063tHKbcGGEH1h+fsXQeu/tK+QrSjsk7kx6/4
gV1IXbDfF9eo9ibGgMgauRFniV5yu8xPmUleytVHwxrmN37J0fqPbdiz3M0rOvC8wAKqW4uv2HO2
zCSo4UVe9hU2hcwOD1/EpEJXTI/wKUvlb/SfimElMZuwRPPy+IpN+L/4DupxLEktaxe389exXCTK
bkPXtDzkeIi64JEFULQXtAt+7m7eewilZBnh8F0Sxz1zK+CvSd/N0kMV65dhU/CLIS23ePtdbZZ/
mN+DIZarFgD8+IkReWTCKNi9DCi3YhiajMse/6CrQ1wRZDirGjVPlhdQHsudhA6s6hnLLJcpJF6I
BU1MyGWpcQJ/iyjP4PHL1HE04u+/lIjA4SkwfP6IRxb8aAdIjKnsM4Wvvmq6bkdXDvPedAMEWYY1
UYNXKD1Tcan0Sa02wte5wTO1OqlNN7NnwWI2eFg38FvFkWRWVoB2i+f6N3nD7STkzhNN5E6e51r0
KFW3XjurBmoWSPelpg+C62HL1AL0xdDo8z2vFTfLsdvpS0lrQ6jJONAh4+FQWtz2lT0AclbBjpFr
dAQuTiMYd8vEq9zLR/rfUl+LqN/y+Mbw3vjZXISZeDfPh4iTPmjrQMtIKbSNpzeWKo5T6u59AyOX
dFv6prlTSLw9MyEcTRIPuWzy8xw/JW+WfI2STAArrIfKdsCmFT94jnIyYyYqn1o0l8FP0vxQiPqW
Frn/U6Gi+CKCvm2Qe6qhRlfITyAL3Q/yr6jE1QunWoccjdaLICLpfyVPiLuymAdVic2wn3TeQ15e
N/oaKc7nZCYmTUr8Oo5I2BIxJtuquvJHAH8BmtXPj83dJ2aYlGq/D9yTgXSnQesNzbBJ/WPGN7f5
GZOf6aiNE2Cmu/+gwaWQJ0iDQs8yTSAxq9XSomwN+vtOVzD1xZydghl95xgNPEjeWeSQnE8OEI3l
WO/Dt81ROQ++5NgjLoO4w25HWXyDAfyfFd5Wh8YcjMOKWKKAnq3ibXudIa7iZ/RmEi0K+PDuDP1e
gOCbMMchJFZb2BuOBv1rkX8D+W4ubyu4LJMSrqOgjkq+26RRt0rUfxMf+9xtXDl4uTvpVAdd3Lz3
+ShWa5SroIk/bq6h1kE43qZ6jsvXpUST9ASiIk9lMsQHSmBm0Bz3XFdicRWcpPAMTwOOLq5MvU3W
fD5jI2Q6SJdAQHrFqwmoru+bW3no01BMY4eQDlh21kLrXlmYZYXfbJ2RRxzYV57EIPVkzs2lX3tG
lpO/TvmHz7rZvs47YRb2++aH9ITBJrTA+5O4lkAFaC43zYDV2Pnd/xvCjRk73eyluq1rl7pHxsNJ
aDHBFumPsCA7zhS8RkO72h8i5zVKSDzxMUGsolKlz29dIG58d5N07bG8dEQFJqWzfruRLu1qf6Gg
//zryQrTSUA4t4zijVQZJfAuO9qg7TgRobVGgUaV3vSIQjI2BLU91sdsPo8wr8PE13MXnepCZ+Jz
Us5QdlwjUazr9SACbcKYGTjpFBmbsxuVQrE7t3nRMwqtXMVk5MMn4spiwUEAAD+YoICGfjc/HDCn
NO1/4ofJbmwCNSlnAFhrQg8QgCMmTOJ2W//UQDNOTwxG35UePWsESi/3qFSGAb35gcFi9pbabYYC
7i01gjpDULKS56hHqQ6dlzgHE5RcV4o/rINNHiUA3WX5163bc1+wn4G1DZ+wCCOqGKIJnOhnYpoD
cX+hOfjWlxZ3t+jfy67pt4l1yVUnDm7xFl1ZKMfTgvwCOUI0CCcHjW1yAfMhWcATZROzvXjlZZTJ
t/GXp1+xXgLSC8q4AD8MN3vQW6Ys8T1X01y3slj4KiajLmnsrGuFufsQkc+ZObWXfNQfpRjr/rp2
wvytos5J+NDBwjGx/3M3LhT1P8SR+DKgIV1CCpRvhl5QcVsXF/aZ12xwmNRO+lXm9yOCWANAPjxX
GAwhiDGjZcOsNF91OZ/wd/8WiaGX8hNDUucYligx4W55cYDuzglTTvUReEBgt0zMH+bkj7h8Ypyb
fzGSLmdQB5lqO97eNJHh0k3MDdSXNWpG4Bhrq03x01+J7ryJnaR1DR3TOPBG2Cc3whLncaZyxRcd
8UTH5loEOasxl+z+fomuqNFsgmicKeIMeuD7Tz0zge3dm9XMA/sN234K8F7bzXpJFRbkMeW1Tpdq
5WucirQycK4KrR54vc3RireTvwYHS1N++RMhbMNCZfV7jngwHUDy/JMM53GlSe3PuxdJAPow4kbX
96Fn3AZY5IoDQAVl3EFWBBuTfb5u8t8VH0n0NYdkjqFdLuZuq8IafGYGxlXj8LIK0sB2nL0VcFMU
EsJg9SlCC5H7hIldqsW3aDFlWwXlxTcctmixj+YqAHMb6Ikq56EXLQY5CTCAVOhrrRbKkNDBZRDa
Fx80Zr9lMiu4o2aReYcV/STF233+5pqUONDyllAmfeys6CHarJnRZ0sBNxG+0rkBSht6pGNPpn0J
etPOXymaZTNucoe8D9srQ7+BV4AHKW0z1iaLp036cCIxh2cFwxNVlPXIx21NYZQlxelH0riYswGw
AorPEskBxFA6jwA/BQhbIj5mkIUQq/oBjnEcLZZ2jwCEIMommv/Vv572riF7MYexvTZ06btnj8m7
CBuwBn4qS+u2wA/8n827dMcNIDZVAIjmiA6rkZNipQ88JbRYFnHVZt4oVw3z+NGn8o0HtQtdJ7gq
TDY9AOK/ZBS3rtZG6pEV+2NJwnFYMxB9TWm8TjZVu+Dv27O4eSFlfoSTZ0zhDvtnywfxS8tJiWm4
G9WL/epE3n6vSuk0EHfC3a57/cHi1MCHOWgRngxXmYy4wNs+cVQ5VGlpRdMlE4jIeJnhytJ26PlX
p0/XcaxJXyXfRHoZfhAFWm/MbOtsSFQXP/U0KUVOhUeGpiTNj4KdOECV8OoGF6OC5g3UQmN/WQoz
JB2p/JLhdKW8jKqh1VPjoZEu1spZiSTCtyWvL2FHo9eCuflek1uZaJlfZJ6KagG7pQspuTo/QUBh
K8VlpBXA+bZnoYfSDdL3PcNmSkB9jrc9/d9AIpjqXpHXUFNKX66ESJQxCrGuCUO+bpJcxyg84THY
qk2Xgv38Iw2D93PqW5xvUSY3pfUvDa8TfeDi5hqPbGEdKBVBaY+9U0lFM/+duEwpQloTZFAVFZlg
VjwtDJk/7WzgiJq0QPTO673+YjuNJzbtpljWujXU9uT3p14z1VTtp/A7jvE9GZCTq9HdBrarAtwq
bRWNwCuRxt+MLo3mexV2KTA2sZHW8ivbarIvXQ1N/Tcizo+pxaQCOHubbeqOXyDsrR2NefQd/m5F
QAZN/LijR0ENjBxZCA4cmJjYxBtrUvP3i6Gc9+zxkyrh8sjldnipQuprysxKhXPlJHml+vSgp9jJ
dkOVAxtQCcywDoj3vt6KPiqPd9XVxh+JFxFW0XiNzL09jJ3LzLyO+YmVYveUUdpwEnLNtugpivcZ
mHkPc39pQT/Gf1MAy1x9QgckwAtp307lTssTxRi+oNhNiYOSlmiLZcCOxp5Ksk+08W0xCX+cnIIS
u65X+GF6bW69pOGBmgsBbDrmVIWegxn7QeODecj3T1ZMnjzDp0NbaloCUUyM8uhAA8X+j6+rQFq/
YCOvDEBxtWaIZz0QShnTK7cSHmVxZ7sAX6mAicLx4l6S0Bf0PZzDdIPRWxxuCEBbtgYIb905Ax4l
WWi5r84Xe6y+FpIsn3yKb7JKNufLTS6I0+vhB0uQbYJU31sVSqWZ8RWWuhDuxxrphoxC5ciJC+ca
8ShBwjfcbnlDXX9NruKySdbuYWZLQt0UlCJkxrJRY2mC8s9Q3MR9TU2BNZskZ55kqdT50l+Bkovd
SDlWus1VkjyJOH+YSU1kXB2HnSatIEMBm8LbUto7fTo1jyP5TLUJchmwDhurM/BCl7gjge3xAbNV
ZcXrjxTV+74z3xfBgKqL5sUcp7AkKjozLFw+cPVpaYZKLdSAzaNcLNspwJiXC8MfEuuom7yv3vtG
OkZ8x4vUoXJREUuowwkVedHynRMVLk5Mi6cu6f3FX9YfV40p3TiTSpGyr2cY986mk9Jv+FNDH2nx
k8pEfUpMZmdchCH97EhLOQromqsqbkzKlsiYtk4zEgbOQlL+XJtQiC1d8/iUhZSlE+GWqeP6Rb5g
o0q+yGr8DCuLQT3xBFvFe+ghiy+JOZpS/0wn7f5t+pTYg960yqOnMUw976QiJd9EpaRjxF0+pVGz
2pkB5saZ4lcp0WMqhrmr2OeI7K7k52hrMC5Ul6+4zto05VL5Q4rX+okb6vDTetbrFwhTU7iyujU/
VL2SK7nFgjDmD5cneywffDskU7F6DoowZyBqL5BwLx8VjygKw5hrVVIJsjgNlSUlIiRp0O42An2I
Ho3fsRQHbxL/N9BPA4VMLaAYUM4Z6CS90Bj/6WcjEsxcIWWIeqV/g9V7V0n5XnfVGNhK6e6EvnJB
obw/j56ibAEZ9LzJWMJ0GK/Q9LQXYOll20iqUyuaB2SfqKVwZ3HoDaDjUY1sxoIyoGTyzI7cwlC0
D6xrDFTQAsVqnGhdKxBS5s0ClO/jYGb3pAAsimtj1d9iFESiIgUNe998sVD9o5AN9u9sA3v4IGA6
SlVMwoSflBtXk+S0Mk9+/7LJHmOFmyJ3/tZVD6LmdJS+GE1nld9YOEJhUNzNLWU9IVKVymf7Cd8j
uzQizQ4TgA7b8rtVkZNIR8j2HJyLYoE0IvRpQA==
`protect end_protected

