

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qYLayuf0llXi/A/DfBGhhFSQqI33KwMvrOjlYd0A22F/VfYESpSX/xmv4drrYl2j9y2eVvFoIEbm
w+C12h20cw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G5xcUNBVOBJvI3bYH0Q1l8FiIlqECVbgIRFOyyX43yWfkZi9ai4qFPc5/+0WXnzy/yKUU40Iim1l
qxqPZyd2DZhfB2htFiFH9xMbRtXOXb1JT7lBTTghC0m72YJtXDAVPJ12FA7w83KzNjUG8dzya9Fk
VBRc+YskKVCNDiJho5w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WTTsJpSW325QfKSWvk1q/++K3M1JfnanKZhiJEhSizxigYRxOs0IaXjxP3ewb7GNlNusaVp9CBRz
xzdSaiNsaFQX3IDAOB3HLtpfQzTHDCMkx8XPVH6QkJFItqWz0jBPLXx01W3Agqv3N0kCy+fUcROc
qCFeNJOJPRKTmV4DXv7n/+H4YszfJRnRsjR1z/c80hYSYlay+VhV6xvnMpHZTcNYgGVyGjeTr8YB
cDl3FO5by3Xt1S/bGaZB4SDoBl66cT4VvgG1peSKu3FUghvPwAiXhizA7ki2/31bKpQUHJiGVH4r
y+5NdS7saklt9gGLfTKI0RIte99C2OKHKOe6lw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vanaqAo/mjebKVXCqEaCFitV6Elo5iRVywPY06caLUkMADab2uO0QwrboX8k1GTZH8OHcrJUwa8D
UR78UKXVwW+TxBPmnh0GVJTrRkeDJ47AXjJ/rPIo4IEcUMxmBjNbmkgl8k3WOQ7Yw24aeAqNzihv
6csqqIrLhrGNP5nyldQpN1/UML1Px9ZutmwRvVqVL0GP2h/3H69aQLgqhVytvegInxKjoY0niW03
gFcYGHqz/Zmm3QV/VcRJmKnf6tiUgoHR5Wv/HGrCR8NsxA8Ed3NPil0USFzSjuqwlsTQfphjKw3f
uyJdNiXfcJsW/Z1AE3LibE6w9v0hiMFl3j02Dw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YCa2myK7GN99jj9A4RIz71DoBjfkKow/Np70jOI0J9BxSKOft6ILYodUV6TX4JgkjYdKLLrfuV+6
STW4ZONd2bE7aXFzNrEl/GPY897Qq465gHU/LlmVQLEF0eEQUY68ZxxCiGiNLCQGn2Y3E/9ZsEaH
EIjcopI9WR8HOGxwZ52gUGKK6aPIoUE7vGsCbWNXExDKg78oqVOHEbnIIwjDE0E+Fx3rIUyiBMDE
0Kl9UacEaaaJhH4zWFFI5x+5P6v5cfNxU1/y2RQeHtLfTApa6FOwlcNXhP/fmD9nJQVkYi1f6tlS
NoSj+xo4THz3ejxmaAolREJccLOoOxAjKNDtFw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hZf0f+dDQOqIzdgo1glW6ibYdjb29SYxr7QsxxwQzL8GsWZVVPPayGtCk2KwC68TWWCuE06MQsfm
sDTHanO4LO1pW8etZMozf3SoeXHzXK8blBKsBGCm6WGjivqZCYUu+DCd7Q1RGBf29yh8KzO4N2bj
iwgIBhZArtwGXtppDjw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LGqkNhLoWXfqWVssWMOFqy+erktYtdmf7QpigIDucSBm3hRq1NqSdAavcIll7L0qkvZ5QCaPdw+l
/LXgZaom27ZYpQbPQJtZdz/TNtn8cmRtcSDH5aDfyaFTuvLCPWhgNzQ/Ivf6h2GP7zfpPS7x++pg
nkaka+d5PHHqFrXVBhftQ0xig/99oxR0hJTjqBrO8/PiHFlzq28aeW2fXqZ4m+QuC3VbfCgLumMI
lwo4IqHMtVWb/jMrImKKmXaEWzAWnrV7Faul8wBmnvqQzlzcA8kxG6stfWRQooXi0X/zQ2mdJ5LZ
SYOt+fTL0EyXV2+LPbQJ+1RX6PED9rct6FsccA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DGnFxVpxFXUpDo2or+5cWWyyqPvdDEBZyhQF8a4tcvdDKNMEAqxVAPqPKVKI85pvolZxRfD2bHPv
ABcaGrC53gfTjy5nZHbBZRdLOUcZfT943hhHu9dZURt68YcKg43T3zClYLJToT9mv9aHEK3sqtce
mCL6j9a28VaSGEJMfN/jaKqlF6LBMI+HeIPgKZjTO2mmyIF8QTgoLta9evCNnvMaziLhxXDQZpmM
Xo0BiCwvIBMT/vMnFvp1aeVeKkZ0y0ySSSma3/ylVAAqFVKG4Pob80EHQPlwsAwnpAi0RJboiXw+
gqA0ZaQh1fuaxBKzHWYsR3yql6/itkL/uRzgqw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99648)
`protect data_block
MhkkFG6GvE7VttYCct0Wzi8ospqUEg8vhNZWLQhJE3oQJFGP+J5PIUHmz3GYcW/Opz3dmoXT6Ysw
EW9ZVi5lCTruRsWipmqwebU6VSrOXAjw5gTYWbxhvx5Hyxkak5eY+mzD8Njth7SeRybpgd5bN1bv
WQVK4vtRbTR7u8+mgDMdfQQ/6XLiqTIn9pTyvA1HVey6aZ877Nxcsu3Pg63b0nYVMdERK75Dzxj8
SCGdScDGANzRyEhfveTJGF9BZYLWZffrhpnpE1D0LzuHgLITqGmixMUUJz6C4+ayQoZ2+AlThwXQ
oZcKrDWg1/9wPKqafOMIltNQRnleFBIMRr0FkwirO4H3Jq/jaoolxXWzp+0Gg4SBMskVtqrCmhIJ
umdQRWXN4Yk41Qndlzt+wCqVfoejBLZRebOi7kjQBbmxQdyKU1qpixgkeO6BfLnTcVvC9ETtLKbI
ds+wOkgw0qXWd9rPD99wCbuH3+WNnlF6DUh3KxbGuF3yd1PKIaMfMLTkTge5UunNpJ9JkGOOzdSV
79p24Aqr2knkByHWyaONuMQ97jgUyPFZfEuXlb3Wy3Fticedsaq1aJacD3kXsBF2luqVqLveged0
T1sb8u8aymzmyagIegoiq3XYOeSWC1irQEfqkKYqpwr8yTKc6rfQtyCSF//f0+BAeEunQZ+wThzU
zf4q6iMe9yjRDsB1W2nGXzXNJQ6CmeeUuHBoDUJey2G7CemLjhOZ5awmHN9KFs1czoLmyVcp4zJ4
NKcODVMyKkXe+dZDLb1o7CIbNUC+dH9ExyLba9gnayQY87hWR7UOh5iQq/I9GrB6Mxzt0viZqHrb
xSq+ApwPxktdL/+qDYvErWL744QjPLF1yLNccnhYwEV5+mow298yZcGodXiHTnzF5r1TYdfUMGPN
3MOJIj3TawyexBmcbCTRTCmY6fLGx5I4OF0O4xFbR//F1kERCwITL5hz1E84rtorZTOsLn+x+tyT
dhBrzEmt505n25GUgIL9nXH2LqcYNDYCy3g31U+gbKRb2+C2AJrnYAXDpQ45pkQKRZaEGiFYljE4
cW8vr0MkEf+9e0I4tKUL/xpqmTl7WHnL4tDEUrObOTrsmUGM8XCiqFlgHLlZNeh4mySQCRyk1Kyi
28eLSVLkNH7gNHXVsU8BstSsm7FU7o1TZvs3VpRnli64XZfss7nqJ9jLqrIRqJhtEbrM/TPi+Uox
ENV7dxhG2+T7d6NKGmFO4EhCPz+lFd5y7LPuJW400GeOSx7HyGY6SaGr1MQlMUeJUYJsIMJGqMPC
+A157x298TfsukzEQOEjyu2OriO4tZiUfQZlywK31x264brP/uJsENopPqz6UTJOz5a6w1NvFsIz
icBwnM6hpXFjzkMjgjOu5EXU60HoduRWxsCVI0d503cjqicTmxQ0fXNx1W1SxFvswHS5XMvsYDf8
CL1dwgcnmCFgOmHtCUQs+RlQ3+6BIWVsOsXNQK4N2sqVGMuNL/KzwDmGZkTajFGtpGvY3MM/JJwI
MXdQ+N6yHdb/39nWqUkbcUht28DbIKNp8Gfx2abC6YXOcdWysfI6EqlPpz4/AKjzYPd/VRJW7iuh
fEXe/wVn9cQIwL/WmkhaXLyiu2+21kOVp/HmSIZn9LmNuimxNkzXjGhmvnhcb+uLPgLzDbsAu9Bo
oMoVs8zAlTBlwrIdyqcNW6OPg2WMCu/L2uFBI034QkVSFu1nBu5Uf/FbH3TdG1ry9Nc0gRFPvTDC
xaWgH0srH7BHrRoNaUGBaozATqgGayAZMVVenb5QTkoiQFt/LMOBKWSWjLXpwDt9yNk9ily3UWAN
g8iyfuJM/zwaZJgr/dODyYGnvv4GCeiYlsO+AG+25o5A10gW3A4hH9pSFuWo9LwvZGTW+z2/S6ZC
aT6mjvkCZEiP8cc55tx9/2YxKx1K+Obr2m0frd4FJUsQfTanl6EK2IiMk099ZV/mbxfjzFxU5GPt
LZYpzzGGzdQextHgv5qNI3LSQavFqXD2lSia+g/yVUJc+njdueTxujYtoraq26yKG7+G6mRZfW2e
70PyNWNkrZ5DhhDijm3Jn9rLsQtgcvFwfQGO9EdyzdSLsS5Arl9b2iXngnAHLu4I0VImXt2Plhkl
3yj8j4x+Tcf4j9N5Ta/UsonPUGeYS1TjTtGHbmk2MjSC/yGSUzfU1uSsky6anWzoDJ6ybb61EtDa
YmGpNkI+QlAoTtUwSy6A3KmuMYbsgY/Y07eTtprz8w0czr6AGnkUOrLLR8I4Ox8K4K0cnaJPxIJ0
tuq9w+IM6WjxZL8X2j+3vJtXF1R8B8NSanGieqBBQ0x0nbuZG6+MY4PkCbJgNkuxi+GqmoN5PG4M
9TC7Eul176CcCitCSHh/TeScXl0aSLt2rRbMLFXmMEUDsGJfwnSa5AuxJKnUOLrB7vR6NucTBq50
4M8uZKZm8/lKnmj3LU9n/NuJ8MbpqyALjXYTPtMt0Lkx7afbR2K6hrDOeEoHhYz4tmusfIVqDtI8
IJo2YljVUV3LniwnRrvDxZvjlMQoNP2qcZ1UdxcGL9INZvXpjrYMhXVkVV/euRXw/aDjU9q6qBz8
Bi8y4+I+GPN7khpKcAktwMYi1DAunobkSwub53Eb8lBN50nxuWODQKgmXGrQ9zkVvevfpFooNX/a
kiFDHQ2du0c4sZBoyyJCqrzkwyYA3UvlyBRgXtcmTtCSy4sCGpBuIAFIh1TvDDsqdVBFDwKoNAJl
ZHsG7f2TswG5Aq+0q6yYVARxHvZx4pWvzGzjPCmEScXQyED4RE9cHBrQOCAtQscHdmLKuoLt1Yte
oBlrbIht86uJjPyEImJRpHmYPB9PftOcwaj9+kSpku+uNo1/pkN/KoVY2DNy+Lmtf1zwp9kAqiCo
SgTMZVjgtNoMcLEYAI097S9B/sfVdNAC440uAe4nMwp0ipwbYXlT6cQV3Ymkc2dn58AxenXwRV2J
0N5E9a2iXpN3dSAjdDYxJwSo8WqZisXEYvyn7h0wjYVd1ut1fe9nazF8tvkjfFdTTxAXnLAE0T0+
wWbI7u+o/CLTBvkEVeonaDN/BlUIaZMZIaHu/ALZscrzJMg4BhEZBTh0nj/bq7ww0yMgYBRJZVh4
j/Ftyz1+92wygc5rp1DnKkhAFb9j1ZfWmZTbV5Z3ndC5jgeeuUD+aIfMySJs9KtH7ZNq5cV6MuOb
UwriR9kP4BsmICnFivEQRiu/s+9srOiIDq+sNpj13mdspPpe2M7/+Kfj4zsO35o+o9AO3Mp2zb9Q
1o8q4tEs9o1rPA6QcqbF/xI46zBicKCUVIDuZneiKxeu2x0b8negGVI65v7H4+OlVKcmXnA5+03Z
tp8sArxZll+tzF+Oi+cNmIny5zyi0a1Ahf2r+KEw6hXvLsFvG85qVpWepJcQXEYSNAhJG+d/tA6h
9UQTY3y7f/fLxVfDAC1oZAipimBAMksLcDVQcTmubt8jiHx+OZ1szytGzRumIC9yLkbfFGZ0tuy7
QEATzPanQXrvgRKfuUQI4k4lUTggMY3VfPgsgr+cJxzF1JOLBrnVHnkjTQiqhgeqsn4G3zJGVm+F
3f5Klyq3CjEMA0DvwmP9r785hgSR84LnzLcw51Zc2GbmJPKKRVS+sxci9cqZN41g0XD+sNHTz9qW
h4cnbtFOAfxMOacQLT3gAdEvdmzdw1qpZqjcZ0JrvHqSa4O3NoN1wWhcW/1AJf5JTo+kt3HwEBjA
KNELtgatljP+JR/tGygqZmjPYeFV79oZGRzuMltZQzGrPm5wXhzn37LlW+HvjQ4824/VAc6vJf/6
uQBFPRYmI8quB6BJSZJbEnjRA2h3UjKOawAO8UNjHME1450DEvGr9ZOcyyyOpK0DpijSYykgkeye
+MjedSIYRZZX1a0S1CRffXArzuHqrV9RVqTNtMD9yCN9+BanRozp85TG3Ygdw/t91XvyNDlBDOeb
iEY34I2yqiuaFHp1acCIO7fpuhry0L95VhIxglv6CCN8sVJ6TfBMR4By7hTCaZ28yvwL5jksN2up
8ryJGwm+AWwkQ70g9mMPPNaZaMAXR3e9j7DzayQAZbNNyA9jcLrrQMTMB4WnUZ5dU8CV2hIdogQE
B0hkF7aCrMU6xDzXLqmUNfp+eRLBbLgHnBWHh5ikOxE3mikGfEwn8bi7CYL/jKd39dDYJQbHQ3Xa
1eieXaeF1/nn8X53dGeqLIlh21VQ66X+y1VZWhS5HGUL1y9s6ew0gTDaGqVUg9uCF3t+zbH7DvGj
sWqr485HxqAfsx5oyGv9jBPrdWMsIPqsbL2SWx5Vw7sZ4VzqXTLWzxPmJrU2FrB+2AkoT+qtKFgD
SYjt6d9zsOmjTmnkFdMl3sLf1hjLn8F1z+ppxdCrOfv8oV7smbqLJQY++6NudMpNuRQ5DxnNb+Jf
eYxbHhpVDE2ft7/qfAtubt0uJ7TJqP/27T57mefJtD3t4L8W0rP/86MVNr0mwedV54X1xwWbZf8T
YlNSgbaVRiAIExorRW6rSKlVdvz3+irVF/u0tCMf6j0JdDWOZ/jThyBBr9yEG2Z9ZcHl+AxcjFqy
7DfGIlqNExo2ZSM30XEfGujtb+MLA+xPCGRfK53kX9yufoEsh7vf1C4Ui1cQMqa5XwpVjwfCAUby
OmEg/sn3IfmJATVfxZpqsZzvU7dVkh2xuZotdBybmWTutPFYsni9S/4kpknki+tbagO3o7JWWSgi
ptj+cISSGvngj2WIsAICEgaTRf6gTKCfACrOgGPN+/B9miPXtadZehdTIX/sCkcqagWHqfBQIx56
ZI4m08S/aJZ1beWAszQiXneBXFgGVLmkb9yVNsu60+cJ4ZKSQtaUNwb3DJ8OZmYkTbqOHZn2eSsE
pFk0OrA57ND1XgdxyBDdIJLZR93til6uo2f1VhZYlW40pGpSdxSsw0sJgZ0sy02gIEge/lrSyZsq
S5LytleMVdeK2eZgX66iCm9pUVzbmqyflxki2nqOtZMYQJqzE62pqAHv9n9FiPiRE64cZB4dUF5N
nJkvXyCax/JYCcBw9U/1jRdXhoyAgW/xQqkINW6oaCOV32sWU4FJPZ5JdZcAb2rDEtOyLQunJo3h
vcI2o7hX6QmilhV6qrJuDD8+5sXhyD2z2MyqD+8uspExMjAvtqD7Ug9QRaZ16nbRO/6o/R9ZDK2A
cw7UuvxIQLmytZNTJMx3uUz9nvGGstmxLSqj/lra4lkR9nitT0tmiBew7/P9rL72+kui8m2wZTuz
4hDmSLoVJODC56QeR9arzaSNCDWeCjQ9U3xx4Btl9EDyqXyaVbVp6BG7GaBlmivIKjqE0yqISrE7
X5NihWijxLne6qdrUZGBHFwR+lCbqmaYf4U/PF0nC45h95tC4nSH90hq18E2dOrE/KiDq9p+6h2X
wjbiexF9kNOmVjw7SGXlR+nSTFO0LUL88ohUyrXimjNbbWGvDaTBxN9kmRecPXu1SUr2jLrRnwlM
Il3dL6A3gCXYiRbcJFeWcMMTd4OeZO+W/Nr9ni02oedd9coVhvwlHWZ9qy44ovIkF5lX43U/PajE
qRQnMJdJkxUXURv0obfyyrVMY2GqEMoQp66BJaigNsjMJpw3p3bOFqFSf0m/4q+j81eeENglArTV
qJqNiAUaMTABno0K+U9GNFMcrX/YFCMZ2JRspzw7Fmd2We0GC4J/pyJmFUyC3I6h/wgqQIRtO+QZ
1H2dBgTELjl44OIW6QJujfxUUYriWjhBxJXPEWqW+9U3nzb7wxweQjqs2gDQ+cFJ+0XEth8fRrva
UHD2Yz/zeFnoFYNpiD5JOnFlPZFhT/cqzz3DbVK4XcQZVaw7x/ekwMJSMi5dL46lUD9gijjT7euz
2hjx+Vvf7oMXwxGWm27SqkCn14IMX6mHFPC3Di4QO4+lusUXb9YmHl68djxOsE5UO7tDStb7On4z
lHXD6mAxaIxkmVn1i8ylhR5lEFpohQ/3y9hRcyGDVSeOKQAhQcV2E23EyLNuXaM4A0OPpyqa8Fb2
EqtDHU1ujwVwnzLdRzpvrsv4Fz/dMlvB+tt/DlGKLAMExgmVCFBQo/mBl/+qcD9ZSKfXt+a/KRXG
8G2VZbygvmstsdeA4fKvYoQivHK/tUg/mGm/X0kCbmuc+7KvTT0FOTzv751EjZA1jmi0M0mBUhqE
R/m2wBpOI0IBmVd7igZdGUygtwe7khTscTMSk7/3Ybh/jMBaNq96KXfWbgcvhWldaeTZEEMgayEP
PwX09cSw2s2DxEX95FHahySDZ6ib6dSDA9AMM4z6iiWxKiAdlhTm1I0C3wL2Go0NqtovpU1tAwlk
sjh1Cr9v+541PGP5npyhpqEb/QG3ZAwhOIpP0sGNQuWuK+bcS/FP3rgnpuz7jj+kaQNHy0Ns5UxM
/teeaIbic5r0EX7N6w30Nhtexzh40uzWU858X31Vv0dx86LMbePIz3VurNAkKJDpA6asAt7WUURS
pBZ/C7ZYig0gkaUWi22cZqEYCzv+a34BkDsjWCJmyrp4CaSCgJRFVhEDhxAy82KYFPm5L5gL2tja
T6NCbknKwZvjY57I5f9JsDQoXzGg7gNSnrjEuATzihemuJw0pOZRGL9UIxj5Lf0wsNigXJSaqU/8
UNmxZCKi15F4txJn3XIFBOky6aTSeYhSQXP+Zv4oJ8HlU83PDxWxTp9Y0z+r3KR1a+qDP32x177g
B4FupiEkTI/rOkK3d/3eyRcMvdk7YWPwNojMyUw9One3Apih344KAAF7pHtLq3Huf2RITPLMbgCn
oyzmAHvu5Jevr7Zlec3ma4po89ayMKs+w3MeC42oGphYq38g81xuRkBvaSkN0ovkeMo/wZTr2Zj3
LCdeAW2PWTfD6Gtl3rD2fTUuePwfSuJj7WB5QV/HuMqQFTJu/tJyKOSyN9llfxatBS3er02solMY
wy2PBCsMt3EvpUD1NOjsky0CTTG+HdyXN7whcZl3UF290QFgBCCw0ULOCeAXsVEkxJGS0fUTfGgG
p8oKmbtlfrtXE6eUNrgcTP+TRP0oHmuLCDk3UhXqiEOJ6X/58cUaPLU14TtNOaBB9mQmssDG8xXX
Xo13iXY1CQL0KB0iLLF9SJ+/zP0h0eXiF+GsQq1ti3J3wYKTWYcNhnjP5n8Y63znv6oZENpZyyZV
uCOfEatc+fLU5Ie4uWUrrR2HBiSZOAmE/2ADvTTCsX1jG6ySMPHTXtv1+Lo/QuQiCi5jaXOMx+7z
4Nnqv9L5IVdYHUh52jIT9ENmhcWQkxhj19bvAuy4BQA2oAlFYDzZXOIqs5zqZ8XdhI+SrO4+LX8o
KXdMFl1kYUaEG2Uh4VI7NrCxNK6toUutDAG/z1Yvlb8wH1CWY8jOudR6r3nAnrjmyOZig0icrd+j
ygO8LwWy+M3l/1TFz+i/VnUEDmkPlLfZ5mnO9td/g/NFHbQJPhRxRIvLYO3ugkiiIoglsKZUhAMz
jl5xf0MVkfDA5kjpIB4mwzSVhXRHj+apjoMVUPkabS6QEJvr+wAcIwMRXTPH/bcaw60ZWfeplRJS
VJX6bCYh7/2xchbP+JJQNuw2lk5YRZEAtOpug9IGTWEjH5NrCkcpfYcbDCZAgUvBHNaPXZeU3NKm
AcrMoZs4KqRjA7SyLX/SmZ0wmJkCE4ldGRGSyibYZqKY3QMbY8cGxWvxVx+L6fLH7fV4IcYcSLFR
JiSXVu00xlwAM6fR0Wzu5p6yL5+1zImDddGX4CPQfa7Fe8K1WP0KH38U0qt7s05ELVvGS3WYIG23
7ABXs7OlGhuYG8gLcY43zZYBE9+P7coW86aQzKUYsz8BlKoYgpt5OFQ1npGP+aoSayliUppZj3tw
Lji1z0JXnH0ZNWYxb66SZOAAsZJfM1wfqCJ8hpQz/aOwYXYAaZPueIy6CjLm2+lTiwCE28rzh0Rs
npz+zA/m0O0wvLUkmDW8H514T0AR4LyrBYv/Bj2DAXjSOvmZn0ucaO6lRBihW/Wucq0k5T+zQvFK
L8un6Q/OvBlbVNM+ah2d4ROffYUWR0VBh+AszPbgyoCQq5xZlryUP1GJMcKmzePZEbz5fdgnWzoh
jeEK+rc4Wn3/fPsev1Y4QK/H2uhEekU6MHBDnByyyVkPeSOg9QDtFyV8BmN2m0MxWn1309KUbXoa
su8qweNzp7ZNsFPSSW/19IiX9RRmUcKSU89FZ9MGCYoboO8uvnyrrrjzE2wUu0VuLD7rZjgVFxa8
TmOdNFGQJhBU+gZOMpvHoLJLzgdnoT3lhDULO8jlqp1PZoT6PSDd/V3AaGaDFNZjkcSJjV+YiE7V
zpOFkEWgwDi4kUcCRCwM95RXTHX7YyR0bqd3vudo5O0/1tMS8hJmIe4F8QaEbUN/qxHnlw2faBvu
FBGPCAg4wC9h42aI8J8DIMiCcvLdFnRvP2oRzp9MAOOtKr0lwcgnULmHp6Ep10O1gIyR2uVMe3jT
3m5AOk7sry58G6UGsfkgmuGKxY9aSSUX/LBZXkmJAwW+ZwWKm5ZNNcDi8vvSqWo20FJ2yPgY+D3N
I/38+VylgW/bsrbyAfsoIdJR4r/ZlmExu2UgWwyH8buV+TqTcheG0yUIFoNoBwsxApFVlF7YmnvH
7KHZPAk8XIDe6Ug9GWc2A8VTbaTyrMtJ4l8SvOyO/Z3FMZm2ApP13oQRfzOrWXEGQVXouA7N8Iwd
GVaLlaJbnRPNQP6UY3LzXH2Dy2dK89BI6tRalBm17tsJIV5UJrnl/6lG330w4PTsu/5IG3nBgKH8
HNUaEl+Gc5bqszpRoWT/lqisgLhvg2XuyHsGcr143d7JNToqttjwtoMwKba24fGj6YQUWTJRKFuD
Uq+N4WjnAYbloe5wkGhiQMCg+kd3zWaRPTYN9F17S2BnkZF0+wgS44a1gIvz2eBu8M0eMBhF7K6J
pVYAUJ+yRYucULry5o8HtdSh+Mo9HC3ofbJ1gujRdjnWDlyHKcAeT9Z/3r051wfV3lt7S09a0NCN
MVHXS+wXYHZUwBCSSvS2A9QMs0MWz+3QLK6QCZq3Z9iBtSQipcxS0fNDqiaBk6GR5wX+6iGSfcyf
dws0do8KDEglZAX1tfmqMaLMLr6xo9URhCIDKZ9oX587rUgdOSOxss6t0KhowzwLvGxVmQ9nH0S3
74GvqbBneXQGxcQnwkXj3Zw3iwxB/+c8wRJGfnRPn6EaZEpdj00hJ5K51ULEkBrI3AjXjaLuMRRU
jZy/jxdn1l/BMpI7wTKtHlmbApl7n8xFHEHaavsbQzkoN3t4bBzbebLd3Nygya+zqELUiBTmLXUP
Ki8OTIBiJbGKJhpjs87jwh0g0N7XRYmcaaea5pgHUDdQti5jhpnuBYCEWLQuLtsBBA1NXWAalUja
mS516jkdgxUsoPMDm68KG6aalJ7t+oy4r+dZm/REWTWjk+jLpd3N6XbSL9tE4RFovfSyZ1XO29+C
5mA4HZWYhscEdTUQhRnf++vvgcz4Nyxqhn2JDcle9g4gVelSMXUqQ90bNnlLtKWFJ+tw08xNLyJB
cmJamMn0kdd5YvmAFFQL40Yrp9JWN1fS8v9F2BuO4cVRvYI5k8eB8qeilYJ++C3hzJVvcvcfxBjy
/Lvsyh0gW70yI1q3kyQcDDG8idzRMbN+UdMqcPkmbCOFX/K4GpDWmxjwcJwN9iy1rfTzwLpVq+b4
JBTlcZ+7U0+cFX1HBRa5PyiTFcflvN4XHmLaiNxIp6bOxFIpl+2asyV9KDaDOufRWhFKdBm0//tI
D1rN7DsBMqHPUyUcJEr2+gKv3Ucf6fhainYo7R0NPXu7hEbXuRZolSmYrlqw4Yp3FFiAP1+gR2os
x0YcVkCu9norT383DZMCi96Jw8h9t77MylUs9ehnpkcoMOPCjCK1oHWHT9VOS7AlhsR472sE9RJM
ztAmIzMB9itI4PkZiqbdxTkqXjlVZjS/YA+vY+6MHBUaBx/tNeTh/WS/1SeEE0k2nqAOHvgN93F/
WQpYqM3V0Ho3Ji/+F8NEGs7pbVWFw7Fu5k9J1DWoSKDpiqJVTFAGC7IHdREsOAleqNaz4frUnD4q
VwAVoxIUxRJr8ZX01MTr6moIfvE0HqD4VlMS9WJxnru9Boha9plZDzfy42ZldhzWD3GwqCu2bMyx
3BYyRFNHtEvE3wKeQtGZwnRMjgWd7IZUGVmhUt4Dkh6XrCmoxkFsf7SZwn1ZgTYmdP9ipbhQ/E+v
SU3Lb/Qtbn+CsJTWPigdq4aZ8fui2DP2WKLxGuu6lFIyjylyW1JaAbLsWKF61mgEsMJox8+scJEV
k+tB3CiiJ71hzWs3Q4PnnLLryvh6XulSgs6UK2FytGvZIH2CxgKLtW8dJ4creZLDRulOhEoAstq+
jX9dkXgaqIoj6huup1dNgYxL4AlblJrrzYx6grZW/B8JjBnv4NLl6GjtoqBxwTWRFOTieRiuPLRr
g5VFT1oO7I24C+NaSWTD9Up4080Jjh3PRIN7LvUP/NZdw22fw4WcjLjFZnpCYkHH/7NbYOaorTZB
kAn3JYmCvKCdwQa8ClJYXgtNE/l0Rf59+iiZAMGbHYcjkvkCIhtBsYNCTJTMwApLXdn0D9Jc5q65
GXKqLCtAitjd/K0L+0pxKrKNcRvvzrz3w1MlSVZ6z5zrCCjl9X3l+Bp+p1oHj8I8ZyKDL4PA+rRe
GmTzXrSVyUa+TUKq4Biy7NGvamrxRaF3BQ1BNefhEEZYMMjgH79MMPYu5nVNjoT/RJlvUJgwobWM
R3+/O4o4fFjhjwPBHVI7NkxgAKrjBmpSe0bkVMooTKHF5cVHRUK0tkMoGbwCz2FOEslO/OJSWrP9
jZQG4r0gaxpL/1Xp69klnko1r0mIGGUYsg3oBM1SZg9phLEjKNDg0tFY9/AG2iaU0YTkmoP9p0Es
41VQhP+0Oa99RZb3zxeTlLIiNGpKrgjqjM3lFMa+PdUc+wShkaJEpq+a1ZEGKuyZ9VJmt7cLF9kf
UlCFtYVPPUSiHyS2ToBYnkXfUWR8DwKneBOJLv7h3d0JRFWlnteZAopEvhiiARdj+xu5MANPc/L8
RKbPYVM4Y/qX3D09rWykSai21qLqYs6XlBVdMkLc/q6Q8OvttPQZGWIPgh2lvJEji/eTMLUbBFQc
3EnraX+XjsItpMlLA3ayfpgjebWNGg94Oa755z+ySQmbVzG6k3poHwoi7+jl4KdUm29AA7OBu3Xn
0k8kBxFvrNH6a/4X/XYQZZwhqkk67aOJ6n/ng9Z5mmlMnXGzuyy1MzV7ShwFRrJHbrJIbLuTaYY5
fsKwr/cTmkPLBnUhJU+2sHRMAC0xVrfUQf/chQJc1HL5fY/6zX13SUMbSgf4PI+GSZub0j1fP5ov
X8qkpAoCIAjbb61MvfLEgTVUcAcg6subpS0UjQh4viwXaRA+4x0r9j/Dqvl9jbNAI5sOIzGcBjT4
PoeNNtVaDheil0dUUwHsDjxKfRdLYV29iz/LrdBjweBrHfCEmmTlxeShKxGSTn65Y8Z2yl8sPuaE
M8AGzqiqu3KBi3dbn/tJ/gia4vqqBp0C0JzVSfMMKZfTrh4NdJxSEDNjwWw5Ll34BgsskK7tuy7p
aWR0JLVWXYLX60I1SUWoVjZvOwMuTTZv8bdmpFwml80pT498UXq9Ahl20HQwSTYQ8LLXuct/cnOk
GmOVyxxvpxdBrcKwCbbVTN6/vEk620T6acfqOUUxZewfKxTmE9hHLOWFBBhzCIcQu6JvNmmiTZMQ
5sh5NMgnjjY4XxQN/1CVcYDHNVEYp7/37rAEOC/CNYubFlyNLt+ahTiONH4km8FK7H2jR1RiJv82
LgQ8ZEjCvcKtWSI4HcHeo6xZ7FILCPv9w1qcKhopHT9b9HSwV82jX9B7o720mRlvRDLTfFe4Lvnk
7ncBYE5ce1oVpl/prBg3r1G1P5gv0Lam+4iTfSbc9ZCOEZL2AGcqlxQ/RlBRGNCeRotDNwHF/5Rz
lAbc28AaFir5gwSR/er9UsKyBiyE+fLgzIsynPoCpRoUmsSxAcZJXcnGLfJOfTXNsab2jKEyzjYB
WLubo4ropk8CiHukPIKVGahNNyt0XjsF3pQE9j8Ie5CtOdnAV+XdPYH2ba7FW97FZo9FImDVRKTI
+O9ekZjKTI562AtgNXv2ta5X/8tViSVugEGAVIiIdRhukEnkoo/q9GrxH7hY4AjryGJ4/sPYMol8
n9h3elZL4GaJxg5bvqq8Y3NC22I16ZXPd9wPEeOFKJvhD4nqVZMn47/ytH+d+WMBXedEqE7BlASx
3Orc2zBAewziK8d0Jk7O7fT/SSy8yrPQtxCGc32/Y8oy9NwjdikpX1Y35s2CPJ410BgXzbNSKzMC
j/oTlY/f4sZ7UQpSn3iEBUhmkvZZaLEW+2Msfw+MsKG7QnA3XWs2AgH49VzLrK/Ooq2HnIR+ClsP
j6u0UGE60wGZWj1zOg7QOuHOYVblLsSxfok4h7URC1S2y+edSfKB/Ybk09kjjiRcQ6bpTpssAV/M
b+BYKaO9TZZy3wE9k7kAhl5bZ7Um8VN19MIEUvt1S95Y/arky/MAP4FaSnqChjx2Bdfs1XJAUMLa
qn1TtcYTlDsh5LRvdspYhLnitMT+FN8R9B8KJX5DN0X5IUp/H2HDZW7Af/H8QVEyCIHZ0KfFk7P5
2V4h6BT1DVFjJ+O5AGgr+y7m49hwy0VWUMMRHpOFqpgYn+Cf4NXadrmPart2SOCruvI+jwlk5M9G
IyQ9tZ2YcdlD+ZHD/CrCphN8fJE6u91JA35ON9Y7sHTDEl+B6bfGx/81uU5mlYUN/vtj9FRa12vj
VGdjlfWHLGCpyZjprspZCEJzL6lTgAOHmP0uq4lL/FkjHbdNYJo6nah4OyDc8wQtSBDB6HTrWHc1
1Z0WE6GO5YTxDhezanA0GNwRjGl+IWcjUmWTCtOeNpL0N/nBHIGgdgJwjnif3NoI6aKIokUhpa+f
NC3RC+BwNbgyzkFJeionAMyE5sX28ERCY+qFAtkqqemiI85INtUlVh0d/MsPj6Qds5OpLUbczsSV
C1YxkHfJeeOtdJMDUZFWxo+icKLa0UlSe/etxhvCKTp3nAJGVNopst0OZgTBu1xeBEhCRVlY6jZw
vXxvZmZdZSAyYPEz2tPzfpMlPtaUWIAqEjqBDEtvcrhnLnblOpE26l1MRILsZWNd/C55xY6PRoge
4pUPeAQNRRdkuMSUSJyyFgaNhqngmXGDvJCiaCLDXZSFZ6Cns17UwN4nAYEhClUz7u7l+ZD3qRnv
zbLZho25JYHGcpNi5o2SD623YMriXoz/rYSNwWdUbg+WCdFiFJ6mXVj7CVW02PBNwb5wKAyuV9xn
kdjABl/X566K4gpcvhItyx8OZ7Yj03twBp3TBYICDMaRMbK8yXXrCi0Rr6HHlptPmB6PmpckRmqo
TH3/O0oBCu8ij52V4OOcApsSxTc1uH0thVKxlAcXlOX1uCv7o6pCyi4AMqZrMcmYUu3tlwjx2SED
Y9j8K2n7Jyx3WHvB9PffwXC9bFUFhLIGgdK9zKm0PssPINNvSWFO2JUZsckB1DxHQ6ySjibg+L7d
R7BF3+mFWlU1PAICrZ4t2YpzIUoRHn1mTTN9Wiue6xjqt3UpMzNK1I0aw9osWv6qdcDb97pVlDTF
H2p8/LNerdm/dhJPCeKkPq9zKb8JC0E5v6tncanu6KBkp5BqR9D2GFfz+Oaj3xCNeV6VMoYHR3wr
nhOwdrNushgPUf6IyCgw1Zxnl7pOPgPv0RzoU5ZOW7BJIsYL/RKgCTLg2HNI+toCXkqv9xNF/3y1
IJqe+GXlslhEdy/P9DWgVYwECgyudsit6Rocz1XVo89GQQJNe1nSvPrfbBVegMeYvYn4ae25vdFy
X9MSk4wPW3vblZQWVxmmJz1AR60DOoC+00p0y4py1TZmSKDVZ/e3uvM7EbgPqpa+lSTIsXkUy6Gj
KApoSz7GN1E8d0p6TAsgLD9ggmBBotFZEX01tQ+65Pp/kvSOLs6TZ3NcR/vpqwA+ApZkEuiRBZ2N
WCuMtaRK7DTYElX/elT7wQYm1ZCibbw1LNQosQ3rqfU4ee7KCp7lGT6Dvh8u7wFI60hIOAyqU9Q/
yvl9/zi6xsYACAeLuItRcT3Eupf7JyccUKJw0W8tha5Oq2p3hFsdpHo/thIwfZTW0UbB+1rZlr04
caGMh6LfyvngNWc/VDH1sw4mSh8OjYzdK9CcgaNK87IQxuvsDbnQWc33GNNwRNGYBhLVopu1AbLP
31+NfSc4gaeX5lfHaZ8QPXAqPqErzyjRZgnX9V8cj21ytBaL6jjYU8Q9xpiuf3sjfB9he3XQLI8u
zn/ONIXKvdK+ddMJ/9MCmjU8vRkW1Jir4/s/9ymA4rEl/Cs9ykE4V/T3gPQxdOhDk4CVx8MNWNJW
Lfv+5HeJYcdkZPx3oZPG3/o+Xz5xwGEy3cu+/v0CvRq8LqgtHe0mDpEbKhO5dwL3DPcWC2MAs9+v
3MP8wSjZfzgVuEWb3ux3oHKi5HocFOlG5cX+L8CauY56xzurM8G2ibGEVMmFvLmymJqNme3kbv/R
Tyo/UYfmWQjnZEly8PiOrjhQDekN6zMVxOGtOvrtGI/0lfpwKoaxJ9hAcFc3hbHAkDQeD575uv7x
nYS8xPS7mFEfQ56r3vgEvOrC1xluCEBy+2+xNtn/T5FO6ZYbxw3bxHvvxYmoeJuoVHJ4GlTgHJXu
1B14ARnH+Tov+j5o9Y+8dD4DWP1Yxw0pkqZ5XMcP93hQhbyjd6i9oC8Fe7FdRX7nQZ3qJ4JLTgJk
bu1yj5ojT2/HfjQhFrBTRv1CwUdn47/3CD2FcjvrBKCabV9LoyEPEKiFj5HNQ6XR+d0zay43wnDP
f0ayAH1M3kD/QJ4ZTBW9loz1p2obZ3Gz2/oX/gVWpzYTFxlZfJQaaYYQaguRaXqJvkCs8veShA4u
2thMNNetVJKZBePLKR2Y/sDIALHlZqmMGP5xxSjtIE8GObk9rmBKvdotsQLg1MCH9WtdFn98XG33
P7VtWrYaz9wx+Wjpjo6MFnzKKjIfJ6D/fXpiOo+YU8zyXsNZahCdqmskXuIt5Q53IoBis9Cg6FMR
yNagOdDsd+k6gGkL1Ths35ktQ5DHXveNgwL5KiXvMggPEGJtI3KexR5h7WzLakKTVOENOd9cVwvP
2zf1T0yMVscM49VNSkNeVgEO/xIf9IQ6KEQa5K8EznFXBNF9BPlSKpouasL/GattJYLYkCiwldQ+
u8bbawNpT/6U1qStOL/vZZBzmdMKhuj459U16RSuBymmNtypr9zlzqnSJ/TDwEF1VS4VzwLFFTFM
0QlkLTZeJuQ/a+vXeP82Lof53H9gq3eufiT4r4aFEDW33JEvVDcuUFFgGlVymfaIhHt1KiU8dvYB
cG/MgXWGcK6UnkqbtztQ22qx7vzkiE29hzRv3hVGIzijq4wVnM3hYBa1mZoD/pfHMWGL9J/TRbTv
NmUnMUDEpCP6FcqBcKK2MptvhSAQvLdvpdmB2lluvF/swywhcVhMH9w3efQNWNHhyfG6VAwjow4p
MKf8de/bTzkZz9QxPAcaq7zV7eZhywulhGe0uNEAJZdUppfPVCJvLJlyIvl98xRoRNSO+Pp3WS/t
ZMcEyPocyi+FgTmQmc8VqB0CNay8S9bZOCiyhx8H0ToqiUSohiDAzgAFrTPrmi6f18xFzHQOyqC5
B9D3PWWAEO0ZhJ9RIix9JJsQ5ggdnBOU3e0jBaJoDZRS9Rt6NsCM+kBMGBvkPh95ATERveGeADg7
jvFK9obcNZ104w1QPcvcC9kHY+Rd4JPYIqNJKMrnBuQ55f5ttMjSyEmQk6wiVDdRwEoIHz6M1LS+
SFTq5gQF2j2ytXI+qHX8xPR/mqc8+95qQ5eyOGU1NxsO4v84jF7y7Fmv+rzqmT6sJhPulq4roEg3
NjNMboQmOWQa7KTksaihaqcFN9bTnpDihWQzI2XzLxxTqsXFrSUMxZXJMnEZSLtsnyptShY1gxlv
6q0+FV0eH9h+G7qkNZacwx3HzdQIoHJH3um2CzMJugVFU8jDm/sUYI0WBlux1U05cEt6GAfcK029
v+VRuxWpw6A7lRNmm1okckkAdD1KqdOoPcdWVsjM41gem3pym/uHTi+1D5P7m1bsdRAVclrY7mIV
XdRzTnw6c/cuOvWgnYiJh6BFqg8JsGtxhvq/cRXE85mYwKM1F9/PPl74zkolEsvF1zUuOxN1pqPP
bN1+4E13Mb1m8+z/0fRXJITJM7S1SFd044dKsKZqf5qYP3IpOmn5PscVKpq/dzgMbY2LkV7GqdSk
k2tS5VSwPxipfj++5Ntjjn/IHYuwKxbNUHHdSTOnpUMhqw/DbhgcttzVwphH5ivXQMwuzeOX4pel
8rOpgRWTcnIB8CChywA29NwfbUzj+XAO1i2bifiHcSvdxM/JNQziEwqvlH1SiaZc+M+VVj35q3lE
nwOViNBLvEMtJUSDU+WtkCCAOX3jCCX+D5150SokCQ/nfywrJiyArjricE/ys7Ii/VgwR5paYUv8
YW2eOPmHkbLemipAE1oB3V56P9gLxoHRjS1IgsjaGK11vqkebi6s63hG11nfQgBn9Oed1/gR2+37
TWIl8CZDe4VzbQ3oebYQx9x5W1WnPsPN43z6DlkLl+dxKBFw/ddvfrFlulUwbx8B0PlXyJ1yAiiJ
mJPSvSb4dhVg19MFi13sEnhq+pbBGzHlRvgfxnjRJqYUw1KXoZEHSF7aqYqIhZVA+9JdGFvGubu2
UE72Yevq+hNoscIrVcBPVswPMTxUdQKmsWulCBDhH5eyU3/WfP/uVBbPrQMfItdh2ZWop0lN48Zn
tPtIZ1K1uwWcSEgwHA8ERHREMEM3otFyT16hA42Gwmo6bngXruLq5ESQ6QpR6NBtLtHy0lb+AKIi
DxTcM3DjKpdy/iXs8uTjFAmGHDHwUAQTYSg6Q2ABHlYYTMnyRZ5w0N8ILFJGlzeG/UVsSE5mCWE5
n6JWYBAII9yKIoQEnTu5cvVwYItNIQ15BcBXZxtOOB5NNZDjI/pAB1zPr7RatsIsVghjjVYb/a8d
4wZb8aWkd0izWLM12by2gjSyynB7kt9FOWmLzhSamxv5pP1ktciBzyyu/8Gi+6wcfZBZdop+Gg0m
o/K3SoDDyb57W348NqsDOjZKoBMSTI3JRySGvyLWCC9HpP9rY8IJP4quYULe/MGCVb48tSZtER3O
NsFdGsk1duHyuzCkBr+h8Dzq3j2ho7ykF407i5rsKejSmSCIrM11oLiG4EgmeLRpIspMcyOOkTjs
CI5K/FrsCnZNNU7RkEvbwMnAoPtJeK/aRdXu+Uctw/C9sHEEkILC4yH4TxITCX3rrtzFCf2T/HWo
Gi/IuUiaXuyC3Y3IKV/a+THyTcTl3nLHyqbXHmejRyPIYqz6e3Q2ysBXqYIPe3L+ONm2pBx0oBLa
cHHxccVX1e8by1qJoza+UFX92Vq9w52N+Lv7aliDvD/WukY0kwnl5cunVgnFVkwtMupvkTjNDqVb
awPHnLmikqYN5OiFjcFy/T9QhywbEvk83JVrzQWekjtUoQVXsrfOiB/cuSo7a9y/Sc0jxK+vQVLM
4Rja9B5OcHYT9I1gd4QaHQhadIiC5fXA/VmbyXbYVJX2itNwoB0R/xMvY5geIWhNt/zJjkm7Sz+M
hpyoehc4ErhngS3Q209BWGh4AcLFuzx0UdGdnouayN2xQ2mnTzJJIpTIu8XaIfcIvrYWQmCw3e3V
CaUK9DRxk94kr/72ZfzlT2tiqq+J/AyZSpvpFlOEMx3NXvs3ImY2jC3KLATTtooXxjiGgEob+3aU
EHP2Hh2a0AHwOk9HWAd51UAv0V90DdJdY5BVVPuhQpA1z3vQAfrBAqCe72ngoy6OJE6xhCGxSECb
buTvYY5mvEyMmJLwY+XMIAzmdvcajORLTleLOdrZuzFO6PO17oMSn7fJniLmTgcE+MY1Ve/a9eZr
m39SDoR4YfQMsl0c1jsCVRCx+eb3zPqweHsMSSRRLMy8ZqX3jm2TMT0DrnYhhspsw67Dv8awFTvX
9sz6SELOAArpug36l2FCyz27MGaXFpF8+9siF9Q93J5TA9d+yMveTT1gupEUKWeN4PIA44Ft6A3C
QEWov79BX4G5o4SUk0ix+nOlwHSApWGhxG/CSvxaycWl3bFVq4Q6eu9ri+kXByBD77+Shq9+ssL6
RaKhvcQ6GU4HB42D9fbTfIcvwJX3MT1YMuKWuGwpP533RFZ7lGNQbQyGHnw992VsSQLgxB1mD0RT
e36CCvRqDjI1CuNlVQHNtrLdgWaqhqCJvbku5O7dCUlRf9ELTRSkqTW8x+HgJOQmaexto8+nlV6B
bTyLifPrExonfYmhx78pBlbRxD5KB9KbFmfPWSZhCZp8U3G/tZR3W3BQeAfm/wh0naPbIj4HrJxM
zdxshdKRV055Kya1WBmzlOEfQA7egvVlgzjEtLBEp5IUa7+eAZnP9u+H4utQ1qlXAcgXeJvzz6aF
mSrJCoSyKPAVlJzLOOTn6tNhhslOa64z/R2L2sAydqhNRIwpnWjr8UVjlco/tNR98cXT7/ClcaWA
qzA5DBCT3YJhRxbeKOuf1T3Z74zdCvNVpiwxcD+9cDEdg22igJbgh71GWVDMQskZxqmsxgG7bKOo
lEfE+pRNYJngbXNLKxShYIfouBlT/CE+USPFs6Dtz2tHs5bRO5WkRDxWiqGltjfgAzk9j+ME08Hb
4fGpxwZS3tg2tZnc0Ix/qY2gPrNmiJUyClk5miWByLr8X6vDzO5GeVMEkkmJ6nogVKQdElxlxw/G
09VRNCfuM8p4Ie7tmlDXQj9RgdpP6nc8J1Wu5TgjyyjNVcTIhg5RA/Sol6AxgObKMM9kqy4Ayi5+
Lz7Wi6LtwyCaz1JK1ty++1oXRIa4pBjfHXd/SjBYyYVA6uOkVyLWJcPzdFjOMYb77dNr1Z4g1mQ1
LcsmHxX/WHlyvWAYe0IudNM+e3gmYBtpPUZpkSpkXpaPcqW71DXlRYL1xQWr069IxKAQO+wzlrE+
GajsOHpaJdj88vD/tmUpo9bKdvlh/fKw1ITyi/1lqPzhpT0VVQuWRN4aDvY9aL12LjY62HOXMwDo
AV5uSZfQ4cGN3QHB0qU1QFoIpPJAdhvaJY7GgolmNpWjCn/mvwBvv2qJHaK7RDZP/wk0QEgfQfZa
nRqBCuq8G4rD9wDweb1OXD2nkyS/fxwfP/htHnyDUh6RdOf9ZuHZiSDBv6omn8xxAVuPpRXlb2bD
pU55OHsf/R2X94PkY4trEobkpWRywspvaHNR6Sqw8Vo8Nod3P8nv+gPIYNU0NzfHlfpQvn3du8i1
b9DSK/uUu9/8OVkH9ugiUiYksJdZ9ociaYO94KAvM7rfo/yR1KwF8xsxyd20qd/zLKG8WExNEIkB
uHxvm90JkUA+RrqgYOS+MuNChWgGzinwcIgW1TzfZ63qVjQKoqLx/99beRGizcEo6Km+5IQl9ZkF
ssp7Ec3dGGLmHgL42Bvf0ucTJiERVJM5Ra+B26kQh0+SXgZwwmr102gjFKkmPFioUtusZFWinJLY
Rim547c9MXP/U5oOGM3rHLMnllDJId62GXNDuGwWwce33ViBZzeTt9HEH0Ceph1ggjRpRzRnIQNx
A5hQyBdW1Mrru9Oq6xmqpe6ZqmlILUF2lurfJcs14TtJ5Hxx9BfU588QkxfC5ERX8Q+lRm/59oQk
FZqaWT/cbpiStXTGqA4PPyyzMeBgfynf7QcloAoLfrtMQ82U2Z78Qi08FniQczjwgJjCrIRg8oAo
WLCzR7WtPoewVbAosn2MRIGJBAkgdYontANbEndQ7/GeYCpkRfzx4u9e1hcems3WuZ+Hn1ZZDYSu
UuK1zjmGnav30kqRYtWJFEw0V1FEoxWR0ZkW1qthdqoiq0NAISyZvwXVYfJr/Q5UwD/V50AkdjiF
AfUd0RB+jBfl1wFJL8b8BtNcLUAN15aBOmxE20gpUatpato5ZmfpIzhgVsLxQRTmHks/vYPWNuNz
9P6Cps8uuBc3VL3oNPSXqi4Hj03WZcKdQxHu9LsuZN5k31SWyiwbWbM1DNn3TiG+k7zoPmMOGUib
gZdlfz/UF8hWLnVpBUDVW+hTVS5V4dcP8siCTrvwEjpo5hshjr7M0AfuDPViiFYqyKpcUpgBRBuR
LPqrYxXWwD6MRYATdTcF+myBExeGyKst7T+RoGdGpqHz3FXwN0BXPk7bCMOu6pVPdi+kNLBnLsmA
FkzmyPZwM7ya9FRIrUbIWBpI4KQAragKeaRQdzJQqiB/MvI72mXdSA88ljF9I5cowJAX+Og6C411
8TYIy4XgGiqAPG2H5uU802T9VPzrACfr5cK6REP1OMVHYMsHj7LsUDm4yMRzxeqrS3pnCdIYH6kh
FR502NrLDSYdr+txZ4p6GDiiQyDiG5yHgDj4rENSkCTY3ZQRs8UaDGZX9BxKBLJjw5IJ7J4vGefM
vJaJQzODAF+2TyNXvrdU9+8pY9JKzlUSx2+TJH8vovMf2vuJUcWKMVrLGmdTkUNwusSoXS0rQukR
y+0zLum+5TiPT2UnJKsogJREyfNFrkR3AB0OtfRPlnpVVW7ge+ZleDRBNI9nIFg8jzLrqrd8kqVd
skK4y/S5CRmGQfTS2ejStGPzs6R6+TEzM/q8iVFHWaWRvKZ02rZNI2/zCLqaW3Tbc2/Wv0U5gs7l
wRQpIok/YYJhmePIs/olvq5XA0rqz95rAvzTMmbZGaBaSaDe8XL1s6ridiy8aW+sSCjqWjMHwghR
G17HEbFzsTBnpD9LQzkoWSCgHuD+L4Pc99Q68/hrIygCfIhab0mVhJlHOytLF3UWMjGjtpnX/1WZ
ru7ooKU6VGBpjNEiA+HWhEQVT4Hf+dig7uzZORTMaVh61mK7U5z2qBpAVBlI8InLuHhSEF/adkEt
jpuPtnRKuRXt1yhpmd7W/IqdyJGfeLvefNYadnHO7iTsTQwYKaHBWQ9aADI/jYPjECDVPrZcLiZQ
9+q1FIoGWkeApIdS1EDvnfrEGci2oPvefUe6LwCK6dBkMmasFh+UCO2lj9+thEewDxz2B5914FVt
vVv2tbMcwSlGA8G5owWaxCRJ4+XDXFqk1O5/xrOHXLaRk8omi6tTkQ9+liRcJ/JQkYbc1WNG7n+h
lG0SBpLJsk25Kp95I+8JZUsT3i6RTO+tVJfVAUWadqSUx5ClniNmdYhcxA7fns/0T+z0YRYO1QCa
gAkWpQKxKFR7USp8d9xpgwITLUgpOgmp1D9g/MNKjwFhHSHjEbnee2KnY2NdN+7Wq5LRXcJcpdUJ
s5bjothmn/q1GZB5tC/0nkEXboh3BiTUWbWPh6YVdcZZB5ombblb5f1Ks+rkgd6aZKgiJgoSFF22
J61BAn5oFFJfZbtOccKmHQ44WgQ5jb8X0cq+BkPLj82dU190a2qZetsy3C/uCuZDEIIe735k93Gd
sbu3EyJWy/uSCLF+yD/0Hc32BB42dotNrhsLFFzvvOlsbxoFlQ7qSRbPj43hs74Jx6jWJM/uJcEJ
YV9hN7C9RCS1QDs2MUxgvi5jW9soj8SmWzMRtC+cf/9Cs8OpZxTdmnYQM2EiuLrAMZbJtAS/QFIR
LTElOtA1Fo5nza4RSIOMHLmhsDAa84nEO/Y6MxUo7e0fPVCzH5EZIG5mDFnOqwldEBeL79QVMSUq
5r8xGhCYdKeLngbij3QWwYV0URMvj/kmeYcxbrTlk0kwZkYyo+kcOFNNkk+odfAktevWF/9HxD4g
/DuOfBM33StFeg3PxMJJRR/qsh3t35dxZtjq8gVOIZcycDhjQe9Ls5MjqNQiEgcrkWG2WLhNsh3X
1umyBO2fWp191ZkapBEo4udkKSG7lrOXWLUDEBIOgBbpTGE6qZioHOHwoR+0+yFW5P7DWMDGOasv
dJ4Ua93lsl2jcGtEWNEh2IdDOpk1uSi09Rh1kp4RvdwVJsEIL2DblJum0Q16oTxS/5QIMMBfpROH
y3BUKk+Ro22pCJuTP5Hm3RM00tvgi9DG/gZcLurCr0qYZMu45i7p7l5byNfw5l+zJw99H5z4ku4M
FNQ6OvfxTkuLbv1CJhTVcUtaAAqiIlANezKGLS59Yc9CA9GkcveB+Akj6YuokM4FMNM8G+jQPKCt
HC6JE6IpkbHZ3VtjFnY5lFcaHFYp7pjSuiREyTTTdZOlNG9WMe2xgxPFxcaWIVrp4bTzYeKRh1Lt
ns/KtjCt49x15aIOHooC6ut5qttRl8Z6WRRwP7psYcQzs8HQnYUD1HbANJHvh30cWVwd6L8nkzxp
ytseJK1cwpT7Fpis5mI4YguV+DY/BpLGcgU6Gel/R55EJIJuc0/O8oYw3qnMLcx/Xso/HYXUnzBL
bWam+Y1JJ3C4vr9wDyyTwUuwlZ/kxzXPSGDQPfEA9mUT3wMCHHuOv0IA++Ieap5sq//WDHAu2WrN
rIoYbBgwj1PtaDmjFfo3KsseZRiSq3SlJZkcWEKhE/1ABxKJ7tv8aNlTGsFeDRVZDHq/aSVblua/
e2a+V7WGNgu3+ppGUIXwMNzTuj1FpCtFHvDxwG4BPGxVI9EMHKDYHOvltq9z27/MMXKg/8zCegyD
gU+bDDlqExawzdIb9ZuAPiezR3ab5jolBG4iPpCjH5vRS2HHaxA5mt/HzAOTQDQsL/t+Dk+o/fFj
IFHRua80Gs8Xlgkb2eTDqau+VScAsm0Ha8J4uD3G1aHzaKdb/Pi5TqVwgRxmqze5/pVViYMfVmuN
UDgy7Gb21IAS9OS6ML8Gsj11fb9K0/xGt4JdeXvUivL67fyOXfwMEj0bDSVv8WB+y0FJlBVRrs28
yMu6ZuEwgU70+6UIBRjIJZ24I/aBveXFZdMpGVaWxHbjYZK35I+EaooFf4eoMW9Cz1dZSIaS8I43
gXexReY/fDdzURjWm7sT5w17EhUHUfJRJijHGBR36KXlhdfATsisvqur38YjhMTVJqypT59PUcIv
pH/pUlxsBiT7bhexaXTt1XF/LD5FMKvPjNw3JkzXz6YiCAB1AYXtZ47pm2TJCnpUH0ezyal3jWr2
1RiEC79j9ZOhZiOO44rEd6kv4gQmnFgZ3WqwF2g+mFyGDKCrPAQlyYGgA1r0bk6I2yJjbL4eld0Q
u/skhEnKA+T/rLLQMRm+j8aHIUnRlrl2f4PcB+PdQ11zh6UORupe+eUqiU7xnHvyL7Sdkpl+x8Uu
Y4mQmfuUmAUwoAxgC8upr64lNFfW1wQMmQRj7xrwA7LwtNabHbGc8At2VG+tV3EkpVWC1hAJ3iu8
acLKunV3oOtnoL2SHQzC2DpgfFlFEt/VJBzge6WveOjaVDFdoh14sCNiwd7eoj47jpdVKkNrwq03
DQHPhcCOiXPg1T+YBrpebxv153PhV02zwCX9L+Ebeu0w/+LDuN9zxr2jBLUfGGxg76jDirL/zHtt
igqekBaKoM987T9nuPAtollITFXxypHzA70rOAuIa5gg4Xqpijbi/JrAZLA+4oADiBs+m951uW/N
mQ0JqtBdwkI3cHP+yu1/0kbhtax3OzS8AA3NfY9Y5LaVkjhDhvGVSnvRyrbwPZG504XSkF0e7p7W
rSOXIm0wCcFMnQKY1RWJkNLxFzSTAQeberwuIYrM6xzGvusDWBqW/uyZclB2Q/w5Cgu5ymkeqtlD
Bp/ErkPyX7KxK9tC1NalOrkE/Ap+9PoZqNr8ReBdIzhdKpVj50sN/mLbbfslwVL9xAEJfAeJw2ao
syx9eAviXc2/HfcwtPBxNVOHwFxeb4vWQ57hRBo61y1q3eUi6k1X483aCHMQktMTPyE63xsjRoWs
Bn+1pTB76y7oNizsSEpPsXNR2FpYZOO8QHas5nG2Q4aYkAt/pp/CIsWzPOcESV/E45RVMrZRxIN+
IF1eRLcdsYPa0KbFtlPkgHLUb1OtB+bk7Z/omZAMKpVgTDP4IdhkInEakkgTT7pGm+wVrsOMz+mE
eUB953a0HXwFvd0T6ibBb3frqtcYYs25jN9fVisox8+t0uXSwzXo4j2aJR1wFoYxO8FErqmxmjVS
jK4g5nTt4sFNN9kBdx7iIcooTLdYdzmnU5bX9KXAC/62wDh7aAAm3nwQZW4yCxnrSuUJP9SyEX6L
XA+5HzGhcaQThxklcwg3e6Zzg/qZeCaqQW3QD7bukKUFGqQgVutN7yMRfpnpXotEOONMCOzGrDZm
VT8C2bo93Uz+M80QFE2eMFGsScIEeJ3X5IRwppMyg+X3QOXFVMm3pghlwHLI0ZB44HypTRkboOlz
3NN6DOgl+NvBA+qrVu5UFtd7loOGhAZX6RtE9fKxG6PFbR3pBTCEX4fU78On7PRFxIO0sWZ9Mn6C
wFJqlg80+UvloxibgaWPEPIPVX3Qwy5WGdmXanrhj83yMxGwbIl4dUF5CBpiXPicmmJbPc4yWs8J
selLaTAT5GuoAEVwrbMyU9ukNUFZpKWnbSEXxMekLPbPshbrZer1XQNPtKTkpJuHkl8SqXZICEhu
Vi0dH/pCi/yxfrItdMLegf2xkG0fQbGMGZkhRtAGpqDmGpdb+n72OAPBGF0f8WOGtE8gqV0OdE3w
PxxkXj2EDjRKiXywB4uOXyTQbL+Y6A+qj0Hn4kbu/p+Bo+XrPX5YtieAFzzKlZSfhEEv7/QPSyod
50EIrdPE2dloT+E425q0UaPgwc9N+8smSp+CVrSajjoif5xSSxe/L2srjgjNvmz9WFks1CnlM+vP
H9guH8rvmkbpYnblTxzEq2v4W16+y3j2BliXlxv4TAQ7kq8hZ9BBWqP9zMAWxK6UZpSgQEHTrgPS
KaOD349RQu6v0sXGNXnsokGU7v9j7GHLBjCo/9vro/RCpbDNrGYGeThEOYg3gUNyf/v4bOt3o3M7
X+9ZyeOxiVsCqnbRmxOZH6nRuVpAvSgCpi8I6c5TAlooo/dyPvpIPmueMyfoouBDpWRwMs8K9hwq
w8sT+Qdi+EhyaXNA7v0mGezQMKRSKTh/HeLENTQVoRoGlJR6r3Om9+OtBtoBarA00EMM0kFjdIFt
qqAxQyUUZQUv3iVGPV/JYBt3C8T5lF4EaSVFmoPgt7T0bnRvZ7F0KiWaLu7s8CMV1CyJqZ3VXUp4
YLY9+BWEKe1gKezitugt9rB0uQ+yNjKDatSFf6F415fmbsjp6PXpGDGIS3DmF5HMdCGg0SJZppE3
iVI1ihx3x+mkjWY4n8+M6u/RlxWq1o+4Tx0GYJfBp+IftQEPMtkPGbkKosRvRVbj7i1dWw3ZN0ub
pPNujeExi4XZCYuB3eFOtT87SV/+EJZzOMi4ZweI3c2mQi+2IUEgKnXTTQvnkBSlBIO35hCHm1EA
as1fK2j576HmhuCwyKvWpsW/VKW9vOtftaXIs10daZRa2nqq5Mr0bdawKpfZydt1M8pNwg2R2zGJ
9149cT38RjXGbn+vBiklvEbxcKawqFrWh1nXVPiBx4ScNtjdsxYk0QfSQugeO5wi0Maw0JnTkZEX
QSYD69fRyu69L1XMxMfzECYcL1Ws5cAHpp7Gatu+G60vOvIODfKjUPnQm6f5jToD/q6iFLTUeIbt
0V8J8SFWtVGKVA+AaqMXRuSOAqvEIoUl3M/PvQMIfM4KF2cifR9ssif6WAd+OyE8rn43tGZM/3Vy
z7qRS+azUOe+Ms31OoMR2F6aO6zyZTvd9qP7bgAo9F+EhWPVwTjfoV7Prs4yytzslGmBOu36snvK
ZiYy86V2tK/D+W1UPMcVmWd6AgLl/Qo4ggy/0CyA9htVZnuJP9JBZ8OrZE52coONxef2/ggmkJcN
zDOoWyFfdCzxPvoP+HtXg0tIHGmo/o1x8iztHZJ1cS5XEc+x8ic0gljRX9WVljjUS1wwmpJzxaPD
BhTK4tSliCFUcjbxHIfMAY3pqeSOMHPqKNsUctG86zroWTbaVLlB9YjJU0ErzW6I/Q6x2ewmIc+t
yXkScnfiZri+JMuQQxC/Pkurfol7RbHBT9s25G8/INnutu6ApbeEbFUiXPs/RAHBr+1Fe4PSbldv
XRofZbwWMIDc4ftTxwZvI5RgD62qFnCdlwYcZV4B+ZhH2ivD9TJt6gm8U8g5zxw8quslsp1uvAXu
S7EFxfdODQJscjB832A7gp8DmseuWr8LyqEQZcBp9txtTqATx1k/6Sm6R1EJPEKrJFYMSwhl/i/p
ZDH++6mSqGXNJ+gdHL0tEapmXkf9rqDXMcsfxBQwe+B8q6Y58pknhKeV+7FGFXmDes4rnv1tva4+
lX4l2SrOufzxbFdNwPhMkKCu0irn5ot9AYqY7PyQ5tmjj5IzYvg492o+zu3pTh12QhJIcCe+E3u7
DjzmTEWyzWezFvAlYvDJg3SLblytVmg4vbjF37T4kXZD2/c7qr5OcKLWogdUzTsMTu8lrS73ZKte
nL9+bApINEW45LbpInKuH8xofALRa6gttSnwYph1Jah8v/c6WATAy5WtM87Behp2zrQ7Q9CBebqJ
MY4WJiSxn4CerZLKiRFyj1JQezjBYq826JCNiGPozUHlXPGptXLSVyiSs8ejw7XDztAHSQfx020b
l/SYbdcryiY2l6S/K6dpzZOFMkWXuuc6PY8yutxrGC3Kqo12QevzQTWOrOa5O2KrolO6yfbFyL4I
IefxLV0Zjcx5z1AlRytEmdkBYdotZjT/HUPJRwqb3Wdkhfqd96rvK9Ctdaxg+D7rOwTDipDBN+lU
seXHYBmrOUIwKcwfAhqrZhtca5RZ9Uf14/lBaI64WbhQlPjgr2IRn/V+cwiduXLdhzxlK9Y3mPEq
uGVq+xUK0zEJPyCRGZHi0FFdmbu2WRA6OwY3kRLct3F3qO1Srg/qxOIM9iV0JAVpWSqfeGvDOzmq
xWpIfvrtgKZKPnwe8ZNFUvqgoB0NXurSSVXNUxVRXI/wpj8/KOZLitCr/Hn2VGKvkp8Zs2+95zqk
q9cEsAG0jbrYP3ij3LZEoLsm+sheHetuBle6ZIHhI+3SUEQHe/kloF/2mr0wpdnZfeGwuQ/iqcIS
YXlAutxKWMJdevs5rdpjjsm21TQjDnXSlKEFh6YeTV8GGJE8I9/YYYk01MqbtLWvDTBT5/Q5mUpx
OI6Az+wW2WK14+aNFWyIXzrbJHvOaJZVoiE4qCVYNN61ebb40zJH7C7Gsebs2s6tIoqYcsAi7vUL
rvEcyUHBb7t2LXoLHVDqHd4uGdyxUmMRQ7mqvse/bVj5izj/X2y46wM5t0trPx/HopvWPhtLJc/R
CDAvaw51MX6Blq2T4jjE6TjU6jiufjDOYhYSr5AxHVIimJsPIWVLixOpBv49oc9tff5nZmYFG5Zc
vkKHEFDVZIluBnER53oD3kiOkMJ/YFIHcQca72DW0J+JGmfYkfTwWfrtzRLGqK0rWahk7Wicf675
E9+utMNKccCQrnvVQpzPP78x9/+zWgBxtx8Ggp1492vGcd9awv+ynBxjETtaxClwHokBj9P6lyAV
RBr6EVl3MK/L5CGipg0DpeNyhgPrVw5tGGNGdPBGbWTKOM05HQYvSzm1z69TnDiIdBmJovg6Mrmn
+Ak0x9M8lCh878y2aRMRmW5I2JhUy1G1FpOAsaD++HgCtGSYCBWR89/3NfhcPXLiXplBtVP56WBz
mSOBfdbOAhSlzFEf9uc5A5x2BSoFnvmkj1juTmY236nRTibJu1Vt7f2rhfUVtEa+Q+gM9Hpnj6pm
wYHmLJP690f8o4yKoI7YyLBhh8Oy+OnW2MG1PlDRqi7ylw0CeKyPiQH/nkDg547gMHzanSeVT57I
2FcF8CdTtcDNMVrXzShZ6IqyFEK5/zBjm5SjUxa9/pcwm23getL9P3OAr0Fiz3bbx3fkpL7IWlV2
f5jhooOSH+qvET3F3WgyhnQpEGuwm32L2mXyxdkSQMrJjLyxc7b9qc83+ylH/Gj/WYZ/kfJDEehE
+O+I8UCAV72lJz9p12nJfkrd5Sd08drHLhj4Kc7rl6P9zgU8O0HnBKOEcvZy4nmoEIx1Yj6sHBWn
2tYuL7tyS5kkz9VfwSYpWstF0TTTORBbUcWLQ1gVMFzUEPGlrW2Sktm1BY6Wmyi0X5wu9+c6r4BG
ft7QoGOTiEu10ZIBI5zgtrQqGgrEIn/H+aQmF+IytgCF/gG7WPr2zxf5ZNJzcxwqq3SGSBl8B97C
jI/IuE5JTPWbWw10CdwcHcg2Fa2cmYAFmuv9L69gcUYn69SoOTdAjBogEtg1Mhp+DW6JwZzaIlSh
J+u9HZFtPHg3Xb7dM0wqaD9d8tvfyA4AN9yUv7elenhPhCHc5N/evn/mVd47mvfSvRYVghH6jJgF
JxGWr7M/Tz+6di/L8QriUBSJBIcc8Vs3muxy5rqGRIIRqprE9x4NJvxuvNxfDBxgiAaneg8x5upS
o6xui8zIpIMyqTbfIIIiHzksJOBSMBi1WtnZnec1Zf555nWEScXyULhK12sra50ktS6eIC2qOPLB
kmJz47PWfwDICMWxZcLtj+rQZNM8nwDJXv05rjh/qDTIqTaQAIH1LzRcscfVazOHeMWT9zzIeMdf
YjPjAXzZUFAsxQtMKAwXUoN/4ey1IzY+tqbweuchnBwsX0PTOaA4BCACGkyMlAkfz9xPwJdoxyvu
sm+ediATKEmIPlj8YG+CWE5B/b9b4gtdlpEXqnxgqapnK/UnL42unt6jJ0QJumFGOH6LAS2G9rHM
8qB3SoX8VMlV5XI+wdxa7J8SZqsA0lNcSg9ojzV3uPuojBMhTpQgmi8tZWolUvewzlUXBMAPU/is
DIDFVq1vKAyf3KkG0RbqUjn3OniLqiFFL2MJvTFxvdVjMG3eLAFGoRA88Sd0fVgIG3aDhqAufCqz
cKVZP9ISaEmRXj8B47RKmYMPHADXBIcw1q8VXqEligDdqPTDQ2PPqAmY1usi4SAmQgDqOu8RwGbv
jFfqAGty5adaPO3sFbyMPOCarEGMdKkSoiDkInDkAsf+MVld93ne46+uD/N3me7WnL7EhBYinqnb
/b5Lx+oH5AAjA4FzDOhg/VqFHqgzo67s//wUUd/b9L0OhAoCFBerE4xbZw+/jhiHsrYWBXNfWzzB
JKAMhLoutxudio5XkDIO53ovujq3472i9vZsB2d7MCIQOOT+ht5Cn33KR6xyVCN8KTEK1SckYJjH
MXHoV7ux2EWDuaqay7Pa8kz8LIWy3lGSLxPCmWPsqmvWm4oYvmt2B3GCW7cJ2XGiDTdpvom30dtl
gCb3xli2xLYr8pAwR1zX1KhSi1NzcxjogHpd8CnjKgJ2R48wq/y7exDd9wEP4Opo1c6qyK78BMXw
/ImtniZnrmDKuOfcKHUyHUP2eB6CJuzXPryMXs2LcNoQfmVqYsGTM+9TLgfcXxypHOcsc6rx3ubS
PoIzlPdpDrvjEX8hdbR6zX3V9Y99ngh7cRVJ9weBajVXDHnDa0Az/EGfYEsaIMLZc7sZAOy3JRq2
f7vvNwRo4d9MjjRvTOJaAdPdlavpEwQR7yX84iOqOeQaVVkKPufzlXm7lhpkzHtRrLBDttU1wZgu
HJKbjbN6crO5l3yCvbfij7yM55L0TLKOSMgTLeaRkfX4RLBUANVwcI/uhLX2ycg2s3JVwEcMIZs+
wh1hCW/t8nlODKTgokQ+7699FFF+DIGW88JaflihkbJ4bqOJZi4wzGNx4tG+IVQQ+2tovLbK7/7R
naPGGtDcoxO2d3CtaUkknBw4Lg9IQwXHicU/8/fFkuXKj1nWLFGy/DcgtUp+nWPHk+eGPk+5/WJl
igwVK+UKuVoIoes85yjX/cN70D/esBTPs1xxECTre8DUyN1+QJrl7oDdpd+jMfV6+2HVqEnnnbqT
kn1+PBanqn4cqIQ/YVFyXAxqoIokDpbhgEJXcGoukaMyCmih38SajK3S4qiq7z+OIXbVlBtNU4sU
pYOomv5ZO9iEduFlw3UB/YTMZb5k767MiLcbmGinSNbrxjJQ6A1J6yh9dcZqRsJF7y5Aikkttmzl
yycu/BbC8fqk9RrtT5mt9Ms/SeiFZnR+PZWz/hP5QwN+nJxLD3f4kkH9qcxYf9NyYaKqQzjTS5sY
6t8ehDuyx2PAiG2lyw3m4oJkDSW46+6jCsB82spZ9+ZV8J859P/hf2Ndb2n4GcKgZ5o7ZCPSYdGs
e/rlCRPOniwYtZqT4vo48YVfTgSeHW+d4BZ/oQHEqKTH89fL62S+WlO35/WsTqWs7UJzJQSRLjqE
PPkemRkrds81oRuYlLpyuq7xS/0nPxGJA/Lufhq6JxAFG8f/eGpjuh+pKoqsMvKqiBpkptiiWbER
NY7j5/dovl38g7lfObq/Mpl1d35aTZEfU0sLkisnkF9Cmf0ovLqKa863jYWzpbQgJWamhclsWit4
i9JOjbyLFAWlZXhOe9XxmH9EwUflL5Tntx5GwTfKzMOIyiK029iGaR2tSAOvMbvS0rMZTIL9FSgP
5hehKAvpgtBwfRxmxeDMEz8LhI2C5e88k70EsXmsODh3bsPxsBaA+OpWzS/y4Of4NYh4ZLTVKmSD
1+Qy/SfBXlzP7CFppCM6hpCvjM/2iBKg5zujxU4oPcQKQSOGtAFznU+ZSsqoU27ttgnOgMN0su4K
DtbkjGX00QYnxO6yYLi4rh5dvtVY3w2aZL7DyMk2g2qSvc6WPUkPGrW9JLg+nYdoZY3FDNhMVUwj
RMTBe+3zi/vorxDT0bOQCZgXpoydexZf6+IW0GRLkNEMGODJywWdi+PFFpCX6WGZAxOxbb7RMBrb
LjXrsbpk9ouJzYCyh1jJ1dKBIRKQ8MI0kDSIZyIrQ6kQCdhkPVkcRqhaXKplsSMm/2xdhoqdYYmd
F4jLDgqVLWc1Jg/DK17VXqNP5INhSCnV1skKd7kRtPUpNUayEgR4WSaGIi61jKYF9zrNeMSZOfR6
SihASsiTw+IjD45RMCmmAIw0eq6Y6Y7S8FgPqL/eTz+bUD4PGRUCGFFPtANLXzlySeA9eJZNEhFz
qkR5Zy1rHlpNmXQ/B3y2wwONW3IUUEXi+z6TAtB/UYNrZg22aUSEXzF8lKbrFHIuQ0VCk2qKw20o
Goplq65RR9e2+fSU9YV2yCvQNQKCXsKjNmG96AcxXYBCpi6NUBcjm2Z0Sf+LeXkgmzHWoP/FCGQm
4F0dKSVgNMbibaK15dr+jpj2VJvGe+r42GZ+7LXiFr8fD/1wAdu89b7NUoqTkuTXSGu1nQ+6y7C+
WlrqnF/9m+/cjpm0dnm8ZiYPzl/6DFBSurQPuPS57uZ0vcj1R9oZJtXa54BI3O3Y16VSPBEqPYyV
nxkjzIKS6uloEf0BmWz9AV9xe3+adFurGDJlvgmYDTRcWPg3m5N+LbIBLyRPHDPr0gv3zlvaCxac
XUL5z9Okb30A7kf/5PBA31M/RiU1lDrp3udGKuwPcHJHUQlToB+dx4vPx5L2/2wSRfh0x5MtraWT
AOFyZ8K90LViFynnhl7vCM7JJdL/QxCqKKX4s01soOa7ctlw2WN7Pd2bVPrzsm7N/VPv7Mnsr2hQ
07L/fQxn5zoOPPpoiabmn7BEQ/LxQm6+00R9M2YOV8jj0ziQCKwOPfu8KG8w4ecVyDp65MoCWwHJ
Kf/LqEjGaG/mGckxYclwqLUNd5tHFFHYLJogveysQlA88eSCbgHtbQrR9+r99/+eynsjhZVDgJiG
GpTewt0NRafdEEfKfhF59HScclDFGEOjQJqzLSVXHPJPWRslL0PsB14cleA0/V9yCN1RBKcM7CAQ
PBvXsYQ0ivxAOA27PibQ1B3lvkMrkmAXIcjISuX2hSsOpO1mY9FJSvrO9FOL5sbkWrmT9t7uYO8R
bhsMGC9pmtVk+Tl9DviIfV5M41guIn9sBwq9wMyX1GpIn+LfHT5o4ZsGPlYq2kD0q+cvSCth+leR
KI510g/84CakjUDiLYuATADCQB34HnXqOVIqP8dCNb7HG/1yMHeyF0hi8cKcApU/01wim3kBNcnO
0d44fIS4XDhSRSJFnbgEUuwF6l0NlNnOrwhsWxh0KPutnrKByMjsrc9zbX3eD22ZHCdsL4pFjo/b
gjxBf8xhDaU/e52yEykS2tA2VQSloeApKLcw9UK0K9LN9Jvd4e3tGhgwetbuDoWfDEiQUlBInm97
ZEdAUynFYn0krO3Q6RFcsPAloeWW8RJ+BMU1vsUUOZRKPFYFiMBOSz41XEeqveK9Oy/MbpU8pTIG
l/RnFrkTElAMtYLRWfbDZF+fJRsPe/8KlWmFdloL5LHqPj8HGNBnJKLcY7julw1+EMuZSCHG+Dc8
G2cpdrPJDKJygvkSm5Hu2pZPaE5MC+foswwaykHs8kw8oYFzHDzpSBQFONpuXFP8NcVDLY3MsZIl
chpJ/tX6ks5CcBPMk5o/H0U53W39oDFrofnXoxiEo480QReUPcordOtUvAv7UGTFTZmHDl3FMCzq
R/3DYhimQ2beds6rqS/zoY/mnpX2f95Iq3f9oKbpAPMAUZHqEn53sJr86MKwQodc3W470dxQWLR2
sHpHJOgmbISnEivL1tb0qp8md1Xbh7z1m760BBkr9YKn38us2X4mc9AtAc9uuExR0a5ShcH9Uvb0
mB5kY+vSfiXqFQZLymsRr1aBFzUB6mzS509LmSRRC765R9FmQOqzQjU9fCxs/YiiHIIA3U9RK4qH
0X8kIuiZWwi4kKPZdYkTvRn5ooJjRLJzwMdJBHu2bp4UbuNSN+EtWFpG3/QQwKKmYVAhqCumcUQm
HHWrPtDQ94MyEXPGjCdWyszim3+KWcy6do/zIA3SVJiIiSoYuf/2+03cFPWtNZCCtSw6iy+/eVXA
bhLjeafFogimay7FNfGLaEdO0juEEQRf1GN4ia3sS+q/L+dB/fGZJUKyQevPCD5LqaxeJOk2mz5z
oPmAniB46ux6u8jJ6y3ajkhJFhvmQHDujk7hM0qyW/3CDcR8BBoxmMkMVfQgslvrnE5uOFc7y0aG
cLA7JNXy+i6rXsSe6VlfxKHTSwbCu69GxvOYpwsvqH7mxph3NcHmvGCi+aS6vdzRg2nWRoFuwTHC
zZzlozWMpm0P9OdLPQ+RHrp4ltyJRHxBqAC0iYoBFLU0cCGEbY70IZyvn4uXMJJmq0UjdPDwhMJ/
HQHUmC/A4bOHGPFbJo+uJMyV7i35HS8s8+EdXqEWN9PBa2sIgc0Bbncopd6NR8Xh3aY7raQkIq0e
cwUwpYT2oou06fBb/S8g/I1S9d+CM90lQMU+NJM5p/gWpVnrPIfv6tepj0yp1TuF++24Yh3NlNN9
RjrBhAD/JBfRI/e/Zfr1ASG9tFek91yKXXio+ztKRYZJf750+nkZR+suaHK4AvOUqSB/B5Sm0Lvc
kczZFb+NyH0HnRlQMtkMbBbpjfOT/ClFFIpBzbu0W9zMmCas7HtO9UfX5gY+RLCq36jttD5+iskZ
i9TeOzmgT7VK8phGkp484agJTLsuA0R/ejvIxLYqtgIxAMivCQmU6LbyEehiYOMW+/5Fr8nNoNi/
7ORiwVMXB9RJ6oTaL8NbDSjzWPE4GYkyTcnlhq/2vYsr+fwdrF2V/W7hIRjZYVzemLTqO3NzGMHf
XGpZwSrVMWzxFtyczWiBb/in+LZGt5UIhzODpxRzqWKMWZroNeT4K6Vl/drV1kaSuFpe5EP0wFjb
FljEmeSYr6h/hseQZI6YvUqdtcsM2BKFVajwSKfgLFlj/a70sPluoKaw3ZiKCigfrDqKCpb3Cvyq
ND7fTVh6+C5hT+M4rat/gwYcL7UAhNd5ZsAm91P+Gx9YZ/UmYwMw+WZxRbg63RMIsPI9H5GqTTPG
hsikyTz8SuTRjq8rd8mSOGS2wFqzOB3zpegPNNszseUPV6zZ3IuxxiEu+U3StAb0VGYdczR2KG7/
C1lR8U/DgqqQhyXpZNYPiV8AtfvA2Qfg4Y90xGgXHOYD6aX4zjFfb19mBXWM/0ijy9xTP3MNab0E
kVdtqQJ4Cv4NAUITt4FMEFyqMsGoopG42moSgp0kAMtYdrHxNl2QL6SFEMT/3wH0gXb/zn2R9ZRX
hRJL0bDl4DN2DAJXybZoowhJ9r4eoNOqcRArGvZgoni44X/x8TYtkc10e3I/W33alTuhSvi+deZ4
v/bRP7nxLvesDNkTzN99+0k3JcGYyS6rWmBJ+pOWgWQzgDv3gVCM0+HEkeF+N+KA7CPIC8Gx7tIW
77D3fQfVvC+q+DggrF6lIkB05SEtVUB8LWxO6z1xTmRk+3023D38OcPt6iY2o71ti8YO7t1o4UiR
Fwf/A55WUwqyFSiNQPMSVZNB+mgeona2IXgr1ue8iPe11YUC7S2GSYDXheVOJoVdqStNKtRrQZcN
npsRK7p+Q16BqxIQjOJ5anW/EvqpizT+WhFaOfSRH0TqdFDo+KMbmSTqKMH6qNDVk88tltSQKb0g
w0Cy2B+9bh1x7HwlA/44k6oJhwrV6/MYZNe2kjElVY8RwoAlb2QK6Bm2kzvlEBd7liIob3IQqDSW
UtN3PnHsXzg9VrDeiLyqJf7TDNsLXm8DnvIBj8IS88GECi1QR7WGJCirxR3mlCvDMVm2XceqhYh5
rWyD+fENP2+AjgC4l7C6927r1DoSlqZnYYYsjGaPPEyfOhqpoJpoibq2OfUoshZn7fYAShKEpw2m
1yGWAVRw/YmsQLwls7PghkGt+1ADHqdQoTZWOYbrgoKRf0tGNw/qsRg8pp8iGSElKuzojtPSFtR/
6FryXEdZ4zbYgmPqLrttrH7fnLJLhrtAssShimHpkbQwdv4/abBuW8yt8dCunN/PKJ9N1rbHou2Y
lt/VYV12XmR6wLkLnWxV4Li+QD7uJNcheW0ZCVRMGOWHFL6BXD98bnOu13TaZDn9Uoy3l2DiTune
vI1I5bZX6AbCDwI1xZ3rLEEccezikGaIHn5yPo0MenceH/OKEG2xLT/qnm0WNweNUMgmJy+NUAgA
qlSGQ7tTiEU3RjL23vCekN87/VCqfBAgOk9sGuBzjPBynTlSr2ipDaaEWxixjiThFdwIuvJoYa4l
52CNEk9oPkkmV7WnTRZ3HNbzHzIUA0UYx+55fb1ut/no3tzo+J3neDOloVuOvgi2VxljRou7FfvK
a6rKRV6yhPHHxA7CKDMEL5/ciP3C0fBCUrpncHU0PzOJXJd9ojdIYZ0CroP8TYeDkuvSJ1NMQLNk
iK6gOLkCnDwDqdfGTfqgzsqKkNr9f+QlB20H2ZN+NdSD9zznZZIltA5LkP6YZR04O4vMslU22vNA
uqixlQ04qFVqZfzh1Hy00U84i0mMNRQLfPgupqKgvpCeeM9YiU0DItJSglB8hQAdCS8XW2C9mhk5
+t4dW25LtaGMEAlJOrWTyUxCkNXzp5i415LO/QqlZz/+3qvk3ajOUp/l9Jq7bVsuw5t6zb90NHbw
/kyPY9sz8lUkpEuJkW1CEz9s/rWVZYywE1auZwQP/q5sxZXZvtL54sMDnS8y1PdIAkzgz10R1uRS
20m3r2fdAmp5JgBGvlOMxGrR/skyAei3CrI26zxgCu4/4TAhBaoqgJNch1heEvhEPt2iqwp4Oe5J
6x0xh1sp922jbBRvof0/R21aoOR4UWguRd5Vp7cEt63LvkxH3GobM0gDShMDRnWEdHHfYrGBAtHa
ahAlmN60eO2h6iQwcWdMx35V9Xi/KMXGfFEVam+Kw9bzx4QdqvU7WA+I6Q4mPA39wL8hmkch9AZq
dvyAjkMYPfOpeR7Ik6A8A48q1DC4jRE8eIzXBk5PCinmnQDaPzO5jHwBhx8Wtn1zrmUDtBBWz5pK
cOewa97sD+mHOwNiRjG6rgtg2+O30pZmnFJ4BsNCJH8yxpUyaqrqOM5tEX2cijHlQC3shW+kVWQ8
dE3uVDoTNCkiMJCOc6IoWGAIC22uO5UM7ZFFtYbQXuD2BfaXwKPknpl50YcFtrfSaKsj1l/+aQdG
6mjtxSdWoTtWXuQndHaaezIcbliKx1mNojLOpv7Q+YRHqjmBfN4gn0YudF9RHrcft9nKGC/OiW2e
ATUMKN6kNNeIFoZ6YWrr5kADsBiI9f4+LWJFfSxxN6KWyj9S2k77x2AWbn1phNGVIphUl6924OEE
pIoYYsDp/SEQqV7gKyqx6J0FMUQG4OaPmEFLId1ZlDwJzHOgKN6BAxRbRCb0iJ+49rFHOs127sCG
8NC8vrpgmFU9drtCVOxVFCbPe671i+s51JDQsncLTHPXPfoWUg/UPcech9X8lICHwjNQnosMdljw
7r8+DBsibib5BMlwBsPXGpG9WOII67Fv+CFEfroLWGe9B46fQAZjeoCweeNmKoA1j2E7IeHZkST7
k9hUX5Ss/MJdF2b1Y0vSTadFuxYNCErEzDLPw2Fv6HW6kK9ik8DgO2leBob4k33YkeetMjP8Uu3U
V4ZcgWfXlHeBcl0/1SGACkmSeCNYtBdA1PSBeAsv6QOQlzk6qYR9vffy0gtcAQL1cVC7zmZ21kbZ
hWKDN5l9gpuFdUd2NB5nkShtAJeGtEeVHzrsFfvBQimxFDIalHJw+wHw9Qbqjdwv1BZim3BmpEJO
ikpa3/F26msxIcYNvo7Sscby8LvwiVzz8x2xDLj561G1wx9ZNuvPVqSK0oTEIyp5mZ7XPw51CP+L
qw7uvR7NKWtXvwsSAw1Fc6nIeFexJABR2C8LuNmxB0xPYBj79h75z22FAje2ffmdiCil5DntkYTq
bYkGAnyYddeBT5ks2JqbCLoenZdKE1PezxrJ8LqzbsqpZluPB13sDuJKDTFICN/lmQl2tun9tws9
M4yM0mzj1rqM9JdeH59LHxlKYSIfjLJtl/Y5EoqeLYAEAcv7U4QkGJ00RSOdvToS2oR8z5HGtOTY
A9oKJk7gUFZwTC0QtIFQeayqUogx9D6GV7eJahcZcXMdjjZyjCyULJbFb+zKf9i6LD7e271truYp
mmmsxIGSISsv73qgdOQCEfPuqHFdu6H/tHwnGXAt8+lZ0zJfu0xr3yNmT4x/y/p9FUOs6MYmL2Cf
Hyte6nmS4o+E6uOO6utMIaqXJhY57WhM+RunuGtjdneqnJ/hhDD/toVThVZC8JuZ7Ob9x1IsOWvG
WC7nYHdS5xntLNt/ILa2i4hJNhOe+OKMW83KnE2Kp2OwPuLaB1qeje1F1NABvk25hk1rqeuiU+7x
Z1iFFbDzPPTWjLs3GQ+5h6tPkkeoYz6x2ln1ATUP+sy0mHlGNtiB8AB6N9jT8jGFYXekewjWLF6k
6B3ukJ7Yf56t/twKR34ahMRBQV4erfiUi7q53UmWgYBwaMEvzRclGroAOMF7LU2Ho7JrLdAIdvsE
btdQKiHYazjkSeVsUjJEiLhXB6TdgxPBO/Xq29J3V+qqjMBYBqJUw/Ikj4K7KgebitGojqzOn5cW
JirB41n1wtagUd5vt4r+FPuRHMrlIQIFL6e4H1YjfpKdqK/bE4IG/IEyFWBcLrOvwTHaOOgqV9oy
n8rELMqnV1aCwBsEAk0reBGpl5hgY/qEUexzEGfKnhzcvmtM7yQ6YHGbF3KGMzajt4LYcyWQS4P3
marnjK8reSvCXwNq54j5TDxpW5F2m50T9eJCP81ga+2ZeW0PFSvYjCGP+ep53UStuMfAXV/06EAg
QHZlX2Yb8zm7bT9vOiMWvcDsI7KUNu87CFHKSzIwZZeoWN437dalS3MGTXxyOcJiu6HIqO++S6gW
Zi034GnCQKb55+uukO+mqBvD0q+d5zABmDCzZQGnJlHKDKLeAoNFAHIc66+Bh2J5AbCZcAX3CjPE
Si5K87wz2wMn5PEC6URld6qgtMJPpJu3qYMmL3HGn8/3ULmH68llXuHGcPA0wohBwP1VU6IqkRQx
aJJTDXY777/R1xMXU+dj3JtPvxoGRHlle7RAZLPEbj1068dORXxjz+ay5oKh//N+9oar0PnD1ZYM
UOkYR6mbLXHjY22O1SeZqBUuFzKG5RAmtn3YcsEMmVo5VagjvF3qkNmaq490hT7IUhdCysPuXqsa
um0EPc+6OQgphnOyCQ4NX3UQfc7gnAGXp6Hkq53tz+tgY6h6J6zcmT8SSS+1rRBe0L0fMEyt2grd
YCXwyo9mfRwV/JHK6042mgUCo8aGdcNL4xS+nNeeqs/ORVtLgGXia0rb4+x1LEScPWsq8LXjaIS4
U0AUXsCh+g8tuzWOOs69J8gnQ8BI3VGJag0eCa+2XSFua4ynTNRsogi64nnndfhQRDz5u6QyzU/l
yleO7C6Ma4iOoBTQilAM5JJO6JoBuclKmIQCh59aK+K/aGGxRySOG1sRpvov17KmvxW0z8m5p+qM
FacbvHF3S+UwYxj00IDcWDNIN5by7+sgI90WhmkrNFDx5NWUbZFCqPnyj8LMrOMgatWwqXxZgVNt
iuHd1nMbmCPc7PQPKRDGf06SSTAhWM2CdFOwISAkW47TNmB4SvYmTo8FmWBa1f4N16QFX6c2a8aD
IByO6siDy3X9SrXGjo7gbHQJRuxmjsY7DKLrk4BurDZi2yLQmILT3RsgLMHzCs/fDSmPYNOvLBw2
Vqpi5FI9deqjX+QN9uhTbpmckd/lk4wTCawyGf+yMsSGmErmzPdMM91P6f/vThlioWJEbq3TyL/7
lziBKjcg4MtbmFzS/U1xr/AEj/brZagkvzje6MpTBbbs56+WwbFi3lWwP15Eyc8kxz30+LFWnXly
vFgzcvjzjppRcA28ItJVk1Fa//Sn8wtTCuilauQpv4XR4dv6WVv1ViHgsnHyWXPGhs7RxyBRaS+m
vInKQcX9pNdShaeoW9muaUnweN/IBxqGkti7YfXXStOTCq5Vbwi9Y5HvMQe6nuj0JniZFQX+Modw
dvVTvpbefO6P751i3bsQobGfI4bm/0/yA1gp0y9W+0v7j8gN/RIKGHFnx11bxXZmsFHdlxy61EIZ
LilWmTgoN6TXKwQrnjFhgNUEAARkI5Yu+1mcd/srMzEhmPt/KjONXTd7OgF5Zc5U1o2wZ6Q8LgzG
yUvaLHtJPTNVjiCcR+YnOG0k4WMAC2V1ICvcXzAcx9d7m+q2tVVCZiWcAcH22HgNDkqVhF6giYBy
T6iIj+XOcreu3Zs/5mbWLlQW+PSNkp0mfIurTtmwQkJdCGW+1r34JT00WcixCVPUHpicnf9AxStx
ZlorRErOBnFh0k9pTXEdNJr8P9xE5k/+n2veke+cOm8/APNjeq3A3I/WFr2jvthINmPFfscBe2y+
ACZYWjQHwPRbBA9+kXHjIbs0OeEbUV1laACPaE2Jeucrfm/0mfeAfe+BxhRVheaw99SytGya0eBz
HhxxokEA/ZF8+hzzHiZ7qC36LOo1JgYy/JtVmhHLbsBdnvecd5znH509jZtIZL44vxgu7iXzqjBM
FCnXKsGWzAat1yZcCC6o79qvw4GX1z+JkpPHJO9ILsSev0ngx3rg/fnxJseepWwexrIypS3Xucr2
IWGQHU1Vc/idbgxJt9kwNytKCqrh6YNFAs8Cj68t5mgJgXGSPVXS9uA61DN1mz09LHEiDcnRJfC6
8QvN9LF7U2jPSLSOCrkjwU3pBCrI8ZmFbUr+5g9lhUdh4tcIbv+urvc/U4eUPLF6rns0syNs0csA
mvgNpEBUkaQGfrFuwfqOvrCjtnvHRZln4pt0kFO9FrtddWpkHJPu+7ahyyMNrZPmz6eOBYEVfLyM
h60G+sLX8Y/ZkNe/wSNvqch3+ZD0HdGTtnHI24dZK8CArJ2Z6qSNcQkKXN468VVYEwsSl7NWgX9r
OsZpQb9c8Y6bfGaGexFIhB1zAngsNefKoE+y3DhwRVDBW2mU8cljTFeU87jIhZRRNRZpI8bCaUvj
4xz2FsUpzz8M7vlD0/tgBhYBZ6jnBRP+iIAnq8QkMEW7lIOUSXpB8tOGij5hu5zVKHA73xxeFRhA
SYrRMaW2snR5OiPrpOldsNkrOb6ai1CYNfM7oGHy4UmpaDS4KHOlWG8Xqb2pxS96LNEYeTigoqk+
P5vqT6eMSk1ptJfTtAPiOxajvHTVBDDWMi5W5JH66JvmXora3qk5KGKWszJqjypeqaclHB3EsrJt
bpVcjOD5ytbR6wInchbVL8M40IggPG10nbQfhGuALPPdyeoswx9g58I5rnMO2fpwiUntRT2Etkrb
RW7Zq5Cd4EqlzU0ulXVyFv2FGtmt2g/QnUDNe0rtZqJbMks/yKhHegRr7KQ1+2xn4oabZ4IxJam4
xDhddmnr9pRFW/iipYdXiZZ1LBIWmBOi//PV2O0NL0TXm56WSa0fe8aWDG7Pg9W29uYGzoaatllK
0eliJGUGnvc4xKe/dt0D81xtLoVs0dztX70gqaVI/U39eRfx/U3IvrX+R+HgC+Y1/Nh3SzLNfFs1
4hmbiPJQV7sWVjXDO8C4UDZdJs0QfIHbjqWhzxYvQjJl4SxqcUo3DOAxZkFEZDOZeAMOENSc2CC8
KJdAfYKvnLiMgKR0Q1eReTqobQrEQp5VUsrPkW7DWkSt9M7aPjgQpu8hVn7nlcR2nroCzOBl7sRS
FlyUGYHH4ZfSUKczp94m+2BZpxe4fpbHBOpRCd5qu+wXY9kb6fGehVlLWL6gxV5Uu+6ipJtRzoPC
y4KMoaYf6NaT//dlyWpItBZDo09ZXk4R96FbxpJgqVuxZKFTjFVYfr683P/vaXbvjUOzIn4mWydl
PMDrn3UhhghKsCNY53m4tPJPoisnU/d2xrvCG0j6G4k2M1sr47UizwfOwkj4V/SeYpEFgMscn6bd
UZ/Zb7S4ODNp8IQ9EuH/HULpQ/9MaDNW4OEYJG55WsVNYIfy5BNKctTypDjqKhdEfYPnJQ1Ct3NY
7WIF2Qf7ymq4yX1yenCSRgJ/tWsxbdokCKlIV18/5r6iBUaBQm/EAPt0OigJpjpYhBIewF3Bqi2z
ItU1l9OoXOJGp9o9oD2cDR0DS60qJLzzvoG6pO2iiTDghIO+NOCchS/dy2pKKHzWa+gtcD+OVNSP
1EZZPsBl2nYJ+qJPan6EeXfgE2X8v74UaEvkxEbkHhPp4TioP+nO2bVml2+479XoSxBDx4Za+3SB
iiHblmJNa3LCzT6G/75kpRk3Mf2T1npjds/NUePN1avMlZmtwfnFy24W0l7/RmPSu2QI7RAxn8bg
6FI382Yl+SLSQDBzPkOiWbvJBCr62u41mNiGFIKYE079ovJam7VgGdwgTEGoR9FFZZwpda9zesZN
3XfoQPEJEm5y07R7O/q2ZQMmb+YEc5jAcR4a9nUQnWtf1i2bPwbz+qFK6CCpIOE6N6bi73wOHtiA
CJfALBWKmfWz4nm09ICK+DVMJd90/+9EzJhOUSL5lZWgd2c3683weG//ymls/Bt/+gyzF9kDWuuE
q2VnajOZaVIRiIcp1K/zZ0iakNZwvyltt33REWqfFWmkbnIhc2wH39Cqlca4QNr0emOLmin1+hhE
tnntBGLFp1yg8A/yAjAq1dMaG7IUKGiLiWtBubG5YKeFs0SyGxD+OGXIdLoGGqTJqiXFH/oxDfJx
MdWXQOH7GVwyorrEl7hv5cbJE4SnSkCtg1Dk8bxGc+MnypR4pjg9VO//FSuzT5FXnxoTiaHCrqQA
p3/7uNrTV6w+5ZLBe/Eo3uM/DfJZnJNP0fbbRwT4AThN/xmE/Q7TaBKZgAABQCBKdQHaYhCQXBt9
KkDEQqZ5RRebqRpg194ynkhgTSs9JOK2tjWmsV+LnC29sxsEK8VbEZW8vzZxyuCtbglbKMgiL7EE
JSbKtoNpJKa9aEVOQ8LProuqrUTB5YkjChas5AaZnz0sZKw2yauJTH97xOSTDQPwvQdXspwtud9l
8uci1tj9m8qWScrgXrAemvlwNZE5rirW1gk1qvT7pNKR89zGKS6MGVwNYKwwj6Pe9LvtPLflhcA7
WyoX6SX/pr3uFmmLiyLkvH+/TagoH3F7hxE/X91eZRPoUaR83O4p8lc33pYrfzLHTIeaezqWYQop
DMIwEq5CP504YP/dVH0dpGmi0pXJQuqDCJFMoQibUdBSCZgyn580yRm9iieMrBP+Ioi7k8g39feO
YMVzatCyiDF6Pf2/Xi/Cq0GmfqDwENoRqnNrdeUFRj4mc484pOtKmIrK23RdydVNTzsJ9wPcdvV4
zEoDQZyzv8sHdVeugd2jg718/agpt2x1DX6L0P5PatBbnaKveg5m5ur2a5xCad++owds9UnqN7yc
CRwZl91AbzAtNabhJrlp4TGXQL9nudvthjq3dagXBkWkNLyzIleaTHh+kK1V53oFZq/Crgwo9vLA
MPoEBBytZxdVib08Oslfpr7UQ2qlZh5ftD8hCYT+tKpHoWVAceWmVdkFMdNQlxNlBwhT8Z52Ec20
So138NtKhgh323bzygtVNtGuauktH1JPKw+yEepCYVra4EmsJktmo8UbGFJBhHHJs2JvQYT7MNTM
JL0iS80qzJ0oGoHIK3q3xQ/n5ZPoboW4FK2NiItygMIWq3ylHlNdkSgbr8TBLZ6PBshMFNO6C2mA
NRgc44HpMkp3VuiX7znBIehJHZPOpQRk0xu6hLJ0Maj3ShU1+cgua2T+Pw505Aw02YBsQUnuu3D+
5hZiaJ5u8x8v3tia+IcZjOKyFPvSwsT3dwfxwKQZCA4FaWTe2eQy+Z5K6oB6tUq/1tsm5VJASusV
kJVyh+8d8tk7LXVQpiCTMM/jR6qAH2+3yAN0KKs+7AnTmZkc5ccgujHCA5gKb7BOC0e7yyyVul9R
i5SmWXbqXmmeidKZfsoD3PZIdY+RbNzo7JQJtoH9kvLp64UAaUja+nLLXqpSkHSir5HHKxCxRfiA
3Xu5dRLNjllYkoYlARb6micjVxJg3Bg+uj9Jg6r/ZxCHnkljWNQdY4mEHps2Lxt5rTj7g6a7SPbv
3sxduxEnzjAjPVk06EJQJwNWRJOmKHrodxk1U7hsSNtIRdw8bzL8z4aJZ2q8UvgRuf/tStJDN429
zytsiGRX3MQBBB0VDTgLcGdzkhDTRh6X8UjDtw5lQp6izjoSdtU7Ip8n+qxRqiN1YJBHyG5e87/L
HDrETRURwWY9PMvMvdkKobKab8KM93D+pBA9II63KI8qDr9xuJ6GzXvMWKZdmg/Jqj0sRP/brsDK
t3+kHRCju4ds++cF68IrbE6FkE3x2cdtqXdDPGURdAG+snJl7HUNmnmRCT9sQ4tdH2qNxtgJAAia
/1Gpw7VqFIxtxo9pUCK1/6anNGWJRYEigMWPhLYq5OqMePy4r379wYBpLBt54YQhcqi5NEabSzAP
q0xh0NnJXEsS7Vdr6EW8IC7Q0CcScH3xAMOYaFSltvrTMtPj2RthrZKXZFF2wNoxp6joUiiGR1IS
4qOqiLkKmIa3l0tpufmalBk5t04YJzhU40oC502J14aKPnsInAu6r11yq7VF72JhBd0pzNsyuRlI
1AyduubkaYfI75XEVGbEFPPdPS4Jw9TjWvwHRAvcj8Sljmi0GgUYnvFYJ2y/e50zJoYmGI72rBqW
/AoT4t7oIGXEkSxByp6UHEMiCjZnrPHACkl67mRJSBOzHsqdwSLuY9L9z7T/GsH8nqvtD4mg8aUI
c0mKyzibu6Qg4yliZsuzdlZIqInKpbMWiFjbYdoQfTvc/iSBpHrHAIXUM1mOKOy7YOBYoBZd51/X
E91vqg7Zx0cYCnGGJ8cWZprAKJsdEM1SuMHmK2g8/RGamwePwKScUgcDuB+n0E0hOJEgHTEisx0g
g0tA8Ifp2Y/JZs9VbbWhXieA1ychrKeMi4RMnGnf7kPNFhN5adoyOXciT9WO55lO3Navck4piGDs
0ubrFOc/VSo8WjDGllBBNZIO2vaJo6Ebx65fAMKfUezSZTHt0Nah/ILe1z/Ha6Nq7W6Mn3WVdrPd
BbKz/MorvI3E24aLLiXID8Bd/vpjEPA5nwY98uWiMQ3hWghlxVSD3kNWoNwAqSt3qVGju4wHBDqi
8fTvAx53bUmeu8792j4IAi015yN72EUI2zUINlYaM11Jw81a1YyYa8ZG6ztgiSXpZw0lA3YeBU4z
2CPYbhEm31D4eDZWFfsZEzzC7ErDCOfVMCAf7X1iAYvMchJMU5efAVvzgI15CsrA59rZiKgaBOwi
7fcEIEBTEEBzjX8pDbDs7J2NvoWhZe9SDQ9yYV7mSPnfySD3UrKt9DMjcDOJ54IxrAOuOmn85IVV
Sc+Z1quu3qIDwFiqpNK/POYXbWCa8Tj6G0yRFqTxOC8Ct40TdgzjHqlAhhdMCxjWQ18RF/WXV+19
tNqftnFa0UwdO/Q80vSbOlP+frEeVdxmkm1BRfwr+oiOLd39vPVFQEi40HX/Xwwtgj0MtGn7E2XI
SW1OS3fnxE/3kR30UnRcVdzHymkn7Qhk/tllw7NWlWBRjD25PtV2360v9XqmF+L9+r16VD5doclc
37RAdjjMg7Q8mxYv+kjlOytdaqPcSeazqIUrsSD+gmOWPnxDDo5ezxiXMK0BfuFuw8e6u7KvhA6F
Cys43kbm+2uNIMI5ke5q78uCFYW4kP3SqqC02PaejOwDgbx2DWQi3ZI1NG6RLU8cL8tXvjo+C1o0
FOnjPxWQrW7p+murr7Hq1QVtBWIjr9oMbsR/Zux6/HoqgC+rt7vxFr0BhxfnNGuQUV81YOHKGKD6
i7FDxAAwZNPG+g+o8icBASpWMRGnRF21Di7feNcb3F8L4q9B3YScGGp9EsI0ZmiViLznIlKxMOFa
pEdud/hOjpQ+yYCVJ7+dkuYzTQNR6w6vydL/04zQIjvh4SxWMa2uTRzLyldRW4EbT89HMd5ZAYdv
ejY/7v5tX8z7cIGd910MW+GnKYw+wNhi9HGKitNsOd++3qvHoAynYW1JoXBQoYE4k6ZYRItmWk1D
iIQ5Cv+vz434orZazTCmWn+2xOR05CcwwCHfcVm5bwk9YYKmts8d1yv7npVjS8GtYYHPcSQh9Bxi
ww6NAZbLkjtnkEPlmz3w5jFaM1NeLuIo22cK8Fc8Mge4BhtvoGASU7xoZovM0B47mQqGcUbOoUl7
p8CQKiL3VKMJ4STDDPYvZUMDy5zg9oQ5jkewriVKFX228GhPHsqBJIkiZur0yr52Rbx9TevNhEL3
FE8271bTmtpPUCb9uW6tbg0uiqLT6XyipeNvF6oKH8nS1ntx5Bd/uWN9NU8kFWXLMBLFv4eJlSGt
TxXqh68iVGPmJ5r5OHzC5fgI6Yv6tw1d7QIBa398RtWNbmTW0fiQqx1KktlozHFG0ZwF/tMMDyfJ
JkozaEAgs0JC2iFuRZnvSgrKqyWTb9/baDtF/jipzCEjk+n/MHFz690xllwLGTw3z+/Wt+gNC2Q+
tNpdeqZRFV9CJU8Kvwh/Z8mHDFPgl/gmy/Ta6z/IhjHIuY8MJtuHHpoY2U25hQiAdZG42W36+8KQ
uHr0s0Yow8kwpoCIsbVnFCwCk7PhYlG434pFUuo9FewKjzF9X3Svgc2NabLGso7xw8vYlHqhc+w7
n4gD6Yv/32DwOidHSmv0UdV1bYru+S7bLkWhXAq+6SJNyvHLjYI2mANZDyKhJj6pZPNRYrxDGbkW
JobfsKwQptmjkkZhXRAiW1t+MdvEnvz1f0zsmxxriW/qv1D3Bz40gM3qW1pLcop5EVFOEq7OoW4a
oiVFfhKfeJVbc+rXWrC/hGkbg2csPFLw0SAVNgdLht5HE1X8lmRq+lY2hKMfu15HihQNy65Qd7W+
ziNLO8DAX9DI4Qh2RbN5sH2G6Ae2jy9A4vkbgX3Dv2/Tj74mCFuX1rScetr1qwAzDcPANQuJ3Hj3
6pgRDn0RJ8sIknY6rbd2EIrkHMPKS7ME1RS7uy7gTJkQz0CgDArxkrQ3Euo+184OkDzaMHKbM2LQ
4crgKch1JtDMKGKj2BfTkQZQFt8StWHSUV6+bM9DQpUxaaNnLSJjQ+m15jE9LhB5pF8NaujQwPZW
IP3o2ymILz1PGDuFOoTJqphnz9dA+/Eujzb3n1fjUHYEC5qDqdHg5ui2GJVfawwls7z+oNdKjwAk
fqOScUESo7Tt2SvcpMOIeFYexuevg46Lqj1JDbA9daG3QAEFdVd1sKaj99Gu0xm7ir+x1pKEdM/C
dK2ADRpb40KaCmRtb6dV7d/NihrenTG0Wb7kOAc89ft3JgNJw2CQIt9WSSBuTZEyOuNpE9lCJ4S9
fjPQE1EKc6ZAan3ljAMj9yjkNSnbTMyIdNoL3EUzuS5uIJw2Ra6PVECgVDVmfToG+fkKR6xvwy4K
YCJrhKHMEdfCcaTwjJCgQ06IviiM4WsGV49JhILNStpmpAh5MMiwLfZDX32HH4reeChwUNsKeaoc
SoztG942NqkREtHVvCiD2WW7C0RkjXekroG3UNwv4C0ZIdiNcrp4mxp2FumebIVw3Rzsv48VAL7N
4AnSOB5Psrrci/pfRWO/WxxFr0nxBoWUxAHzHIJ/oRrDhj5UKH1I7pvSE2r9qqJZLl6kHPaQIBIS
qFzKK/wmZ4WcTNTU+lkzAbwERZzvjcYAhtpH8xKWy0U2tcDphzOQtohCBubvvw+mIJdHDhCJQ3tk
BuVNUrU9ELdEgRy8NMOGrRUeTQRnrZ9kecowxgwIjJv1po3Yg2ZgaU4HbbBPuS54WfmjP8GQnL8Z
ePddWrc839AUOl6hgRurY2XuznW1/Ga4U8ZqEBOW0CEVx61GrNGXa1zLPIbsdvKz1nnWHVWna6VD
SL9HUgIfBil6ELEAMtFBabpTpYvUNxywmVcsM1McosucXS8mgKPkn2Jrh0O0nv+DqNElz5UMKM6i
bCYrkKSeadb76yaIoTjCxnrv4qWUKm8fa7WARHwv5uBfiEx+HqcGzu8CznppKztBVqn8gdAKfjCZ
VP3c0qYjUCrE9+3qb/regCcUexl3y3OwHjHP7IEdxLoj5JpWLOu0Fk5nVF5ijK0sKXJraTIohTP4
IGGcCAOZYlLmathGxWlxbu6YD9uyY7mD8zxNDOoVsdreaOHg+nr4qg8yDThX4P1Mxg85YLTo6is9
UsTjARUrT3i0XMcMtCG9MxIkVLFrXBhT1nLLiWBUBqfPMF+LkmNGMr52EfUY4YLih+phcBoLOlpv
wkJbeORgWxrVvt7A31vgIBeD7eVfNUgbP2e++ovxUIUVfRf43K8SWiPviyAvotsPla3Jp5TSFGsV
pWPNKULpalE5xflZKdb3Va8J9OYut0ylfZDMP5X+x2I03bT0R9iQNh2hRYZ6tEBobCLT3TvMDT1Q
oR6QmfU9vlV/mDyEDqL6THL5AlGPe+iyk37XJV7o/RPxrEn56NvY6P4RosKe2FnhGdUo/63e6EoV
0qumoYhrxGK2maQsyrN4XJp61GKVRyrUo2H9Bv9c6ccFGsSkoJdJchentLwpHO3wqg3I7YBibzFh
0gShhl1KgT58JPjvK39KtJtcVKfEYkYlTZvQVRaHY70LsupnBZPNPWLzofCRRkFK5q/tPqn5pSGY
6Oalx3JAjtWnUEw7JD0MLNBmx14aLY/vjUN0dYsb4q5BWw8asgHRmecRdTDz74T8ly7YUIG9bdcX
1cyODZhQZW4AqeFZmEAojdx1TG1zup8GzLnwEPxVqo1m0Yoprc3FPvIkY9KrrpWtSDbbTQ1PAV6z
S69jv4j0eKrBIXZmVGF8I53WRqQZgyS7Am/IsRlf0oqdtE4vGU9ENUeEOL1atjH5zhEqeRL+P7MQ
RrN4MoYBhUmza32HRwKljRAjzgvjpBLVHauGnjr24XH2gDjQ4f1V3TftPaJi8rC/lgU3kAJvUOPg
17o+FyXPZi7uYJKFabPkZ8mgXsiwM1QPsvR54iMN50r2TqLyKTcAMDAxRzsLLNgrLj1rsdK+rPIy
ALGBPXRWlUbSOIzSd3tvn9Au6wF7hTk/6ezDLiemKfCdvDeXmrcaU7mjVAfg32SP3Z1K5Y1xzQvM
9YxZ+YQcvvyiEDL2opb/x2dzuDGL7isdCjs0ZdyWXfkTEcMaigIhNdwkUlpCnk2r1Ek5PpYO9fJN
XWQD3ROzv2JtK83y/0NvtnBNTCPgVni6FOD6rwuQAJrtX/7a+tvZvJ9k2T3VdP1t2JLdkW74YG1/
Igal2pt9ARlQvBEbxueyjXSZ5Yzsdhkg8mQdnSD7+riRfYx4Kq8kRNhPf8G+8P8ybTTu1maoOz3r
5NvP6NQxVctQAyTcvgQU19LG38iRLU1TKBgQ/H1VDp5y6yzZ5CK6Yz2X/21D6XPGHs3d4d71YuIN
5zcIVK90Bn/JH9rG5WvRt6Ndse2HKW1PBv2K1Pw6M2qUONH/sWNndKxQxCpYAwuyNvUTINjTybHb
LGjYN7sbW+U5VsOJXosLtG1+BmAaeaJW3tUPDGTI4jrV254qfjczsex6F1PcLpaznFRDupgOL8xH
KjrlwUeEdb6wrzbJZa38jexMQiVRxVXs66z61VXwJhE4FWsXeWNl7sOff5WaER76yksv0BVi42gN
RRNL/UZlr+eo79p6e55R6ljzLkF+t3aJlIokCgkDHdJuPhpNwkn2ObIQyeNIaIFFlgB8neIev19g
elxcwW9XvwTpNMDiF0TWZPeF4PK/uypxB4E0zr/3TvBlxW5f9dSdHXZcHagFwLZri1mVOnBbrCyL
qkPhRlnK9qvMPeSKsFlUhoe8TKwgbDwJwFohnFB+mdMzHa6wBgEfrP1IvfLpgSmi+CmCAUp/cXYu
pP/hFcxJ4Bi0ylT8xlGGX6dmJ3AZY8iPTGlxAA84HdRqBP9+m/V2YXrauKKbIsN2G+HGchvFjfBY
rLsMe/GAXlwH95WTrGr1yV+yp6AFTVUtE3XwxDAmnUxbcb16J0MFr9Wzb5EsEvhhNqPAdK7v+379
Bv1ZA60LeejRXSGxl8l/5SuTzpPQuzv0mdehYTEgPuQGUUdYGYlh0xbiTyW3bUNjQvh9WV5+Tx51
YXeUcY5Uxr5W9CwiUOmq2LwZegd55+w+PeU0SvyZltmn6OP3d1aLo6TTknc1yGBnwbEdohj/NwdH
SRgcIG/ffxjrDEYlUmWQw94XfzzqSTQfgevjkoFoOYQDORHThmEjqAQivEqe13e0v3AX4hglCNSo
6nK3cel33SO9trGQmoGrVs6S/S+DnyErm6FgkIKLJgpwFjrncnLow0AEQP+uf/772VyiF+F4nMgF
UXhYv0zti3CSkFVP2f58B2CcoutNpXMELVR72MB+YJzH+EzLqftbDGVIyk5E4L+ID1qSYovd0w+y
dEXXmJRMhaPs+dgbmORtnTRBGULlDS+D/dhXBLHVy+yjaP9VIzsQ/RUjln32iDOq0iJbW0VfmaBz
6V7aHjqiqLg6V/R5BEeOvRpfnltsHw3ytvMxXm9hVJNrx3fYDzD2+8zn8AhXdq+fHHnxe/UMaG8O
C1MBRk43u9Nd8d6kM51N/sMOZ5/B7o3ly0zy6wgK0KOBggIRD8dR5qvPeA/lQy0sIrpksaz+8Kfm
SnCc6fVwlm6NiyGYpnAUTNesh4DVmHXIqE4hFQQyamog0IDb7oMIi+EGbnUOJgCLyHKTJMhXXTSx
tsnjDqfV+xXL+tCC0lYT3xKhkredQT4VPkw4ruu4FTjDlVTcFJQg4gdS0uhvvPIDaxyowqWvOGXb
INcIiUO2dN4WK6foMt86N/jl3ZQwy7mb4B1x8LDh2QVYe/DtoJOZ5kFWfXCJRxPfIAU2kE2vk+Uj
yESj3lEwxPLTS+r/9wTW3KwrCxINKv5n5fnGTTO0Gs6zX4JMmWl74KOYyRQMJ1VdXsnTO9uGZwNe
VqAvVKkfEjgjdpeeDcBOsWQlpm1b7+Zfg5jSvBbtzsNTtIUu4t9M9HuiPMRt0rwMFX0f/Z7oc4WS
RSrZ4SYdi9Bg6Jr+CkkfW/WOgp/Jmnefvg8GPXCabsGEGKNdPMzPdS62WFL1ZIpD2aGqKFrdak8i
yW4eG/mfe8F4eCdNu2bQnvCMAGcKMkRf+UXT2/GskXT5Rgswcpoe6nFNKdiO9a+zr2T7rGa9ooN9
6rP3daxlFbRovSqn+H91fGwplfoc7fQazQp7eoLYDmEYFda8CbiMYV2wa1VKPhnoG7/IgJxsg9GL
00kJ00NPaeUvcJ5PoxLaME/vtDunP/9ElFr0aG2rFYbCydyPXq1/3UJcVYFGHR3PgJOtEBw0P6KP
z2Qs7M2+JARwiSnXCI+AuROZZr+JUV8gMrvL8INGSuPUBifIwSGz8xhEYiTVwRdxaicyxoI35fDu
1CA5ENWAJ9eW+z2mzP5PoASqFZCNg0CxBp0yepWxTJWTGvzGFBkpdWp+WernjrHifEQJ9trWo1KU
hWy25Uw3rJOpZev19f7h/sWsQ7h7IR8Uc97lD/J/thQouecxwi6eo/WIfYbLg8s0AoPLBFLWuEgB
jThlh9+IMRwy4B52DqPJwcQh9mw5w9tIVvWzxaKD0sZ7i8CDBOaWcbAcDr8WT+tyXFvmkLnCSkWF
pADivRyYo+7Mk4tY0Neik032aAIN7130tOQdAw1rwG2lwfTgfP/52jKFezRrey+3jsEvW0WgZ7Fc
k7/0EtuJlLCuoIRAGfui0QqxYf4vuC3TvOkwh8mgEN68vH5wWsY5CEeCPxTwtoYfBtB84eTnz/Ot
FvKF9gbv0I50TLm6G7sZdeVPx5TdCPdNUeGDAbzV1caZTPcBoLQw1ipJ4ke5dGR4Pa0UWsBhIO4B
3Ooif2fv5pKF1ZETUMe3SvAuOlRhqgWA6buqUolVi09AaH26sWZIdioGTp3JWMsGlpQiI+h+vDif
dMyy6wSC2wRwx1FQ6TcjurArDuEDRm2C91bi/M+vbditRMKv3vpQkBLuUXIiO6/reY2KIHnacJWq
bt0nEjf/zVSTJTDMR+xlfjaAUjeiqNLNHAGmdLETG1DjUqgXLknV24FodloHgXOyxfjYEjZl50Ol
U+6Hl8efypq+lXTG7jouJxHUweHH3JSUkzyT/m7HYwMotJCtCQcZjwI3B8PPU0KEDlDmGFKrQ1Jz
3dz6vSjVvrJnPRJk8/23V/dEVDDm2MI1MoIrzxMu7uQkW8EICUKM2nnqYQ46YyGLleB7i77IVJbr
uOK8HRwkX/+KvIQq5DE5z5mzL7O/4iYvL3xzLb/P9pEyeUOKgkcEE3AkwJEsfg04x6gRyt0Vn9Ed
2Yq/F4DgZX9O2PA15CmRLa5LdEdusA5Diirs9O6laXKOaJmsVAGHIJA1n+Or+QijX3/O5+DGvDPA
ZhzaPW32qcAVY8cFS+A+nia1tPMKyLJdn+x7rFzFdEGRJVaM3L8dM0pXvW0EW4TLsjVLEG/NtEBK
RWssecB7VBwwXqsY78qZc7ovOJZ2O9mPv8UTcfRCjsw1/vWgSty9POqNxmeoa7yv+v8FYHAfZNSQ
AaxPrdpd3tizsxkwmbo4ELPQ16NO0YVFHl8jjkF1rdx+scdt83ovjIPA53MASSQ4uomyTM88z096
mwU6p+s42TdYLprxeurcibKsNgmeTu5DsCbSIkHOgL3zcEEwwZN5XBfwlq/+nmSfYUxm7XyKlFdV
JWH+YCGw47ULn73XB3FaV5tsbHXlm095uPicdpTlztp2+91m23NHgR8bsnXVSAnYkNG4lBPB+om6
yAF2+8no0HfIpUacmxM0V9uTV8fknU5A7qnDw72OzFYefCRG6rYbeehetot+fra2mnsOoZYSb+AX
dlhCAvGJV6fhk81di8LyizCgOZhCfBBnKtfwaGcgTr+njl4EwXi8fjMzB8zHYnQ5A73iwtUtKMGK
pRBuPQKeZ/J0pRsWXgAF2cDJ7IkCbTQvjhYPNoEnhSvdQv/wnHESeuyNOpx1M1Aob/R9pk587G2h
cRt5Tm88VoimPPxstKMTX5/OmjAeyzRU+EsUYx55ACrJN64wDjFg3mcLfgWFinvk48X3RlGzHdNU
Rf3MJWNcqb3wnuxgVoNn5/eGuxj+T6Dzw6oOcXUN46HGVCX+E6pHeH4d3HVr69rGh4aYEJVHSA0S
idnHndRhwzZevtX56ZNdWlHGafcrs3Cg52e+Vc4QuSdMPb7PGtaq2rJFSItKilEcYpxBO06TPTNF
xQDn2TGGSl0Q45hgbzF4sjGhSQXSI0ymzXLrBYH8k1EElMJw5KcjfADZmjPvQIeNmFIfqfzt75WE
BDRZg2I03yszhtndmnbiO53Tvj67Af0pi5E7tAjcu50u3lC63PIsxm0p0OPOCBuHMJPvYG6piUBO
fYCWhpT+t9MWV5D/EohxGzSGkO+fTjfzVUO4QkPUI7KBYSEaGYM26b6+SYT8pnHZO+nTyGP3ZZ5N
kecH6/h/srBa28IgmS+mqmMS534XPDqn8cdKl1FKpRVeRFFHGyqEU7gkD5dAjiGYAcufzbm5OqIr
0qaeGOdz7BwFR5k27Lh00mBmVCGbANYB2ZQimYsy3OxNbfr/bv8Pa2+ZFx3g5XLRU/c/MHeWws6u
noyjWiSmEvvaFubKNn9JCxrRNAd9sDGdoJH8aPUuyJa9mi+wTcuq8J2l0jumeru5gz2INkVxKh0g
nenaYKZmLTb2aTh23nRTa3uZsRx2l2qZ68SY7kFvQTbazpSBYnsFJtUL2WuvPEs9w4JM27mWZvS6
00BgyVnaxdQMVCoCtvxX/IIe7GMev8IGuQK798ZgCIMr8XbYgA9/YuIEH1SCCe7mPFreBLb6ZWWX
GsCardXc74v6gw85OpN8/MvD/rNtFfiet/47dOs+JJzPkNp9RZOCdPPXtNsC2boGp+us30WECY8H
eRGxjeGZMzy0VuQSiOaPeVTZjZicLY7IT0GxkFxb1ft/lKYB3koFuGVT9uC7vRWfjS/iA0L24Q2M
34qhSHRl4hWhPZ7WkBgsIqthdOJaTltj+TNAnHeQCKjZ1pRcEMyujcR66KMfwrb7H0WwBXSfohKk
e6axJlbGIhPIDTkRrDZ5vlO66HNIZqs2mJGmW6aQBXw5DpieribCb87uJFKqLa4JiKH74EkNdzpH
dHSooUWfQdpSDdE4wRnXHhfohSzzWTkFafu4cMCISFPMV8Ozss0nI+L16I0cu9cSIRyhoii+BBbx
Ar0v7/qAxK3h0kn3Feloor2uMAH8SW4SnPBdplKHwFK9ieHZHPwNZmjlrq2JWa2iRHhScakqxEUI
yzTSbuiFt+HH3O1d+Cd6mh6fP4HQGTolzTvkk8iJJ1nIvXHu83UeIZsBJsJeZXoj/F3F3RjiGn7V
o7RAYAr90Hir3i+Sm6Aata0jdzSLieURLiqGfoETO84ndCKqSLNIi8oJhANaL0RlOqeU8lr3dl0Q
TdYiKSCbXMfbXgabuemfj5FpsT9l08LSY6N1Q40HYCMTNjLA79kAfuA/V5LW5z3zak0Wz7KvXrC5
D/nT5dE62kStWE1ySG7qwvjN9sNh4DlQkqYSo0yU8Zg8BjC4mmtnmTkk3CmGMF8foGtfwt6qBR3D
BsY5OGw91qV2G6hyjZElnOK0bAKtVUfvjKLhiQB5ndXlT8b7Il8JnFbRNKt5jMUBNLYblHldFY5f
gvOa0PIyiMpyEXlbpETC2b8xmsqsWkpb17UfHrXmk/Z5IkM9DcZ2+RmtuCm07NSv0QG4alXAMphw
Qc2gFQM04DPaZE4gk8fzEM6Fzf/aWkbuyhLAqTNOGV14CmXr1NmMqLNyeSBkAXPE2ee3TZ38AwEV
UQ9LHMOLMyPUe4hGw48fHbe+sahKLdmTwkCLO5gW8cyt35NetntBt78/sQau78/XVZflvqnG4C97
7DUG0o5aCZRen68A79+YhxNdAuF6sbT2hbRmqbsseV6jJrB8nppR09iYeEoNcuTzU3EojepoTJ00
zhd6bvzyarx8ZVPm6aqdJa42ahurKmRgLb2bioOjZA/0jYHOa92bjlDOb3usX86hbojCnHUVM8n/
Sb6WuTTPW90t5Gri1edTasATyKJX69azIIfEVXMqHwKivscFJZ4KwcrNtJeYY0CXx95inU/Z2k8h
xhvMIUHHkHDN7Aq2PZqXkdt1FFuvlG23HhbkCbKW3jQJ2rfRqbKGuu03AKF8lexEYHyqTSc0lteu
n+xLozXMyB9GzMKuSREjvsPHWkwQGexLXHT6vR7VbarLZmlvMnm3RGtHJ/kPLy8cj5uyo1w4PDtT
KC4hN41CnefEK3kdLcDiat7REPkYvtdaXXQM+SfDeGIeZ3by/TBX3t0bwrpIznmnubdZSeGx4Xsb
NVSHUB9/1d6SAKx2IGoDJUhBfouu5Gc4J8PgcKkdWLNzm+pUVuq/uBbw2n6oZZSFA9Z1Ap2qVI5w
QbsoW7p6bUS+uYqhLDcpZNPJsdg2WNpon3Aj2T+Av61H9yGLqoEvWDiLvPIW1OO9SvVtVHLRI5CJ
TGP2I4KU6yQClxOJ6PQSuqx2NgZCkajxBJBI5e6XdqLnQkC9nlpAbHb+HT82vz6+J63HVMzy3BVD
mG5Nv9U0UGTllo51tSYFzbB8Huv61KfcfDaXarLf5TterC3mttoKMiQyG/AlEHTT9++2+D5eXkc2
jX52wvwEdymL2pgdkbAQr0StkSnH5SBQlrhY3Pgw9uJd+JgjpTeePyzGa1vY+Fv0THhYjoqd7WmH
8KFQjLfm00C0AXX5NhZOObN/PNX6qmqYUrgv/HG6E3/fN12f47Ipf2h//nS6WiFNSrgfcGMA/y+q
HwnsQI+hFkVMJ2Hc4+t1U3Ny8Zntz6jIGmIDSlNMWHtAkH2i1x1Ja7Pje8oJXLnQLBomliEcElzg
HmvVntANaIU8h82GvDCvcJLdcMnnFMex4RC0bax4Ao3Wa01USApMnkfpPCNJFvxX6sqqMIH1X75I
V/3g9xwkASPovkssW5EsQj0TbmaEcitzCRUUxcRG5Qr/mzpHHA3nGk5sw4xpJKxz3BuuGz2dGyoq
mIus9Mxfp3aBfKx9DmdI/ETEdPesD57uVe97jM0dqwpaq+dZDT9RAMLvdiKWT5cagz9RE59hV522
RWw7vZG/8Fh2ehmouv8QjF0c9HOfeelJ7rQJd9CJHptEeV7YamSpQDWZXrcoxJlajzvEXC+hVzdW
JuC5iNKa/2tSE95NX/PCRJLtWfD7l7CoUZ6AneJf9Z6bFa0NEBQcfiOUbbWlqNPmN7+FukPaNd9D
fLrFEoNue8nu74lLCRMlsdylM9tGVdZVZ1wrooSvX8KwN7t6subXLReFpEaUaMBqvKpI9rfYbppb
/d3t0bF0W5Tz7ALUZ2Qv4LKdn0TseOjcVmX1n43Baj3e/zsSOUoAcnrYF/hdU8f9cxe8QOvSPAmH
IE6ntYK56SEl18ucN6mfWQFdVwMkEMvv9yaUtpTyj75a1ejrKCV3+FpISyjxh6icUl5FGTuJ+OmO
FlGIGZoRcTHDFbKvYej0FxfIHu4CsbuQ8xp27upXwn29fSDo+WatTD10JdFWIZwbBGPorgJByYvD
X6yo1UXezCXlk4vwNGZIywqB889tl2x6TDEkGfI4WPNbhja106zNXISj33pYUZd+xRWmYshfSi15
tOg/2XmEbWJedFrLVeXXsVRJKWstWDcsrTx4CFqxlnkDUZQMlhP8XeJmTTPeZmSKXtdos9Wx8Vcw
8VK1DZIObUkWnPQRxZbucag9sO61uVu9Gfx/ApmrHMtZYMGE1QmHyadXNuZTPuF+VlbRGw4ify7f
nVGbozBuAV3LcWcNv5pGN/jwX/olpS7hISS6efn4iOkuyZpii7/VwpgsQh5tIVUmsveAIV0uiNZt
dL49TS7SzbYcUGSdYcz7E4xgFbUXJkPi80Ps6+iCnfes1PRigEPKp/WBpAiPJJalihxeN0PMPRrV
FvCo+RqAtvpZjAhMWyHIaEiNt8TgSfgk/ldtVT9WijJn4S1iyZx+hQqLOn3puZDDxBB2NjQV5Gj1
H62eRZkrbM6npZYa4IrKm70BhDrUxYpny9FJgSC7aehWYcSYJLApgTzf5qgrQQiIQi5zyLAnMO69
QjabPxQ55EjL6R/0FRAFERIy190f51alhZ4PPkZTyrV+lndcGUWi40K2z5IhACyRG+hjuCHtb0VH
ac9inFtDvNx6rW17YdNd9Ar1ptBNzxXPYgezb6FA6EO19M9bsaR7VvqkpGwTQSShIbKGZL6ONdpN
TqIjtwbi+fCtzlOyu5hOWZ6QLdJZufUJJglaj/dbGccEEIbKb5Lt82aF7Ymgqmldk4LH7aryYmFz
axsfAePIdCZzKIpxqA5dJjt56IqfTxbJS9kWIeKoU/YHHO7pCeSowHDm3lMd8n+OvSv85c2pGQWK
h+zcR6UyoMrShp0NRn4g1b8qT/VODHd/H3mA5OAJgmhKR9yiA5cL6bkecN7hJhjjvZjcy9cEma47
nlSZg4wEgtLzNL7XxygnRxeygGJjYDZvOJHNe8uFBaaeNDhchwx/2E5VO0yJs5w5NtRBhv4PRMIa
SkV6VClshyPXUnXU8PBuaOGuj383Hl0e0He0IfeN19XBs03Z4mCxQLRPOm2CYOpk3IhFPHpzwPT0
3Nkr9U3mkyUzNqajHPHHG4QmCIndpT6/J/TOQfckF1ganjieF5K/receSuLS2r2hnVfK+8s2C1Ti
evLs4qCtjCzl6ZjrHKr7h6vwYUzD8h1xy0DX6yA/0p3XTno7svv5526vaUPALaQz+cxVeIhxgkfp
6VcImVx7OhBpBG2Hl1Q0PYmRWqRDIun0HaOfVHB56YO2Kj9Nn/wej5UXgEvVBYabJ6mEQaL3gtf2
KkltOG4K8XbR3r5m6hVAUArEZjVQGnMnssuylqxRMddT6W0KiZvF/GXBTvZ6OG2M/DscuY00jEsw
MCVKrOXrn0DcwBl0pnpTkgA4tOjI7Sf/rSg81/X4XDQAtR994sUF+mZz6/Gpr2/JrywzREJGWnt5
8Kr1WNwaqYgDsEioA8MlsYkGmNxL32orL0fEdjgnIm11otPJJHg+/iAUROcRbSLh7IAycgllNPmq
d6AgIOiHDr5wQUc/lJNIyLd+F6lpxR/N1lDLbk323uY3nYEYrj9t2G+yaU12tEFjsQv7yNHyPaQu
Y8a6WtBrL4C5RwRq1rX3YxOQZvN8447U/0qxQQdXTcOSgTw73xwO2r+0Rn5RDQkFAvX0jJjouem9
Liu04h6LTJnihzLhJ66T/AIux8xoykBrC6yvsfpBXq09BGhYuZCJhdNBT0V6qLhhHUiMvp6QAf8l
KaAmeLf7s/3t94+GdQbhIB45aVSeQsfNXQSabj7WXenSYtAA8WOEKWF7lZTWJWDryM793oAvUPIl
IuwWka/2CjrEQbnWHwp3cU35tp8lqB3wS6lTyCONYuDyibmJfcDJpVPcxXyjwDdg3ZnVDJoU/H/2
0n7JDkB2+fWwXWC33k8lUyd+VbOQkkJwmMF00OMPrJTHTggm29c8aDIq8DXLyJkmCAVLmHuU0l+u
b2MtqMLvJ1CyN7aF7DgPBtG8MTLikyIG9HPNliHOILrpAI+cyD/mUKT8+kQpfBa3T1Tx/sp7Jl9y
xC7h1nrKXTfd19vuGm6pBgVKByXOyCpEyD3fZghqswnFl+gy5c9DdPzfIf8O7KAlf25Rlyo5Aob7
GaesY6qq69TGS7iDbmA8btJJpa6UWDmCE+QmODx25hyy8EgNMS6uVBEw7HIywwVJU+YpOhl3MA2g
RzrmF8PaGl2k5qN/pvZeHchjJnVjSpqrW0Wp4qDqAIlYvqKr3PdlX8fgVT7uF3IKjfcC1wJO/sUf
JbCTu6a0THvbBoxhm0Sc+a2ubzTdylPa4hThBSKS5G7a+k18Av+Cezyx2DblwZ7VdgbMFmkDMic6
boJd+aqZLLNf9ypHoouPMU96/E/y/c/FEdGSapBPgOFT+1s2DE0aoFC9FUSBvU/Vqn84biNnN1j5
kRTosi9MU+ve6IZEX5CNxcmImbELApJjwfcBUEfSD8Ex9AoRq32C9ksu9fPU5E6NsqNpwAwgFwTm
R6wX8dRrvkt7yJ0mZMenBa1IUAagEphfrgMKfqINRg54WnPZGHYU9lX9p1YNc4rKnAbHIWpnQfYT
a4NARcSl7AxrL9EnN89J354pw3f56h/5vk+4bIjLc8UlDI24fbgUnfuXqoIfuF1hjMilaKkgPYuO
DNEA7+Hdh+DCIjNO22oLBsiOmLblWkcnmUFewrlqY/gg/2Q/IEpJ4uT/mY7F7uLdgjaY+32NDViu
C+BfIYxpUNbbZc3Dtwv4TVMIhOpL+MMHb1VgWph76eS4Rn9yNUP0cT7SzuqzAkVToJ4b9ebKlTD2
6dBs+3vnO1h9nhVzqw2F9X7jcrQ5uMJ9uVJUjcT294DGdKXKnjPqCdQfSFV1+ylbKhWEsAf9xfmX
eQ3hXDeWoWhAN38k7yYbBJ09KuWLVlvhd+0ASAEeVT4iVRlMGzaHRYKi20Szj8NrjnXVq2/YdAKT
TqT0SrijYase4kYYroOGmD3CmRRc1L4FTVe2mmWGgpihT2A3Rs9J9Bahd/laLW47uDCb6ljkv2Lv
i1P/oNWvK7NoHtdqCvvI3n1Acy9wJEFyomPpLILZ9DdxmuN5PbOHTbeFbyPfWY0JNpgbpc90/1W1
OOLq5NCIJ+cA649NNM/mh34iDwYG6Wj9xx9qzC+XSiDwJRkFUJn9EjhO89X2P/pGNZRxPzW9Q9s5
+xRKEx2nrZ4/I4uDV6CRdj/Nfs4a8TyMa0EvlicoCK6nS0ZfKPcYyEfq5fKpf7156A1eTelu8Vw+
Mxs2WFYZFZLkEj871M26hC2iO1Y9r4f3Py0HCkmMOv9+sppIT7ZSauT+D6xastd9PEExxh60CXEn
f52AD5YJkIwsEYZ1cwKNHbRspFCgqId9I/evCQPxhzLMIL+TJ7iccEClhx3y2wAZTgLo62kxGD//
VIpNC5av7mZyQ37n9sZx+VyM9IrRy6tRyM3tC2s4jhIXa0QNJEGJwniIaqj6sTGywWeg+A7zVjGx
7glfLkx5IlQsLP3MI3CldNKxvEb5XDtv8sVM2ywBYqTOxlq/5PmUPkC/pcalNHvYZ7aWgsB8eAJx
C7RSv+7l9eYnYQecpGe7pfzNKFi8ZI0om6P9SGQ3SfQ+0u5YSQYchr0nrhNkjPWWRIRSXgW+7mc+
RbUxdqoaSmHrCIdNYtlajLlSLQ7CKaU/5nXk0SDNEumEih9vCv/P+zpxFUyxUHpjhoe2s6Xk5IGU
646hpHHIr/bkAOkV1jh6gsuDLlElRW/l17KIdY5esBulqwXxl3Q2YcOArO96HqMxQM4t7hsHiyEA
+b3bM6/V5fNL+uGoSRLd/j9tjmKK0FNGj+pQnPRCRZSYTLLrzCzA4ASMGo62GwzIIMO7ExFetKHp
PvmfEVDkY4An8zYHnx/0Klw/UyN25SaO6+N+Ddw7ohhde9Tl7ZHxG0gs1xHOtlCcgwGEEkMQwMFb
9Hpn25c+/Elz34qO9lBFV/MGzxao2BKjpzjynCLPJBATf3Ih61rPtUDrIX+5TH/5CXYuI1o0bKMW
dxPJzG48zKYFaMtLJcmY12ekNf2+djEpMzt/JmYAfQYnhGRcDQIIQvvfrfp6zZenbgxcU030WRku
PrgT64CUhCMf/PkGTE9goTorIPZMSISe4e7g9pu2fRdf1tgEfPaUmIhjJ/xvY3SCIskbCP/AC7bT
uyPVBm1Cg5LK0hSYLJZzcTjhyP7pM6J4tO09Wf5EgGu017XrSnvGRaLIdPx/IjxKuv0whO2ILOov
8RiwPmhbOnf5m+lbLs6aMRZmi7oi5b6NPP9DHD9jYNJFz2X91xMcsaN+3ef+vWMD5YOKOU5iPxwP
vwCbvwD9tEfVxMOQyxQa61yucGh/3OJgTu1SF/Am9YVaysJtQDjTmETODUIWESGnfXrZGJGGu5IM
Uzt9CYF5b7uKCCuFEUCa8OzMfqewreaF+ACqVN1WPX+JZc+usqhnfzHFw2CJwcgW/MSHI+0LGJQe
ITpm8SAnEpzX7kc9Btqh92xDXgXQHpqHUKa4frHGu2whs9wvaob4bcu5nugvVIxMRw6bU1Q9GAJp
Y/3RI7lREl8lSABH/t/I+m1rOvieebs+jPgiV0hZ29S12jnMHhR117PGoEcW6QXzh9nOFeG94T6U
/+jK1Rk7FQLfdScG3Sz2HKnlAYrC41HvM88GRcX0gthjALGgQKQSIFbdK9pSflef/CsOvYNBZZ1O
yQGJBjp8aDLJmL21AeS5PZ3IcGzNIooEvcKfg+evSTz4UE7m3/TTY+H5gdfXQSmdb5k5QSH6Qqev
YLEDxbxrd/I4dojN96XY7+sS2AoeVa34VPVkjvlCShmVItQ3BitelCcM/TpDpSzE1tikZe2FW1fL
2mVBEk1XUS+qANTiBJZ5MNWN5Y/f3fo2QegmaLEwshZZg5JawFHG3kb0GZWJVzeW6QE0nuIW5aB4
FOXs9KVVBDKjb/PdnZauZZ+HyFcoe4slWImbzapX8hSzaup3hEnQmipc4LDdhaP4b168IjZSI7B+
e2eYrHYa1Mylo6dvMvVYrxNJqTnONfmCVFcEULWOYxtGtEwmdFyrjA2YKAqaBnXwIEXtmrM+6FIO
ZPnrZG3ff1nb2IL2T75V7xu7+LCzwynPqhKE7APgcJbJLrXxp1WrQHGnjDerex7dcmetBLuPJyYV
B+BiLcOqqg3FGVG5+O3nP0TUkub5QuoqI0lWI8ds3geHkztAVPh24OItd7mwCEZfzN23wKgk0U8H
Ubu1aYcrdChm2jgNQwVkKKavFqPopHfmdWA/2TiDx/3bgkKy36ypLPGohtalqCbFggWGKOzlJFTn
04DXY01diIMC9Z48sEkR1Hhm2NjKNYzFmqbuo1SiyU0zYZqLgfC7oYhNO+wzAQRDnkZDcYd3uL8h
rpvCvYuL7nmWYz1NekmjBe/u6Zb/mzRYsLEW0zZ1xPZtuEoGU6bfyJAbaDcFGc8cx5zJ/s8346Bk
QMOCMtNDvdseHZ8dFHhIJ/QF10ZZlWdbp5Zno2Qpc2skw07p+9aFCS6yTgBXg9/RMkgmutATX25Z
z+ucqMYL0LW3Fs4+IPIOI8O2QzIQq2SrPqCqqnkyN7NxDHZ8lK05J2aP9xCbpuVgsC9YL/U2iqla
nHFUied7093wv3yeYAKMTXjAcg4RGk2WFGXPzrTQiqiDeMxdTmyPr6vNv7eTsaAyuGIS4Pe2rkZq
LEuqouxVeDoyHshFfRMubsw4BSRt+nwqP/vffGZhr+5h2RU4bg/aDQi6IikCtruqixPOoUlAICH+
xTUCvcLzsPhtno6zhdkzhLiA7uoYF5jgHAuJqscUEKYH98VJ5eujiVZLBM69LR9ZkqXtZ+x9AwLq
4d2xoBPyMKyRuSZoGrmV74Bv2LTAjAYfzzO6Q4u4DKAazaRxwgrjTKe2gESEPfH5YJgg497++BYu
gwlshqEMQG7p26sG/OVp19CF/babSeK4lRESQqvMJ1PuVYFC2v8gtMcgpniBrP+nPmIKzkH2EeM3
oM3Ny7hNGn5KeuRPEkHI6CRa+QfDYmqEq2c610cVBDadehu1qJG5ldIRHftZkyWAZA8ntjKyhwuY
3o+FI3lKaXRhkOcmNZ2ovpKqayBDoUe7dAAlUxGOPlI2x0fXvkWEPkt/oDz3CPSwIYGRzClSO+sD
P4QsY4Wce+une1eY7pPdhfowHI57lbWWDq07EBIedDAja1qctCV1OENwN1yQPEm0nUUhFjeivRP9
uiwRSYPFxkPYWcCdwrDaKRN447icMiIvIzofM4VJ8FWbzuALImwabrFukTkC3KoTkMVRJKWpX7ey
yTJ8JLp8qTDZX1kUZ0Gao9CawbVyBV19w4NrExJoL7lGRJNm+MdmJnqx/3CO03GX8O2oawQwCNUL
KR7S8eeXFsbbiBhFQVVwdoXC4CR3GSP1uirkjnJhJcfrKjiXEm0CG6R4C4hVKa7w8QTdF4vp0pSu
lLp+iB4chMtO14Sjm2OAEDsBpsCs0cuo3i4ysP5fEOhVZGNYPggP2PsFvYPqZWdKjIxTsivPRbXH
gxFEBBfbrYFcVoLeXCswAZ2pXR7Z87d8mDxlCMm5mNRy2VHcjBExPswxBOLiDsD4gacWnkD/tIB1
Fy9+607G50bZ9Dbvi5bwfZwHWZJjCc9Yo1VZqql+jHU59j/Knr3H1x4F/pAgogqBPl0sklGaTo0g
VKw3AjdsP1t3gYWeReUQObYdpWQxCMPGCkxmHzNVeIAnt1z+o8fGstGyriA0BtYftgGmvasMjXKl
Dw0/yise4VyTLPvEot3poREXlNq9eC/NMtwVY4u/SgG2y5le4wkHETlZGx9C0zFXFKCeXrAKi1Nx
c/jvO6uNZQ1q12+K2q3L2uauULvYtjkHp+RmZgdjYHiTQERNLNXAY09plBI8Iif72GqBUtjflEWd
Jl+SGbM0ZMUfIYFzMrgAdb1e7xKwhz0JDeh953ujTIgcUh0miccUqFUw/kZDZLMZy+kTh5xBUNUb
IWvZkwg2OLe494dmm10zbnbh99L0UWfEbF4Gesd7EKBFZCj2xCK+o+TAQlqsLbrUgCL1qC+lb7fZ
lXcpkOntOcPMoUqFpyZnzAUtK89yTdlsy+xjjjJfnFi20GV3FRPqYxmyb7SRM0MKD4Ai/97BRXr6
JGNSvJHZX7r3UviDTvjvUrLI2MltnE/yvHxTkrLMCDtzMP2Fgv8xzraPQg5+P1j8WLx4xJi67cM1
Pi/6JspkpwBMfSxP8OJZaBF6blvbWecCmpSYL0o/uvQ2Udt3hxZ8SPvdqGdwdZR8HRIKtIkH0kXy
T8rozrvVuVRu/zmJSU9l8P2BygXtL1Ag8qVTAGL69tPYHTCaIYnpfqCfhN8Wo/MGTYVnHUbFU6S6
mYNIYuJ53cVY8Ob+rk0pPlfSr50akuwGCikyv/btdv9fBHKVnlAAcBEX8KHQ1VTGBNe4xhGrwcfc
Rc1AsmiGfUHmkJ6Q2Qp0CsKrr5BGlSiKosFwPifvIBsefwX9Pc2bWNcL8WvQKKYL1iDx9uwwNYQG
mKWmeWDMTRLgaE72JDgOBj7PIrLebI2isMcac34rFg6isd5auRPi4wGOADFiCKvonCHYVtVNnP7r
oxfAiPXjlRU/YijIkmQBGXFzUSZQPpCKKadJzMN0BqC+3OmYmFbeV8VTBikFvZgeykQkqQAu9pBv
St4kjxh1CY1wMcrWBGT+sIRisiG+SvhyatDWIm4DGD0xgExwR6xW6NqynY5k+joeLQxkuf1wQXDN
R0OEpM/gkPinhXqR1nSmErcBRjtjSaI7shKcDYCtLTLdPnKTDOMWFbY9jVCsPM88ZSnx7lIvtJad
TGl0mUxQy130Q3Gm2coPRS0PCswS4ag51btRfj04jTXtqLx7VudM5qemm6aeAy7KPxlbJiuaKIV5
d7YTZvp/KewuFWwicXAhXVUDWcIGld9oXF0u2loVm/TMRXhuhZCzvv7SoG701ySX2SvIz8yk7Kii
XICbeOmVbr0KJsuSvGWTiHeM2HM6oCY/DXM8ApH+WZhF4L1CzdjHff0XMM04OQb8FvCH0zaFaF8q
mhKVDV9iKAkHGKDSEhQQ6G6PyRNMzOGGDoUhK47G5t1zlMsFNWImQlIdMG1lrr5Njj1++gESPynH
O8Ynjbr040igiOTioo+6fY3G387Paa0+u7bNPoLK9WnILUVj/2C9d0kyH8SLlGFIGbNgO6BlRPXC
lyhatwTg5RoUsm7/E+D0GhYVhU57hd1RGCpmqbGb/yKxEjaVm829e3MOc2509+mqR4+GzZqOYrJJ
/TESdFORGVRlCW8lYEd1pCYiy0gv+WfXG46o3/XqrowY54ro9+PtjbDhcYIF2f97T5Cx5W3L4iwR
gfHCwmT/b6UGe8AUbG5euBtxB9wCKYv6Th5jtVcWNfWZUf/2CWWy2Go6N2/ScCJcy4ya3rOe43xb
D4r8VJM3ftp+vzln55mkDT5QLwbTHMiJ1HnK1A5B8wneA2WxngFKFPRAxPpJNNE1d/EmXl++H1zE
Goyca0Fxgz2KefwBzGXchjph/6hKkYfp4IQ8DBmCXsypN+e2Ms66RucPIlS9gbXnORSxqslkvfF0
n2ywxR5NUphfb1p1u/K4jkCOE4a/en7Sz4TVn/Q2DpvotcGRzyXnbTaoL5zkUTUtbl3z9Ncv0k7o
3eoq5ZFDfi20Qk0q9nk/Eyog1WXTdnrlYeQ+ZMg/hKlbtyMBZbNJ4NUNijxGpkL1R6GXoHHCRYNa
WezASfrJvmY5n2/B4DvQHccC118mZZ22jtHihCq8nsFhU+s6ebzZjpHlY4zjx+fLf6YoFFDBmba7
8r7vRFhTjCFuqTZ+OZ7M28m6kG1pJOeH4lcHDwrhdclKIndO92F9eOw6SWUOKyZHexBQrrzJeL6g
SONh+U0d9u2m9OjmWYIX1GJdZ+aedXN/1VEF3mYg3CBrHvBoC6ZG4zawxn/FiDrLC82uwetsyV4O
49UGXQldBN2pQf+/S+aE/xgyqiW3vIUAdx+xjJREzIXMbn47u61LPC0ArqmOZlFTpve58wGZTkZB
Jh3cNFuK7Wkl/C0NwEr4q+V+nM+ZoiXbLLnpI9DlzcLMGcNymVQ3TILn578fIgN9foJeTIRlanTe
5Qgycstc7rY/0CIdndFUITUNEr0uGvpkn6SVN6teJjtJkNoaNfZM6nVk1mtQPR+jOSPVShM2qbz5
mJdivd006aCLL3ujJkcaP1cYTPUlqnNXDPJxHyBJJBYqTpo9owbWSChJurKreVoZR4qselDYy2nA
sRc01fOVCzltM3GU4MzsYdbKweCZZ/4i/SoNcxS7Iu9rOBV/kz2+rSWnLUytTnrgKlTxq0/Bp1ZN
KUAh9RVRyvaP54UGPJUDoHWaKSPpZPGVEfq3bNuu/VCZo03Pzh4/FkXpvmTR7XPEU9tZT5u0EPrE
sL81U/CMLatL52ZJsyEGgCdT1hiyfuh5oB5EnujEf0TtMjEfKkduY0FRinL1/78XLGyHKjt2d9VR
nlsVSbn/lIePPEaR9woguH4elyPRWkHnxuJfiisv1uehRxF1wW3L2THDMZdjMN0s8bz2s4UkW3HF
tQGq9Jt/n0tWHBMEojkduumTiKq+w8f+dcZxJdrbSImWy4m8A0tccC0DnqJkgGD4UGLC2HpyrC7y
6CjTQZ6/mYE3+2N+6k8c5NLsJn8fGAblvKH1GHSxvt2/O2YlrT7Bk4U5piUYVINzBliEHIGRVNRZ
fh1T/rxfDsvgLWa+jDFLwGIOXPfShkRfaWozft7XixQ17pbqClON/10YbONNt02V2JxUQhWkTul6
tkyoulGIXdivM7t0wWjyJAw5STz3n0JVj6BPR1audtQU+D7xIfO8I1/7WhJOiUjbYDt0hVe8ZHxN
1Dr0hnn+WiQmRSkiUntXU/mMlmjq1OUaE2cUaMvZ6qlfsxZ3BUOW/vn7zljA3cTFQyroNdhBRCsx
73JEqO0kQENpZjn4ghjpOORvJa30CoFIlg0eieTomDDnWZGryuACbZKmB/jpFQXFeDg3vHOcn8YX
5+w02lv4F8aFkieHwRAPKt08A3NBCHDxtXdTmYTJeuDIG1BP8IKGT5tWAF4GfaAvNwWDwArdIb83
2NvajFBbJXq90mccS6ViOrqBH54t4u/DY0DfCWWpZwHokcvlfxqc5jloUx79m3B5+jDTaE4JjqxF
4HLe+qoW5NQPmILBBg1G6aDpvy00iy3mkzeiS3DJX/iyNQG9bg+fsFfJRfoGyXcqp2hMcF+5817c
nPol7nEbJ3z8eDyf6RKAwBCW0+9C4F5MDhDc3uxMXbsCvu06g8tNnSnQ4VTzZpBKoVwvbklEiean
Hgas08Xi+StQBlGVBFA3zCLuTGHn0ADjHWQGRCfnjEuMOSiaIhjHBXe1V4rCVRa2pjsEbdicfyMQ
GuAqbkly5OY38alJ2x07avTyD23vFMPGVmwGP232nFV+RFVvxqdbNUWeyCmH6uxg0O54TJUlAKLt
7B2lwr2YnEJgkW6LkeqBaZaPNbYwCRpLDtVNFEFUcSIVxFrRz0p7CVbbFvkee2KQz4FpRbo+Rh9L
7YZChb3gn01XvjC5SGRRxr6WhuBbFSO18nITjpUTil9Dg5K4V6It0gU7HLUoviBEuSOnhbGn/L0C
Xf79c01nPFGNY56dE2ROy9/cgSej/kvFDLoD0vNk8PVkp0mYdbrJv9l6odOp4LJl8XSnYBA6aW38
wFCdeBzkQf9m9EIOwumQ1cPfRmlEWgdCG4ubRdTHaPeqk2IN1IiIMnSwHNcFcJfNfT9GPKaTkxr8
o1dDU+XzE6Z71gikoV2DOwnJZcuGYVzRlPqB/DXHce/cPiK2DMfDEx96fTZozEFGJZ6wYRbfMlnb
zXvgqCQ5d+2HaIYXnlFSF6NMmEE3PbwSKRkvBSWvzEv2KTlNHnL8HMQ4B+Ui1LFJOzV3vbbaDA1B
PB5SPsIEZtymI7agcVxcBGQImPsP9QGCkJvMnWN5kyOZPdudKQPaRW51BHC4Nf51tWY41LbqrG1F
0gRN6O2yZ5MLYZOaRWTX6tlpD68v/7nkbTIyZL9n7aQdobIPGr/Bv8OekpUtDd4OFxviuMUHLuHl
8OeAAtalsdVuWPeB2mHuNnRliMrMkghSbtz6xnXdF5y2dIOQmm0WFLW3id0l4t4ECOHxMZKYXU5Q
hRkyVVTvAqWKjEZCB6zoMUTQm8ETVXVXrtoUXiEyppz9i3dcekE8ctR0+W+Rw4+k4Ib8o3FT5o3E
biUevS0FJ/MbcpzL6m0ZZcL7ro5YgK+/wsu4crHIUtJgVxhH87/77dTgHR8z4cQy51c/NVHsMia7
vpGJ8SnHMr4L47oCbjnFcitdgGaLcAnoOVfiL6v/ApkIBnFQrim/B+P13CfD0f7lVXNWzrlujgvF
aMb3JSXdvsduU2hnHOZdLZBBPB7zV8orYsYSxuUuTo3rNdcobpABVck1T/0zhoQ85rMitDy2DOYg
2A4fm6CRN46EfAGFmwhPPI4VwcSBSo08CYHtSrTkPf6dLoxijjzAQM5jjvtgmD2jkLUqehDZAczI
G7K42QhOsyLZeNKNIInynAxQmyYg4okSp9b7kko45WtTUtxSKlIplXm15/r/JsDj2UbA8Gjprf92
NeG0ZQAH+JfDC383JKB0ih2YGC6bhdq3YhvlkYXVdY9++Bf4MMZEjQCtYv5DT+PDJk5OZLI7kX4m
6q23nUTYWkR1BXAYAu9wBQstJf1O2T09GO3Xn7nNd543icBrf3TNfef5ERwSQopCD9fomdn2lmKb
CPAQSzZRdQdhCONFZMzRf2fHkGMHndoo5qhsGHcRyECXu50iZ+GGYtO6E80GD7/e45ixU0A2RpWA
x27wFJX6AVl1h2jJQ+QDklWsfDJsKoePfDHI8v0oSbsiMGKBW3LUL7zKRJKfbVrkrNEv4w692NZG
k/EbJdspH9TvCNX9V4KtvuAgZ0KrXOVyq52hLZ1/k9IPEoX6nmAIhM43oFsYHqJLy2hcJqsjWuML
vgU5KA0heXqLIrqza085aZZFzmV2Z2u83tjWfccMEdloepGvc+b5I/2rlwd+pNJhNbO1VGUyVB0l
9hrLZPSzuaug/5D+tJYnuBc1iTpoCnrfy2yuyvh3x+sKWYmct60XYE3X1cDpeBhqkiEb2HRf4Z/k
w1FvhyhA0go/gVttOAVPV+a1NA2krZQiLVAdx+y4ch6G6UBKWEDmEgTi+YU5DXatVOY1D/aTN6Zx
66AjSBVa2WiRTyPFyaeevZl805bbpjC6wlk6Hm+rlsa0tPE6WI/zkKD7Y4AAylL0//rfNRumanER
vOGImPhnxc428kJ0lCCYoLSPX4tSCd2GID3ANHSIsT7Xq2bShcLfraWx+LfVe+VaXDhayF+Cs2wV
6EMjdZ90p8ocz0mfsR8SQvl+v1Oh8Zheyq5BaFf5l/qPINYHfx5dCRb6RAIoRfaqg2k86uzeta8q
ZYxT2qWGpqpRx+J6bibDcBmY0AYzKxHmAZ1vrylvTlJdRq1gxBnIs+phFoMzRT5ZSxT/ZzISzuAs
frBA7KjR2uSBowf/rjqOQD8FgQbTmcA39V9c2HVG9ZEiT1B0iEG76Cwg+JAF5j8173B6bTM0Q5Hv
RvhYSA3k1W+gSSUu8H9tEKKmCD529XNNYYv+qyJeHqPSO4iZwaW2fsYu8vrw1qbQ28dwuTj46Drf
ljc2erNiUsT3RXAi1kgrZrsgiU3upta2OVP3z/njd+qPdf0OkGGJ11ZMIWeuDhLulKx4uNcWGROb
nViGzcqc3PGLNVEEga3oG6ltn6cpTdOPtsF+jqgBFjPpPQAImVKQL96CYDTQ0lo2DJ0ma+hAxGXy
FXAMrE85gaI+vHdztFc6YAQ4gVu2TG3tMKfdZJcAYdzT+wy5u+nb4CKwz7g71q6ynYmxDm9mX6FZ
GaH9e5DXIMmpFkwZiGjc8+8Z9E92jJz3flz6bb/ki/iPpkQ5imVfOiStnHw07tBj/HdHT01F1ZQ3
rNBiZTUW2H3AtsfT+8hf3p5MPQr8cOR0PLt34+OKayokNwuHzXviH1533AL2R+LBJUbvE1dnPIs7
SQFSnR+L4XU/V9yq4eAOvXxuIXMPsN5LZLoG9eKAE1ZhV9GKhRetQXxgb5ESrV2RqTD/292Mc+Of
VW2wtBFAcGTn5CTagURMxTD4aOk91tMRP1XHn5E8VDlFNHZ/+V2TsCyBxbShawGdGYssDyEe/Y05
DHWBy04Oo/jWVoNK1vxtivWVBBrrdADquqvIRQEkoq//UTDiVqv6674ArfGpo8iunlhn7429CWjC
tz7A7dsGk8qWd3qEvpsBidogkA5miVDTlxLasvei50sK8L/XjLZEhx7OKgM0Zze4VVJcZSikng/2
A+ZxeVeB9EzcPLgBXXdrotplmRtvBXiNNbhekkKr7RlTX0hmYz//ML5GbGydIFvkW0LdL20yEVI1
Lzd6nAK2JP6ZBlPA8nNPAbG70fN0/bUQFDtjWjPQq4puYld3yGrmI08c7P6CKUkXriJ92XJq/NBd
P6zqXSn8t4L2rE8qo7ErszktqMvNZIUw1cXOuKsS1KojzrIbZkZo+yJZsnwwuf63v6iHHCXv2+4c
bPr+voXAlQZ65rk6i6yZkyjD3xUJvevK44YibfeXwmWnYN+B6us7QrC6au/IBs86lTUmkEPRfxS8
lCuOC5zfwSwxh9u43vC8+uVboZA6u7RAqFIo3Er/4lGr1nRgUyCjtF/yE+lTZjRleBDzLoi5RAdm
rLaHzIFu+XtHmB6HjgmgvmBCB2hcjYMTkUS1EV9auky9gQoVqcqzDzirvKu/rRsj4c3O20FwRGnn
Wp90Tmk5QmsOfAmSXL01nDUIWW4mg4Ere2Ij0JbuJ2om3Y85vS8qriKzfldWYD0LZshFSRcelxsX
1P6Chfek3IrIDYXzY5Pr6J9ovijLNn55hDsjpOROmge8LNhbgduTWCE8wR/xsdGZLSYRu/LgC/Qw
89jZicTGzdDo7f/EXM7FLmP14dVjLYkAIGv98jfBwnSS5WwOxSS9vv6f2LO4f3MFWZthUSHZkIn8
Qhh4IWQWUCHtj5qVezUs+Iy/mOmM07j3JB+yeUGOcjP31wKm3Osh5knAlqH9QZ4Ok19874RnhZBh
urU6WnO2Hb/UwbjU9aOMw5LhX/OeMS3L6h8Ap1u1wiX0JLogeU2D0qHEoLAFQ10aBMVIPrvNT9hD
dtK2oLMywlMv6HK/LZfwaL9ldoO29x1DKKYn4qlJKxav6olmUfVZh+44UBkDkgaEVFtWSrx3QNWF
gIaAlM9d64nOYZlNLJP7Df3baMZzIPUI8vtzgL2IY+dk3bG8jf0s0u6jzdwj4jrNb6d7pJcwrPru
e6CbP14f9uEDTCDM5KznpO5QXgZer8w5Zuv8XbAXpOi452UFOh6RbXSIx12B4T7aw0+Boomb1woW
a1p8kfQVz8eu3U1NlkSatpg0nELgGpEWC7/1yq5UFPilKgvsNpLVaPreHhJITc8psCvnZPlssWAP
pQ0pb4aR56Km9sxfQAcbiKTKbcLo5r1g5fERTC1P383iIqCkBF1MaSkZO/W2OGJ1WbGPLhHWTR5a
NM+RoHEn0LAeqfhoJwXH14chng4QJwggrPJfEJOza2S3mAU0NbFsLAndm8o1nhsfYZXG/Ahk9saW
zLOvhBvbPS1F9Lpbghn/INKkHNHJouNe8Qlf+sMHZOk+Z8zKheFr7LVbAXtnTBUflfHDF9y17Ojh
YYshJrffDS5Cujpv1Cp03AoL0nAIOxUHYSfFCYlqkNITJAN1l7hPuOWrkueRe/06PINIMVqn2zOE
A0WPZ4JJvi4VuSJ724JJs6n5ZLJilvxUxX3LlaV1/FaYbf7H2Kd4tUy0p6I4weRo6KEE9DJEJcls
GpwqsjwHP3JfrqRbzTHiTD6Bbt7EHtPP+vDBgdrNNUXOoA5bL7GXiPplTXEQXVOMCe6zrKZTA0P4
FhEvjAFBwA1NLp8liP/2yi+7zseFMRHXAsMB17gWDTbDDTIjJ+Z6348zMgyQA1QsBcsxuCgPdpo+
fNBxI1pWNG/FyjJSjE+tDjZyxgA8/ETfecTrVq2SvBKdBySCpFGJqffG/+/Kiz7w2jn4chL0Td53
PHfkRVY5GpktaMngSGu/7PnchOeau2QqxiIuv6u9NkJphdmB1fQAqAK3bjIrV5go78hKUSJpp9mP
XjTMC03wnUSNCwlGGM5oEX7eMa5rn+ZL9mAVQ2xLZ2nIgjW/jzDcav1Amt8YgkJD1TDn1E49jKeF
h7CDTP1Nuc4eyp3m3X9BhNz9iZKL39Ho1NcmPiobG98GEGAYluY7kNxECkOkvHNoCPT1RZ6cUvHl
RMZhScqKmUWQQz8fUQVRkEE9m5SfDvJgkrL1q9fq/Sv4z3Mb1fnUGJe6OjJ6921j3JA83Uff831d
PMpwRYK5pw/MEEZJ3ds8Ru1xTuRbJH+Q7LY9Z9vkcSIxODxO7Np2MQEgpKiLgTETSjcGK0L2R80z
ff8a7OxJifwWquZHylhjoqUPKjM0emgI3gajmpTwrTDanx+fUJpLNmpUEryCnISOiaou4hVaNvAM
FVdv4Kmcmfy6egyHKWqcme45rTKyId8OlgSVovtf5F/S4CnwX9A75jdp6nlH/n2GWkFN7K2cvAte
+B3AlBWkvjdx0cwvmvQDMT7/RcV3alX/oOb83nXmSHJ+OQrRr+12CQXMuYuKhMIITMIozb+fEvcP
SBnAJMQN5a7D6m8SgkJ2tQj4su1xRmiCzuxzPZfTDt2ly3q3fzpPEtYfMJY4Jyf+DgO9EaiPOL9/
CIqCOVVSiGzboh+LKWM0y1NQFYObJDNAyDw1sSGzszaClpNfLO4pvkbuowWXURh4Kx/I2lX4xb3X
mD0mqYr67DmRTFFNGER0+TaEvjr1swzKVd5RoRJTBQTZgGlDhXW2PFZvOIyBIIb9oAG2xAZ+yOnb
MixSZ+ZYBnDLwFrHvPRe3OgG7Z5kRXeZpa7YdUG5QQJHB0HabkXQIyJHoSMrviwqHqkQLIHmVT26
+1Lf1S7mE+GVC22XgN5rymBlW6P+e9eFOol6DYAGndM8zGnifH/cMHba0sEm9YAjdlExPq8JFu5Y
UWlaj8tcsngPOjMJcqTtm5qket9XXeYIpdksVJePHVS4aKUV9edn7ptdBDaTmjWm6Zpl/Omz6V/s
jmx3r/bVx8w4rG1sH07fO9SgpZbTU6OSiOquvqPiAEF2aioDaKKlGcE8fNf78vKItq8S1WrJsIVw
k8Xw/1SJEZWwlwYExwDCBSyzwyH4QZ7jRgy2kTACFLOAy+1BOsEji+TyPULSrNvODnaUZnuhnGfS
aHR7vOtgUKGHSjpJXmXpY3XcAmKQ05pFRIx27uiRwyMcVCgTlFmplL3fNugBvD2Es5X6uSne0/hu
eiAUkiu1Dq6bvel0KghFQxxr/+jiTsYx3DMDA7AN0EExpQOIjiFNxDnokKij5A0i4Y/SHE1HD8gH
CTNU1JzAAVg52V3RsVHGyNs3HcYflnWhV48Z4iPluZwoEgmhpyYS8DPFX6tRNaO2zPFoNkk14Ltg
SmLTcdFDVbtpUc63XSE406zo0Scqhi7/fa404DnZvB5tjoQB2L47oFPP24Mt2tjBSSE/8TkmhpbC
BF0riZL8xGwpFNTzSBeY6BTRnA3H0FbkCS76gqvlHcM5bn0eNllrwUUF1pWl1AlrbLTlZF1POxcs
P86ByHLLkzYx8XWMbgo+F5vSkFqmOzvFDtLfQz20aa82+MsSz6qN0MhTSxteQoUDEfchBTt58MM/
5iWzZKSureeNbWH1abryCwRcEI1lQcWGWj1LeksvpN9kjlL0+JePknLRLl84xMvaToZ6pJbgsbVd
JIgkmco6Jhv3nL89+ippCe7YWFZTYd0afHb/WABYto6flgAle9HXpRkFpVJQtCfSrDXopCvAjaP/
yHPm3u90CQ+rM/lGfG3y3313Wgs7DdYQmpTYrzP31n6fdlE5gdHYu6Q4OkXt5YWfBCVkvJM/yga4
caCmo7joy44RacHToxezRGWOEutnenXJ3h8R2V9ATvIVPmm2Wktlq8zIjFxPnjaiN4IZjgA+U0W2
rhpJagsABpjkzd1vj7u/vQJrr0wTH87yItcXM0OvyOfKniZYiP90ws5mR5nYVx3q3kMztelo8mEZ
7JvbeFtad97PQTjolwbs+9YwfepVTz0v7fALeTc1NN77g+ThUcCPBnCD3RC6xfbPhbg49EuQAv5q
0pnriJLW0GcRRWS55+iSw/HYsrz0JYXSHGLK8kOFCHL2+xx9zlqJvZB5vqWpJeu01KnPNwHGhCpQ
u9uch60Yp6TjOKlLrxm4xwD4e6Tsrmd0EmUDGK+44uxyTIq1Ig0oh/Fo4PWaGNy+gIxIyXSocT8U
u0Z6KIWs2orl8s/y8ijIXtSSrKRD9J62qED6isjsQN5bvnZ22Q7TW2Xl0xW8SUtBhGiYUyPpLZSY
sEaPdER/vm/4hO5r+FazsMrd7DiSATipb0VVsveGSZQv+NroxRefoZtCPCHTHp6XVVJoAT/3qFBT
QqJ/y8eLDuMbKkbH1HTG8E3IM3MCYVrBrdUmG1Bqb747B7QVHTRG5bubE2aL4K1AJuzKQjizLJVY
RVReX8bdgSlI8ygY6y+w6zQ5nX32GZryI1iHklUVC+PM9K2YV7hvl9xsZPAt/fRN0BxhcQ1jtT4V
mdjzKWF0uOZmZx91U9p9hoj/R/Scwxj5lCXbX6O2Y8/s5cgJkQ07YlPl6x+WrBQGrk7KI9SqGeiZ
IlY+iZ4cNZtsbw0+7y0AkAVAWrHO0WMEEof6rGzbW5dg9iBCEGnVKSb1vLzOctFhwYJy+ZGnMydG
KrBXlsyS1LzDT/Z9qJ9dbyuusc9LPIrf1iZChSLVN9OoF7KH70g8+CtsDkwqvxgiyciZtPG+thCh
v5Flkh32BukKA2ffbGb68Pb4YKmw8Fr5fQgXfZKEPF73CCGo4hIMRho2d1srnN8TzPgTM8s4GYeZ
BrKZ0ROk3F8KMMF8JHopylMjhJxu/Wf7tN/amI9OyL/MjL5uFiktOdDD4MzpqxvvIPoxL9mvEzeR
XxkMKpMiIJF9pzeaHE4UCAPaZrCP1gQzaWguHHfndoUszQIO7tUNdUxHLmKTCujkrFCw1pdE1WDv
Jj/ZX4pSAYBaopghskHd16sVTc0Tsd5vndBZS+V+UIMv5xcHDwx/ZsqOugYQlsXWi793LVvqCB0p
g2jQ7b+KsWAqu0yrrmZTmZWEYLGFRcs2qfK1Zs3HAOwIdMAItMzNnZACDJLI/O3SrOJzbGz0A2/e
pJgTg9G/50WQ9sq32zAzAG1fznFr5zlnezpcZu7hEij0VQF9vqQ+NDpGxNWdAIrGqEqQWPPJNDH+
ESTlmwazpKAdc20HuAeS25uN73Dn/CzxMcPm218X8X6nYXNpzjHYtRusaAnBKrQ6QRlL/UedGg/5
Svg9oWKPQKKiHKqBLnNG2pWQ3mtxVzJMAGaBbezsnQ/C+GAlAIrJBfFWtENnduOtNuHAKGQLLRW2
fw3A9OSMNdY5ytZyED2wdObW0scnzIfFlW+wVj6DMclN5b76D3dhSxe4UFEDbl1jvtXBiS1CwINq
gyZGTRDCIWHrdjojILErAZx9bKswzcAMNIAY1rK8/c3UGyiw6t1eTnOgCX4BZDm5tfUs0lAVGNA5
ITFJGyxR7Gv7lDSLfeSHwJHFqFlEP1U60uJsgmv/KRCirV8WE3OzpDpYSgKkNMIiBW/Ue7GdoQEL
F9mjm2Kt4HVURZFjHF0D010RDiyMjrvNLYHgOZVw54sTu44ijn4cHfmATHvXscbxGqmic10mRfFD
cdVHp33R/yadc9NiuNdzfD0ff+Qr4stTW6IbGQhnnMZiKAPo6HBvBUaqLAYGVBT/2x59JP0ad57t
1Be/heSNgieD38skqdkxI8sTgmB8xSW+ICpaJcXbnOm2c1wIFVwpol/Ay6UmzZ+qOAHIXqrIdC/e
qy8sN5sECIepcapYpj4vvhdPFyBuDSrKuKXir09XEz74R6tmwwGFY9dYNyB4PmZ4aiAkY9v7rhOx
9qGMPjJD0RHXCFe9DYs5q5GKVYRiTzJfSbpXiGI91cQMSWYpqrn8Odl1y+lKJkNf2mgltkTRdaHj
Rm+1J9q0LE+4jhaqZzYuaiqD0AfOeq7KNwxDM/dBhINmlvXKOIJBAExx3M86U8Xg+9s3g3LlJP9+
3QZzxtgVgvTTKidt08VoajzeHG5sPwKoQQgUGPSP2H2DD73OtE8Nu/VCeu0+d69lAc9QvpfJPni9
S71xebZCaCmQLiVFX8WJ8r6G+2NLuf9tzBcZdpV+SE2Q4X1VqpIZvgLLQmz9t8l5LsWfH7wOCsSr
OexuXKx0Oc//esNqELLUd3q9tcM8meewhd3pjlhDkSoFO6+yHWdR1Gl98G8MKLEwwLTpbEDjN+ZW
AT6uS82EnXlKr1yZnNHurqkHBv1DGJ40d72TIFe2LC4rwZIKPRcpxtJGwUNUFPa3OtmwkJ7Ad2wE
FVIbYuBu3odxmCip45nnA32ysHfwMNA17U5ih92Eno7QzhYsFYhYgaJWz3W7EmWZf/fYTMuiPrQl
bmBqpohd6yIIwOV2w9VDmTSMcF1PYP3E8Hne75hm+273YRLIdeIGKs+3agu61GBCYZnebZuUE2QN
2CpAahCwkD5x7FBi19Dc5oh4tZc5flRt5wRahbIlKc93I6gPpbdcfXMXk54DDRRtYLhgzMyfk9Ex
l362he3sVo7SG+waktSXgNPsxnYCql4uIdpXDSOsyfORNW1wmxudq71KQRBgp/yl6nOnpeScp8/B
Wiw6pED6CdGvhh+pKbc3IM0vQTTyv1pKKf5wBn2Xs6T0dxzpduJACSrp4jyhdvjkx7gz8Pqqq2Ag
smzUzxer8RojD/FkNdArDhOwHaikxn1Go0u0ufOlpmiB/G1dftgW24ILM3UWLQMyR9vQmOYp0Gz7
wvjyRcj57NwHu7xDf+d+rYFa/5+nOXg5X9yBdZSVZt1eb7fUY+MM43NoOSE4P10yBb+CXGvTLKL0
YCtEOfVOfZu0Bro75drwnVBf/wmS1MmEZ+tkrKzhC4ED35AY5CAJ7oqYkAzHmwd+Fi2cAkN0//Hx
XtZIRIc071M6YAS1qPQGNSkZJ0sRQlIAvsuLd0MR5EBey0pQ1KamcGDrLHbtpW91O5wVuV5gt98H
hf7ki1rRVCA07+mMMBms/7LjUwDFsyE9oJaz0e+JuBCpqxQyWYrie6WpnIxbzMhVA/RBD3/VXKBu
6q/IgZJJNYHAwj5hU+l9tPJOr/bgZW+V9GO0Zs/g0OjgWHQHFgCRevgMscw+D6iOU3M2JpYXgpvO
Woga/GSZKiO9s03vUrwPLedVTgA7OzaoHmjdJIYdSGUwnUnDUmKuk9LMNYX/PFvnpkonnAyFSLi4
AzflUHNhLYACBhfU/7yrbR5az+Knsnpd3jW/RgupXA4RwSPiWCAifsI9SwMyP4j4wMWX9HeYl0C4
EJFX+dmyBp0MtqjA24vamIbh5XKfhfQUvZPMqjaP7DaNA1dtWCuVSGlxxEa1RkznDeopq6RYQeE4
NzZ97XDRJgiM5qUHONU7xXg71LwHTHQRx3e9iuZx8czvKXDG0fjFQ1ZHUoPpXrOC3wJAyuM53A9i
0l75J01UAMEQPYfdK4fI2FBzW7Yn9QsEF4HypI4DmTnNp5QS7DF3jzkp2JU71nJs9G+MtOnAOecX
nc3NhRKQTKqzkpCVKryu9Ly1k+88sNHK/s6ZVdY6u21rEOi4uE4EFY5RIMfmDPpS5Nt0Dd6vvWf7
xIp2KKfMI2D0MYPQKItK2iDVfeXI58yFiUNx2Y8p5O6OcBrB1e4OKwkrjCkhTkgtyjGViu4ECh9C
8XRL+WjEZHLIROZ4E1SeyeFtEhxgrRPzJvn9L5cAGjCLj1cTNcBSkw2y5sVbJpQxcrc7hDIgTiXX
LxjfprJvQhUFQLY1yceK7AAtAiVUKQYMlpGUt7uILUT0BP6qXuyrtmjiIpddFc5aASN0OxzvPZl1
iq08w+LlHrRBlEjCHxpC8BnfIExnuEWZl4ZgXa2JyiwSrU4T/GakyANhztJ3IL11iSWtq82+7Tjl
6szQcogWekyfV4X3tuNzIaX9n+bkS0hHjAimS928B4eyixZxCs8rLAjiAtZpknHvu7qM3S6Xg8Le
x4OuFbb2LDnKugx3jndj0AHC4NJdfn/8Uadz1DjCQA2psiDNiYgYMuPuyIoG9jIpIBBn4H7SCLlX
q+f1jjyLBcrllaqpvXrXZJled9E6ynrWXwmAogNOszPCWkfKMOqJpElnxCG1VVxsgkt/AxiOe+dY
QKALEL9jVUJR0vQHEy3kx4etZpXZPI3sk4a/H7KyUdmvpJF8YxmqpoRrNA91ZopjiLagq8RTkUf4
VItM9QzRgiYTjX2nfKiK7+i1/hoR8KgSa63w6b687YCDNYbP9gYTylCDg9FfJrEhSgKubR4BoILl
jHF822YasWXFwXG+KKmA9C7VSZKHna/G03gcxooRcaOdh8t5Rh+BwdBI87zTLA8uiKrXZdWfF3M0
0jwyXNBIrTTEcCR3dMtI87Tb7iGZcvs7S6reREYO8MVdm3r87ytwOhKIXUMV68fDtpSk5BsWYKPh
w7eBZme9NkguBMYvFyjnP6Vf6OE285A704QxtKihwdXozCIfVGRGpr3P6zPLW0widUmun+T2DEri
y2bY+noLY41pb2czX29ni3I9hOeD6XpnmtxLJJlQD9O2l6GuA46GEJA+LYM0kkm1bf5vpnGjNMc4
c1QNR+66dhXL8Gz/v/gJHurDyIWsJNSYCwN3bfpyfzqdFx85l2WvKMhKiq9rwGcZO2GopZZ9VTdq
nw8yiCKiR3xCCllhXPi837LywrPYToFem3u4ieb232OfzgyOboYPJeuDF0GhLtKDiS8u9+pInU3i
SPEbbNKvVMWVxotdZi1OBw5zI+CXXsjZTFl74jlYJEqWPPXWkZck0yQvRImlsyalCainWxKYSFxa
1Z2B/dymCcUUYl2SuqCCBJJptQh1Fy9fheFHUsZybN250ksyeHph/d3VPoCy7QXY+RrTfk+h/vXk
jNUNRx+gtWSo5Ij8bDh3Ew7KEizu6Kxv3MC0NtRVB3D/XVTax23+4D58g2pMo5gIEg8D1pQLaCJl
rurp03lzXOxq7OnO/2FzX4zrBOSmaM1drMrM/37+svEcWmicIUUZlJODH/jHwF8uXRllhNl6LF6I
voySFHa17qap0r6b7DvbSmO04djOEzLoXfx02UkJwXTr7ffGBNShfLMNt5cMB+1HXsi/sKnMa+l+
zHTCNGcnI7GKBfNnGAGASrRLSadR/3igk73kJADe1OOgSzUW1CXQBqPzl/3ohY38m8LelIj4WbMA
qf34wKpsQj0k15k/bXG7sPnwmf/cIApbfTbX0IMM/a8iZ+iXqK9I47rv+oIlbfFtKE1f9LdGNiyM
mzSP1GrweyO/FCwipjmRQqOA3qLtnKQhp9DjHkkY1PvgnWuLRQkoq3nrhv9FVHeYVQMFEAzdwM4A
sU8ye1cgoGx0W+TMUf2F9r2+CwmK8O1dmVuXfsex18GPVTpH7gbupBzVJ5QYkU3BhD4cA5SsG2iz
RK32hmNtXHV9MJ+bINxcN6NQaWlNjaSO9SotmMyORR9cmZmTJbOu8NY/fkLwxAkfvh48RB7LmWZk
JObFiVncbDBe6XXXwZH6TEkR5+6bMfNVFN6mv/BTTuHqEnQvsSIV9ct7gbiXkWt/85Ml+FgvrMfa
4UNTCYsz9S5JRgk6/irQVSI9yBNBwUiYkVNRZl5vLYjwOvZD7dHRWCUOUDOTq5+c1SWwL3MTojks
HLBz2eHE7Op8zahwE/PQVZFBzhZs4kJA4eSsBXH2rqjafJqiz00auGX7nSC7gPUaP3451YglgwvF
59WFlD3W0s5AYlsaTQoXBrCCwm7njLH8amBQe1YyE90fy4Hj9yDotqVNt2pYOkSt7fPpfKYNxBtc
4Z7TAPjWmddUu6kVFyqTh57HeY60ULrvWmxm2M09lyDVrKFMUmxZofmnjp7+GMx2aq4jBKlkaviV
TDRTdGFM8z8178G7T9UUK9a2UkgOEKjBbtggyu3+mfojLw/jyMnOQVpcZTrTLIn4s9Vy1Sx3dl2T
y14+9mCqdzX6c0kOZSgZT0WvkAjj+o2PNgocVN1sCbtacS2dPkWdLSF3R/DRWWS6L5TMYGMp8LEp
PwdUrAM2W+JSLT1bUliBHBr69gczySglUJ0ZHXMVkz4wsiorC+kBtIClUCDz0+IvYL5J9ocRgf+y
qLeb0A1v+y+Vy23YXZNXrTZgKzXAON7wO7T9xXxgpqU77oZ2ATyxjSWkyVESCx3IocAwox0uz8yf
MDh/ofQos7UF2INwDlDxTkyGuhjJX5gpCxrKoo1kSuNUhRjiNCBy8kOU39oLJ//cDh9ihhnVDfM4
UZoNHqH1WTP6nt2q3nrJ0o1EE8nJasBMMlAfRCp53nvdP0DYAo0k01Ji6YOxQZbw8hHAgustcVCz
N108N8y+FjOkLDaXR1NffneA9cPJljim4j0wRtJtlwivTE7Uyq/irJ/w+1elbQMVbWtQg3nm4+w3
kbcMmVW31rR5fivc8pIAgHfhy6k9/HATFEEqjYfmZ4bcm/0gLf8KBUNl6cAcRvSahfn+sUAkw1Pr
cTIfh3hUsNFX9vTd+rD5QeDs0JdNBbg2oTZMN8G5yJ4My2zNabjiyox+DVFD9xSGdANL+N7OiSSf
VRXzsqxx/iuZfcv7kjwEMhuyLRzh4vfdqunR2XGwOy7+14Ce55mQ58iusZBxEJ/Ul5H2BHYITywl
JzmtNDoekaM4Uiku8fzHZv8vA/GUVJs8AtOlEoUEkiZeakKFPSDXiITa0PHTYY6/DHQqOwsifLea
vfg4qhlv8KpsqgEkerJMlw5wBH6i6E3q76tSUDewfzXFD0JNH9+a0j4WK+aF3ZxXIcnZPlnvN8oM
YWz2JouITn1Lteo1YWUOYPMHD3uabjQ/bfPNPCAHRUho3djbvk9eKlqg2p3i9A+tX7QUxfVpDcAr
05eYudGzbmGOX0q0x2Sbkcqz6lH38phQWYxP7Rg3PRWxk8agbJZMhRpRVEiOCeazyBTx+UwEGZzU
ngIwBKLuVniha8A9b9ka/dpQsRy1077OYhopaTWJoO/1/9QFN5wn+ox94GUncnHnVhVHnbb2dGco
72ZwhobrTHhcDzCygei99BeY5hT2QjFPpSInn7NpIu6hAic57eioctB/YyI5yXpow5maOpUWozeY
5XZA2D/JTJEwsyOD8NMO0Nnq8kRm9n+cqAPkdAuuAGBjkKQs52NfWh1XCDJ1NmZd7wl41C5wglip
7Xum0wViA2HQprzB5WVP3+elXAGxrjzhQl5dJMh8fo/OME5T3b14R7S/YxIEAuLanoEJr7rrF6n1
NLzfQdVur2vtyhtxJPJIL/aFajBly9ziRNtIMeHFSzJsEdE3qb2PcAEKM4/xy7zkRMIcsnmABXuL
tapzpHBbO9UOaFeJop/82cEbdzYLEntGT0QyTy+6zOB8xz0LO/L3caVXOFRxq3gkxoMgZumyeBO/
eRX06HnR1v1vmcqeT/smg+gv8E9SzeQSBdJDhmgJP/8yUgeVNcRYU4EavD1yS/r8qgBjRAcBqD7J
NxdJ3pTxnTNUvbiCtJAT95zjj06zod0uOYfRyAFdgY/1ujGp7VPgDFrQN8JrLhSOsff/+mcHmpqY
ay2Y22J7B5fPzyWdEL6B82tfAluwbZmvA1nuD1wQDZSuQ6yzVrfb9Mrmv1Bko2R4Qtnc5r04hUzy
y6HwEsxmSMejRwrByi5F0eWz7UfIh+mlVeutw1KiRZbfyEnr2T7qXMXwK++ag40KeWgiNUt0A6RX
lBjsDL+5Yb8VBABk+khDqDNKJ54GxLt43QHlX7IbnFaUUZdgZJJt4rELTjpVwoWeimbXlqVLrKVL
WZWbf8g97Sg409siZF53TDUkn2icFRsph81ytOlMWjdvyJx2yBoXw52lWAC1PgVjylfDW9Z7/XwL
iD4IwHz730Rndacn0QS728138i6UayT+WK7vyugn3ALjMDwsKwFPZTsnTO8JfRC8LJ5zKiZnAmtU
BJK5Xn+gGxgsn7Da4GDELw9H3WWljDR1M0TMYicmU9rxfwcjGnWKG1pQ9Tsww9y+4b3wOE0kU+0c
Ij0ShqrtKi+j3wpxDmkgXN5hpwzTLSgDnBBd94gcbb40vZJnnAR84qMdKao1Ih0orBpP1R7jzpcZ
PX9EcEWqZnVDpM+iVNr5sV5uoTsEt/nyRbO37pcmpFsJZDQhVrE7tuWmfSWYhwvGJ8yCMPA1/1ht
nIPodzAyWjV1WAUZxPFX5JfJDm8mGV13r4g/NgVlbg9nIbmtyBsGWeZ63ZYUJTODWjFh76eQ2zbF
c2BS2Jxmg7f8lD8n0xviLP7u6mVwQGT6GvbpAwFx57MaPnpUsbOwu0tvzzc+lsy40bRJM68NM15E
SrLcg2o3ZfOKPxG95/bUsuV+/rJfW2IW1Uz0L/iD3EIFxYrfFs2Ra7hdoW42uHanyQnQJkdKGtOQ
O8FoSDD2oK9GnkBWyqpMcqZZln7sa7zpoMmwoAVE3kMu6CzzjsfQ4tuj1SRF7oZAsI26JYXra0sW
+DvwOqGgI0NjD1z8CNEbHpAPM81vmMgCXwBbd+lIKZg18RpSfsCOymPEpDR8IpeQgty/B3p89XG8
iRv0ROtYGVAz3FZWo5HKdyM76tSfgPsLWUYRUqEANmX/tftV6jZCAAXFHWarUpxaJqzJzenkH0En
oIwu+XcGzNjEnd+HRL6G1ycJzyccmZ9xgSrYgLR52fTEvi/as4dWt79dgcoHZyiUsooRelFuRyHC
hBiHe1Jv87KecQvdh+xDMG9H42t6aKd86UNfjw0GfUdP1Aoc0EAaKwesUii3zQduqaMWrny0wCJe
qVt2pvk/0gabcN3lsK7CPS4ibR+8qwHOs9ZP3rLxtqMSx2ObIoXCTMYQYBFPP4VJH2f9VYfMu89S
laNgTkrIHRBf69FJAsu6cVLLzb8XU4l1WklA6Cf0BmmHRtCPYmQ2YptE4qqiIAeXlMVfkONkrhhx
Obw/G/TxY3jnYtcYt78wKlYSYHZfTOqv16WQa/jCaJhWj9KxU9dnsvosqtRsI6A1BRgCYDDqtwwM
GXdU06FxETLMB7C3HAAZS9kjvx/8gGvig8iGkhtJpwkROrzt4fRg9E0ZE3ZES7MgA3O1EJ9TBoDi
ovrQwUaU+WpfoFBnvdvdJgflLf8O1BouiZLQ3mKAYbAVg4ptJ1jNMXyT8lcKI6SvQpMcXmsHWz1l
n7UIsIeOV4sYYuDDSTEQJugRoysceh1hvJwgaMOO7TBLuy7IV3vfvJNO8b23eNdRFDaoq5RMbbfy
o4x+gJtKRN3i/JOGXwptYUj++FQyD5l2CC3xb+sjfaWymiJC8eVYnTMLqByxKKFh/zpeIXOsnyzZ
ayvakHSa7B7iWy/ZJBK//AD4pZKiwGsmMfSMkFjxU6SrwL3uTGZZv9VzghzqDTuRNkbsmPmvahMW
+CZkA0slprx9ClH5gu9/U+hDdaP+8RPwLxku3kCuOeKMxaNm7juLButQ6N+E6Q8m6uvyqdSAPEqy
YWJxnCnwZuU1sJcI+HTZJ3p5pRV1nnY0m0s9gAsYlI+ul+CSAD5VrQQRodaUPR0flf0+plWgOY5f
+V2nNQtmp/v4JYpD5apvcs8EnQeQ1wTKg2XD7F5Nvfz/Hoz1aXnq+fmnmjFgGNx1Q70pMFyleSJb
fyVENzP8NN5ijYcUsKPaYUd7vAioYhASUxpl0BCdDnveujcK+/+C8ROTRPuO4cvTAHybCC9Iokf/
H7nXoI/9pbzf1g3KrSXHTd+qhgm+etAo38uesJNP/JLBoku1DB1AVwNT1muiL2HES7E+IQDvjihR
Epz3gp2JvzSs2iFuhYzzs4ZPwzzgHHzPWoExPxmCp9jUSx/exnf3CNXf+Bx0D1qitzaDfH4XAUG+
/2S/yM/PT97xLJmyFl5wBIhPVDM/Zo1UaAmorvljpXx4JENz19jsTl5Ysh7StkItLSLqdJVSr9NI
gqz25NCPfi1avwT8c8Y7SWTy+kWi90ZB1/m7bqJzgChEeRHdv6q/DZI18MWgslD3ojWQJ664t1ja
UBaxBN5jVwKOIgl2l+kJjOjFs5rIVTYUaNrmmh+QRqjgMhF15HLOdCXwvEvnYp9GOz75X2gNTqev
XZGmvDiD206/ktcTNcTkmAAg3i3D1DvZ66tYbYLQXF6cnMKOM150iEDEmZQCoaM1vH8SdsMT8t1U
NL9yAUA4CmFtuMSwmzUhqyZ46U2TWvb8cg5pIkbwhy0CX0lM0UrI/XEAbh/fZeqkmxLsUlUirGIO
eCHGJRdUe5nmKr5cNGBW0sKP6mqRTcq22sw+hfwW9MapArt8U/6+j2ovdzhDZbyWJbBfssSM6cLc
O69vbbAV53DR2ouxH9vzx7kxm597hbSzwmbsWGqKx8JzXsKlg6GdlDYj1OQbctDudMUIutqRy3Wk
aAk4Qojed+C4U+bhPD4Hq6QmHzMN7r1rplphSOLfoJpJVk9X7Z83Fx7SMXCSkQjg94/cAiJPck66
dO1UUb9iMz3h2xYFIqcuXyD0sZUdmmMhiafArYmbPPKIllrQ03x7MjCp3X2USGVMC58vZJlZ02jb
3Xqg1s+KLz59vLGm9Lqkjsti8a1826HbI7X04hDUBoscd2tNazmTYifpXxcVIExLnHVqMQyBlAD5
R7pv5DXBWF6KYeGjR8UfA0Wl6IrCftNWf2LxklXp+zniF6Jwm/tJw6l6KglQz8MACwdo5xhH49gU
cPQ5047eMiB1Kjj5IBPGYok8+lUPs8+QStY9VPzE3yELoN6DqEKEXCRSjicMBcgwIBWRIDm8zOQR
HxLRIWSyXx4KLBhXJo1wWRVrkIkhxqD0QENagj9qbVqGTMIpm6Pap3PkT/soN/LoWdtITFbpQNPH
CUuJta8KidJNJLedqlmS8xZAnSgg9uDAjOP6i17sKOe/BBYCbmU2HxT+nysrieB9+015KFqETQ3+
Mc5rBbqgHY+PvnemshLZVzZ9QpbCU9QIIRwWokPIYWFVICoj13QjXt3bTUE9ZSwWlTr8yg/S/ePs
kD3UMH23abaHm21XVPApozNBgAxladGDBQmrdZz2q0C90Cmw4NUFht9OSjKFjAeGfD4JMeucWvYV
h3iQ/DSp+nDIuD0yfLJISBjHAFgfC0ZNcUQdEhV547iDQoIyHKUZAX1akwlRxsD26qCAE9/jmBL2
+AfD3xyS3Q6S8HssSb2gZXZ69ZiXtEWwiRSUF5+wnKrJMbn10+IVW4AQ9rnfNkU1b46f1VGKJH8G
HgV4y+R0djOM0TFFljd7RPVQSI/hV65ZQ6E7QoQSl9ietwQ63GeAf6Ffh4jBumQ3A4UTPZn9x8oq
MREK+LaRKR+lTQGGGw+5QFjUGGagALmVggfXWtXCFO+ZSou5x0/lcRjSjcyr3hrbzLEcdPLHsfmJ
DYLTlTy+iOGiDGEooBrV4uFamnZ1TA8IalQ+Vs6Tl8p9i23XBFeTHnTiPgSg3LvyF9LhHKIc49oZ
iNHXJpXT8+e8eekWzkUeGc4FhDax+a3EKelogb8ZVC/0XNhgZpzPXbyX8N0Uj+BJYapxxxOMHriT
WnaZjiLaJre/OxoIy+Eup6vuqXjrfkG9tdCU9+bm73beLVEgJjXeOUR0MdxFgU6CjGlgzVqlplTc
BBTpX7EuW2I/Qw2LGmH+JflCxQTTdG2tJmq0FLZWIgP+3ADbkDcOmJW7ON02/z7YpAh8gx2Ht5/c
/0NQA2bfAlcXFbdvR8SewUHVIAIhm/rSpG4Gok5pjtoHKO1RNBcMZZNTYjnx99PxnuFBDX4UNhPL
5P6aKmVNj4pZTf0YDxQYxqL8Pz2xjFSfl24AulfK4GOVQsXfzamN9fB4gbsHzn7dlGnSFTh6Vb3b
K4U0IkT05IqOQT3KAtdYhH6oFHT/63TLFgokStF9pRBVvs9G9gfg6UjGe+RFazxKDdVaS2Uc/TSh
C9fnniS0NElH1/zgHHk+46UonSBE+L+sHknzyLP3KDbrSXgfBugwBnXBYmVFhu3wIotCPUj4inMS
KTjL6XYnmu5xdR4ylbwuP38MyfqsVlpgRyR7FU8OODyyGFtk77xkL9o0J9lrMOi+Jz0mnCexoeHz
/o70qmuJJRmi+P6j6fFJK+eLAKxaVBLqDS2G7eHBRm7bsejW3/VBUcDS+tCZSEWvrOfaOr3xcbJ7
Pp98T80q5W94hTmyLGkaYcu5aMkMv8Eoehil8+wyOfluMmCkXgNsqmgub5SugD5FdIyrfBDtCKEY
ss5j7JEr+I0j4vCdP1cAG37rQ230bFBIzv0WoLDSPe6yHWpOXRIcjPeLIiu8cbKwKrp14AETV2jB
Qqe7Exa+WLtcYz8oJEQQfic58E9D5n1hyPYIP2GEQuYbHUeShmwYaA55VFcEHxn66Ocl8NAfdl9j
POoh6nwsy/+q4GpAX4SFHzF039ve6ezPH6fAP3eL5fxvmOnQ9O1qElOkTltgW/NUjLjEiRT/L8jk
iQsgLBVUQrngU3mUolRI0Gc55ioXXYmzSZ8WRR5h2H93hLr6ujvfoc0FejI2fnMFgi9ho/+XiS5I
Sf1oQd5rmNAW0/g1ZuiVzFlyhkLH832VPAV20vyxA/rjRUEtqlAOEDS+busiZVCgHUlUSw0L1no3
AOeudZrft0CMFjDAO1TdQkfZLTGcdglEouKG9DdsnONX9wLdmQ/8MeRVtZlWHucrTCNq1Be0Axhi
qHu77A8iNgyGRl1PGbNaD8TmFUIHZWUAh9sW839BG/fR1XukzNSS5M9p/c3faFZvGZWTOlbAvJky
EI25+doFWizS1uVv4m8FnsUy8xCfI9W33urHVPithTs3wZdH/Q8dMxZuv3v3DYMvNoOeoiNg8YjP
/pOz4QirkBFb12FrGXK6VcZpHR3LVphzWtei2sL/ftirp7krk28e8FSZqqYaTWFVcK2XFXfkp4wY
Pse76EumFpH4ZHVuDpnzhh6DLXvFL5CalEq45snEjMPHuIJ6R0LsnyWMfL1bWnd1oNi2B3nksY9q
idPJ0tFTARlPI6qCDdr+Rr2/yGJI/6a/VRuZoSCl+I/2iUFm0hLqssxe18qWQbrHiCMz/itLQMeV
UjLGDolSimU6ZQa10dkUdfjElffnQPgU8jyAimWuBuo/yNbTvsz7ROIUj2kgOCQ5cu3sFSU0+CKs
nxu2YHySBZIEomxdXBThTT7oRhd9/ynx9oQillDl3GJFgvb1czOj0RYsBKF0iCaECp0eSbDT351g
BJ6ayiMKw9hWPEqQFMaG3dtxH3boRLSTWLcShZwyENlby/HvOXbzp+enCxoqWH3WhDdSJdWJAGqy
y8Er57kwaX3VVL12+yUzfaJD/TonotTHkxXCftWVIkvw/f4xHvG7ednbH8t65c9CpB0XK0d89YkL
/sb6r/DW6UqsAE1q2tz1fb2CL6cormhJcmpW2WyGUJ/8gSwDCVydYqHQKUNSCDtDYKkJPOgu9cyI
vqAo/l7p0WQlRTTxAXFKG1AqmnnYvasw9Tm/EOoBhvwSUh5xTZpawCk9deq9HNMU6koiVqTP/YRP
Fs1r16z5h9pdykcrXC61s0FHE8KCXtEvhVHK+YP7JT+vayiKvFZXLIQ7k9uGFMD2yNMGac0DZGdt
LAyOqDuxIfwr5C/784mjM6JHD/raZq0uozvl08heW9KEe6q8Q+Fnc6NCRg2WGc9NgZG9+t35jDsb
3f9cA02gXIMTeY7+X+TmgvoG3U10YjM3YtP7SpNhWYGEKzqzdml3+Se98uwDFnIXtdNjApV/Lon2
K3cNOmh0A2EJ/5iyBW5WjoY+bZbDybxj9Low+TLWhh4N2ZxCfOl5aQ4yO6NdMSKDiguGPO7srwnC
yjs3E4VSZA9moeycD5VOnQHVHYJ6CyqYyu9JzjRzF+mPCmWIkf30SCygsbocC+SG33cGDiO8ikFQ
H3QdwWddppdyAXeHnug8HgpLHrlQYO7Fubmi3yfRHF1cnOwFhAy0FzvNMW5FRrCMimBBkmfjK9UW
Ea5MurHFB0KZ1Yseo/WOOK6J+kYCnOvQsp2bP8J7KIr2KqJ33X0i/iRZgH0gvdYspBPTdPTacnmf
L3LznhFQ5YrQMShHjjp6s4ySvGmZwYfsRmmvIT2ONFM66lbSW0mScmSZ9STlcsxjOdM+T4FHpSQj
zAKWSKYmQwxVY9cYGI5EYCleqNiecDt8Yk6doUcbnhe2ihEKDJxfO0VBfy3nfqX42cJbYr+lcLht
VdfkZ11iGMDT7ajlgWogVsQRS7sT6mZ6sMEj5SXu0LwhowUgKJyUVJ9XEtQcgODkaDaDfRwKXfvT
mOzrB9qnIaWfSvEVBy3rSaHd56pO7+TbjQatGx5qG1US61tavVAKyWIBw5EYErXlZe4JK1tfIKmq
/TfW54bolCt55JmFC1w1LPyLnNvSZUEtA33CRLl+aEOr48+pReYoSMuQA3Q2dtC9qjCrzmUd7rM3
XOZbRFen8leYwFrBVia1o1WITWUb0ldsKYDKQVjRIUJri4VRF2Xm4HIGFTup/qK0FSRT4OqswYPp
D39MeiX2uzV93PigXk6SCXB071tNFGmWCwTscJ9VE+ZIwc6OAwUqrZrWyZ00ph7zFauRLPWngBzc
CmK9sBJn4sd5CV9Q6r693GN8+yU8tLnGe/dSCcdY9601w04SyonBsopk/WTn46xen5B7dmqEFUzw
2vcl1l6b1k4merNRDg/R/KI6V9+q69Ox/QSXGQC1rN4/hsBS7YoZFXtQG/EobaquGUNA6gRvlTLn
CdS2veBos1ff53S6owWzME5HhEIAWRcES2vJLwt4c4mrvCLf0mlu6k6G4gA/RwRxMpemxzXHw5WJ
6gQO4r0GGXywfHnwpHwFK29PyUX+pZY9su77Grtnunopx+BjVdBvSt8D79hsB3vMrxJvgcqQJi7o
Lzpoj7cyS/OpCIqVz6Hp16LPQI0duzAMqUEn4gpEgejXoZ0Da0nyBX93fEKEGNxxapaaXmzPB6vX
ovsdnaerOGi+GDVUMcrOPKUsI5uMbx8g0RBEkPLsAueSCjislCGrg4cvJ8/QJV7xhmj7qlh/EWmu
BU3ZgLyID6FsNFDTM65D/83X1MYO+Vni3LxTJ7prTv2c4OIuKZDWB+Rtjoj7MWY+C0j+qQewsFGR
yQL7psskPkAqinc1tno3MZbGGlNAoEk27+kGW1WHq1EAilJ9OUn1xClyV0W/lbca4LQ9ePEWA8wO
z544YBnl2pwgjR7jqID4wqgcePmcS0J+8RrAhxvfsgdYwQdu+1Q7PWeU/8PQtgBwxrBPsoTuZKde
+hb62J7NlqJF1EW/KoymVNWXX10wVs0ybIH0A33Vl2MzWgDvBvUdbi1Y0vepfduGL0VwGuNNH2l+
uvSeJDqmfizh5xPQjsFeiGMdOULW4FKSgIrT2MK3Bb728lB1pNNVJf+RsEXXkPS6dayfdQcsvuS2
46rZI4XpMf2cYYluhepH3JZcgwWsGNvfjiOTvAiyQyEH5b5f2edyn94BCZWlyUJGuX86NKSi01Zc
M4dWceD8SbRWqXrtepDzMfvxb/UpgV9Oa+V3OUScxtX8LPJnM64YIZk+W39UWcmjznEX+V3QaM87
trKyRT2UTKQ+9gzliATYDg96+SxemMSwztdu/K5KJjKN/fgJze1O4gHJlcq7PavBnhv+tRjtI04V
uFAQxH4uqEu83Toev2Hqr9Gq6bdwcmEQ3EOxgxR9r9/rqbd/M0aFnJjjW0GDnTqLzDbX9ETKAVJu
2J6ROSGzPuBgC6Ycp4yMYSkUU7WUj8LSyOYPOJn/Cl7PzJKhCfKlJfYinXmZQNX4/e4weZmpc/pL
ayJi6UmHd+fW+Ykwl/hSicWXh02SpqrlG4+W1hZtYvDuNGJIpPiBkDH5lkfWYo6l6yxAcJLHqu4s
LLhxNqqRM3396+ZfESD6FRKBCp+DZadnVgDtxocv3TumTcwzRkKyNM4LFWmLeJq1WQH7Y/71yR1q
P9wjFi2BA1FFAcPPJ3iW3YFPNzmb1sZEcgHa5escdSkLoNH+cYZUS6LgWXmuXYyj8pMhmt1PwE4k
MsZKdnQrgMf3N506+DGaZMP3QRW/DEHXVwWvCXDdhWlu5fXBo0dmpjQRGR8Q+XYK7CuO8AdVdCNn
w8CwicNwaxu4vg5VfZGrn/Rf+MTRmjOaQC6WME8+Y8dJ922S07QPBYzkug9Ny+vm9SBhBfznLNrk
irlc31v6W9j9MOPbJhAJC+84hwjLbahLH+TS98WJ6DKBauT8/KZE60wr0ssMJt7LvNKfOCzYTSd3
wwWo8+44oraBYW6/J8Wf+ZPLI2Zjj+5tX1by3boxI//ajzNXBpaHaogjC9yRSgYzp6+FJb2ndte2
t9DCGCyeEVZlTw6xypQngnWddvsIXl6OBjlIXYFqoc+/UGxWQw7VLlrIcYfl6Tfyv/Tum6jao5Pi
RYX04EV00rFEguO8YUs/oNduyYdNEPqgqWNO+n1B9by8lAJG2nOrfNDJQ+l0S3n5SvCrkeQH+SUc
Pqb+3f8KH17s13A3c0PxTuDMzaHaoGLBiqvF2Uu7vFsf9dWI+JBGL8009NK/4bdHaksHUhk3ajOO
hpxtvRdPgY/tzL88Id5OpT7OZInYuETcbD29mwmqbts3bkx25wGmH0BlfYPn6ONOAu1OQM2Dd8jR
eaB1zoMaS3wfhNKh5iPJE6YHq03qTBuNY6bHUsOTYnpMnc2MJ2A9U8e2YNcxtikCpnkE37C/YeSP
HcsJcmPoMS/+PaDgWVZWsGcGijFn9K6JkegzWx0AuVM3SVKPxjCknJF34eEhzNUhD1Olv0biR1LM
JbFc9y619OFiwcBmDB+dE+cy+3baN9MZwpd31tF2BboicxoranZhsWorE/vDa23pVGxVpRqbKqK5
z6rnu2DftW4Pii4VU+eWB7kCOUSUQMdN+hj9XI6cRErnpXsXXPzqer3yjfj59QE9BPNX82PdPqtR
efhc5r9zPEAcGlvtHsqVIdfPsOQjcCpFwHSvQk/cJV8xuyreOfe091UGp5Pr8+uX8KTnQsuYNvaJ
pmStIEdJF3mGKdHLVCyGHb4W417tteBangtq/ijaRByGGU3zgMYH9M47E8ZnGJbRe67L2MaBPiid
3zp+0yJJXvy1+qEb/nE5UvEG0WlnOlqXz1o8qVp0mNrFs19hf8Crq7FMM8cdYK7aK40o6iVwPkv+
r6pexZlFf0tqFzdigpjYFO/O3HnUOJiXKlQek7PZASEGCoaCn4LcdXIQnkcxET2YFsD46PItUHSa
O3JhVcnBwfC5OcoQxxKHcKwTGMP8Wcdg35KCLqRLVW39VbNKnhkchlGf/6TFGzgqlw425JyhuPdd
GhnwZw34Z+AYIipg4FF1gaCg3mHQMfl4/4Os3ulJpzhpxjvrI2kNwUGMUWStcf+lEMrSDYZpSs5J
CuKN8PcJrYy0PviwQM38xFVztDhsunlrEfaR2OyJqSv/Zg6HCakFOobAeVrva00aacKEUJUZpti0
DLB9SAID5MrtrzWNMOK6Kb35QG5CMVV4F1dGHYwdAI4Cn2rQLOrGtpMOSxkm5ou8wwJSSmkJZzJA
gqN/8QhW8NXC8czxbk78IsG0aMDJ7SnbLB/oElOtw4FqSFs2BRTP+mdoW28nvco9ZtCYgWcveGah
nUSzBmf5a+8ZzoNgWXNS4Sv81ewF4Zpe9DLhibdw1rSoTH+7NPCD7Rr93d3oObvN9gCcVForYlKN
W8kzBp9BdRewpE0sX2ucCNYU1Mrym3CewvOI9GjikWlTAzXayXiEg6z+pKwz1aenEM9Gj++jWRBv
F6LqCDqTVlnkhnExiy6UMEGqp45RW0MBWHlrJNmsCdp/KvYjem4p+FIfmyxEftZWtfEd2VjM1MIp
Yxly8mgJxFXfhhpHTooFfPLvjx7SH1miriG8ZGbHPiwf8W+VwA0xAqqgciEhDTLhO5N++z9rILK5
dUyq899ojZ44aycCnrhX/dEtV78HPXSpTTlVP/m9BJegmb703mRh/ig5dEi+MF3JihbKvolVfC4t
MHIITuvF6EPPtYwojdhsnRWhkh/dI1jY/CtAFpXvjPQ5QlAS/Iq4MS4Mjoy6w416NWIMm4OiWB2M
DQlw+IuzcwLi/EHzNOqacXhDsFh3LpDTKzfqg9TjDe72QsoWzxOTmuvtxmt/thLb/w4S2w40N2O5
bjgfwaWHCsaqTmjf98pN7wKb2fSgOuQ2MbUyte0LOIS0fcZ7Hbb+jfVjtYOy+Sp2loJxaBlEW97y
LjaNzE5iLVwKiyCfAq/PCu+ULI6RsqC0/GvW2dVZRF5kxQ/MRgBsxhE2qGCkZsko3T+hQf3YZDyM
6Kl4USfpLsrZp7exJCXh8I7cU2sOkt0EjNsfLR7ouiXGWJw0JF/o9JWdO7mqQIU4/h2LCClsea26
KpAVk+LZjqygoxmjTPBzTkXX6YJ13mWVOCfw7B5Ezyfq/RYTK9JujuODNBd9E3qPLLQhl352tqjN
Kvr/FtrCxrStbDzMzuN6aTzPpa5qlr5Ib+bGYGTkGq2kboF1+Y9wZpSg2KoiF/JqoPliujbmhWi7
OQYr/wHHRP0Gf8/3PDyz3H/TAAi6RTCE2KzPoqaayAEPKN56KC7X8M3XhxKEH9U9Z4g8Bnuumofd
P074RW7K6LWy12aRZ9jhKnplhrmx8TxG2G/8EtC2lwJX3aO+ok0nmQN5UZKgoI8CO2yFdULo9skF
IJryOk+u4G9qCYYvhzDwoUgA262R/rIqxnPfLAVVmpIPqnTyG06uFyZ5xln6WYBsIff+O7ZVrwih
j85+3RTmy2RJ+vZrXjn+6Q3Ke1vhJvui3ZVKNwR+E7aW4eIBkpb8ThK6sHf1zIG2mKlzU8i1wt4j
eYX935u2JCRtRjbQReKBXCG7657JoZbRIVczYtgIXicAIFXz7fN5vFedEsad4Pw1oJmWvMwD9nPH
RQ9yT3vJWunzaPnFN8Lt2alVHbwci12GO1YjicI9N8/sLTttBJudSU7jBhDpn3xVadAuq3xeq8aQ
ks+oAIijmPLfp7lLhK8tWblAIrL/oCU4F5vQJnZKEIBESpolu3EfZ8EpG05PI1xPEHhvJ62a1acI
QNiy1xYDG8OOODT5Jdz7J1Qvvscklu3329gii9RrJBzSGni61aOj68tpd/lmdlp+lLHoWMyffZxd
2KZAnlFZg2bSd3dPhBaBo0YqWPqACOw/8cHj+QabzTHqD4NLOdVOmpVgDVrIt6d/i6FcZ5V11Lhr
vjxoQamg17umgI0G8nVWndupHDZAzMax4E7K3+F0TjX6ULNh+N/UwqHZno12pBpQarscXh05pcL2
BYtB6Q2E3JNz0QoMgQoyYWvJ2/ymtYAZ7pH6SCS3F4U7bR58XgLE0pepEndsRvwbR8i+Gga3Vkga
pLNyMvmMk2ZGASyHjVrcW/FEeGo39IyXbNbEV3x1CCyHWN1ifR7EULHNPkFaQEyGygXFYrvT+4vm
UGoRd2GA8W7zlYcSvve62qE+ahKZTumGyZ0qdl+7J+S6O1F8uJQ9Q31H5w3KqoY3gq4KRvbWbonu
lV7GzFm8VAhu6u4nVa3eZV/tdlGqd0MSDxIqs7bFYf2A2TauRIDipmJWTaJX++fnGeP5Z/7K9kio
fmS9EcnYt5Rr6qXsZBUugjJ6zwld6+J3ReuAYUfvUSAS2uNC8/FLGNl9kJa5xLh7JyPRzGx6vpHT
tvWgfLp1HUuIx9E7OXqDF8iQ81UZJjzNHTFwm9kA8cy2+7t5CYwPK20cvtwqkyvGjYIPfggkxXTQ
WllnIRdVnKDA0PC8fxfpJRPhQRHiK7OQq7NI2oQs5h8V1CPuPZLpq3yCmuTAQNlnluhRbLe5RAXD
kSrYrPDPmrZJRrOUFqLPEbzoV78hNliOvVkFvhIe2tCAhEIKh9rIBhot+4FdrOAa4JaJ+xolNhFz
3ygLSganS5fPXh/TMJJ/4DWwvxJb9cV7R3bhMkCZpcex5NtH57FFuNovruehYSN9ciALS29KA9jC
b8ErD0zTdM+NViyT0TCfVE/UBLn+jDBD4PmFWfdVflet1gw4tAaCE0FW7oogGStIL43aYK7ZoghZ
8r8SuoCoaPYwvQ/62KYlLbzUxqY8QQzDoGbM5xaZwnqha8e8pw1v+mMXAykFLrTW1VKUpGTBdszA
mwU28RmUaSMEfJl62TXYJdd1zpg7crAILMpjJBS46ljqrzWF/VmrXwAFO8/nefS1S84xyzzmKh/6
BOSEpPyb6GPbWxZqmnWk3zFKm7/axb089xbxanxdCTSCae6VNiKDGw2rb+zQRB4AMV68gEprOlp+
mxxleuSnO6EpRq1ojgvPPdYZtZUtIwhnb/A3g5HDC0UuwyLeQUE3sYFzqiLiLG8Mxz+Hw+o8ty+x
7GuL/qar5klczsN+ssGwKeEfVUFcMqwkgtLmbG/fAhj5jRUGunAJTzUEvnCozY01iN8meZIhylhW
3PDcRLsSDqop3HT68eKGIHM7X8WIQ+fgEgeVN2owpkN03ylcTTMEbEnF5ue0WLKv+o6bFkXCkvsh
wEF7m710Nj3IqAOkhF9Zv0UQkrBVFAnh912tdTBGyN3DI2L2M5uYhtmYVSuWMakOGSxFeNyE8Tg3
T17e+I1zL+6n9evBjlwTGXFsRaVj2fEFC6CN9TcvIRZ5YYWQH9cOk/xTJVNrq+WqYvckR6cWbmSN
uC3gZHSWUxibPkEBPnG393rnAKxzQoQ64g0zOzCWh7SLkdhr+Y5eRc7s9J9qfFUlYDF7p+d1aP49
0GZBOjqoCCS5lUTnUeRf+aWf58CHPnmg3+Jv4APKYYCSeJWXy2y3XvbUNYtryIIsh9BeFwFx5M+T
fmzn3t8yiFC/hA9qzR7ZJfto8dJ9fc8AgYfF4qtT2T6BEVDTMW8zyCewN6/XQm5sN9fDUGyn6/du
KkLwZ86VeXQWtJd5HukGgzngoWTRzj8h1v/kM75WouVEZ/d2BIxCWW79Z3FFCi832rrGHZgZXO6/
eZE7WPr6h35nBarx0bZk8BKjuUrVj4yZdgDo17+G1HKu+65eGhaFaJp2y7sUZYS7IG3xHKoAHoBA
pg3k93XgCnQlkAtoV0hwbvy6lpqcFe2phhbLnP5F3cSbjXgruQFVWtfbXNpwYhnSF30/IW/9Bt3j
KuNf2emBX56HgTfxnUvLX4V7SEmMBvcqukjGSjyRlSgrSMd0rvxjRDlR84Re+b92gcCJNPCFHzEl
pS/gI1sLCyyTafIFxz6oyaXwXda1QEqRFiquAZNApJ1pPCl2Tcp0qMrkdPGEgdMTtMeGUFjz5SRP
pt4fpkctIuKW3dBwGHGwrvZQZ61nYRdzAfnNnbA1xOOEoxpejGGwDsNNC+wQ44u+9+jhD8piMVYT
e6kDWHjVFiDnx6THP/bGHt3nVG385MwEUKm+Q/DZ5aX4AIJeADL1EHBmcTnCUG5FtQ+BMQosh1Db
7rByYEPABf/LGKzMaIp27JXKEghNQWWrK4JLyh/GJQnMY6vKIyUFml/QzLVd7LkP6wbyIfNpst8R
RXoZ87NQ6YbsMx/N0rxbvKHTRvrhlkmvyjlZAD/m05s1aH1EronX2OakKh2GSKDShcwHcC7s37I6
/a/OHBT1LDNsTJNAvCmBuzpYMHoK4HU4arFjq7ZCzhLQlzke+6dgoNDONE6ow7XemBxiMLIXtPUZ
7YzSVW0HiZPzJwKA1VI348CniLtiSk31xOw85L8Vdg8PBbOvovudcd7m1IvvULVvMBdSY+F4QDee
hR9q5N22HFi545HJrlMFtPSH5jCotPVlHtnWytv9yh3uO1cNNckWJBC9YCGIzkNzf3rPNJP1id9y
riOmMLmMusNhqRGvTOHmrQvMbbhwbhHTEhlhRGrdHDRpESF4QeU2H7XCV8KQWuvyGfdu1xcrg/04
IOJGLW58u5vIF/uONOkUhNmEepFH+zaTQxIP0SCAb1R2gXvq6IkpkuayVleRThUA48wpjY922c62
HusyKZ5HZRxCaepKcVCMLPyxAsmEZsFnfhsoi3GvL6hc7xbAujA66USag8xnTcWp1WYQk2j8IJqy
AzKjUWoVg0W4MMxhzIc4w2ZtwDRo0IBy4hwLDFur7rkSVea1bCAKszdlgo17Ng+W73hC5J1HcSlN
fZoxRqPYXNcULPeRIGz8SjdjtEA4ncemeo85sAqa+M/76EdAD4exGLIVZP0wWgfMiG4FC+c2u001
+BVFeXQlF/rwTRoVTl6nrDdM19XSes4S/UPc3pHLF7xifU5nAFGSzgK1me6mCibcmguq9eJr+VNW
koG95owdOFVqZvoXzT/iq0WxorTl8SnO32P9Vuho7xDagI8Yo/jOcQfGDHe0A/yTjaHYV3lXAxBu
PP0BVxkBSz5vikbCcDuCOvJddHhHmetB0kIMctb2pkxV2dMHuATvm/30uyHPV/A7m6lGMawG9cdH
K/1p88breoqOincIcAn72elpNpAoqs4gmTGUto3AacNA6g5mNrnBpcutSHeggq6QaYp2qu/xRQ1j
aRkLWn/YBexQMYMbt/Ox6tNarWm0+vPD6PgQONTm+am/5xmk2vJsqbeKeRXLoYa2UJGApAPBJk4q
J8iUmr1oWhLwDbkyMbalx46660PJ475GEk3NA4VzqhMbiP1MgO8a4SsIznZnbeZGgyq0/GoQkPPZ
oZK3S8S9YYCBrbYE0BABfQHFBrtDGVaqzQ4Uwzkt25HUVyiw/2uAuXU6paDu1KWK7xtzxFV2PHmZ
8MJUf8wnTS659VsngksAYyv+ZO5lmVGQICfoa8odM88i8Hna7ycaUT2WaJ4x18y/kyn6fyhtJIzn
597ZEDQ9coxky21IF1SV2opXAHZXveEjf1GbOK6KZag/iqvqKeE+IeLcdS61hXGhCBdEZF++7tAJ
oZTYKTzxbkUwST22QCGxOWkY3CejEO2elcO+SmcsoTGCQayA14z7RTKzqX9Vi6CCIp+yCSZQWmLS
z6T13Y3VXbZw4K0vRQoeEJ0Dr7IvFQrK/Qb/LhWu37YzXStuIUwFDM6k7f0FOZ0EMvS51k6/24fQ
PklJQn0g/a/3QYLGoYreHqC+Wrp51VBV6aADc7wuw3HNPSmw2C2b3rRTtB7SYH18jrpcsWjFjgw9
lzzGzW8/5dGrPqf3wMei1PQ2kCUTcEwipBWmO2Jfl1bx+SvHeFdtmEp5VIkcCj6apH/A+1E0Zik9
CgNBuLeM7F4U5Kpnik1UlDC8bQppTRss3DVM2b4VK/RvRMiSF6qwfIExTETB+Mzr1/mE6/vEZZbo
7K1uHaadYjjkph5m7cKQ0KbJAU7Oo0ZZiHHj7EHtE45omlhIrW64MrTuvwXS8fsiM9qrgcPhDrju
m78t2CaCf06GiFfhCbCIOfqiT/hSfu0Eg9vTVno5bdcRzk75oFhfSpXWafaenGoRr4ZsDFnXUvjG
XUcy7eSsb9GZrp4h13/Vt4/9qeRc0SlwJGBRQ0fzUSNxUvmXmqreuBAI40q3iPhtMXPP0Y9RkBlO
f8Ysfk2ej1YjzrBLO7DDwf/kffaAFSywFAfY698XY+HfsIcsg6eE8GAJ593+NpKCRPRuoZ6ZOAXR
RhB8aBWmrifMG14MmcYO43iuJwNPg5H7uKuDzvMr+Sqz60XOkInVbI6PNQpbIwN5xMMgZ404WBVS
tSp0SrMD5Sf3JQFCTOmSKwOL7K1S04rnHSAusadPqtJb31qHm5jZs2R2wP2hZiyU8J6N/r04vlUC
V3pirOm1VbGB6IdODeuukToguLyumgupLPp4LoR+4BPBIMNIGhI2KxInKaezh3IKLcrvGqYsfCde
pADyT8Sb5kzWBY0NT/Yh9PdGLXQaylj5awPzjUazUIigjLNVEP5AGKc4RN3OYRCZGKW38QDEb/F3
r7CBlDet3LpyWx//zS9PFA7u4903TgZFi3DzHkD/LPBPU14w5ASYV/VKlNtXme05h7WSOaInaPFW
s4gySlC0gP39k55sMmWLP+lxrzE7a/OKgsyi3iinunTovufpuO8QwYUbcqggwN/UGe0/TER9x06m
yUuAyMPYnuOMNsnoMHdju8VgTCCtNk0AvG8BeAGeoqLfKH0xCOnTMJqzL3qMdAJdeJqoM0NHVQEp
y8kV74ovcTLaEe6cy2InzTeOD0C55v9xjA07zGkXyAUbq6Ifu5r+uD1MGQgY/ezRrKJjFafNxhzq
FUFTJmb3HHNvNSTZMssH3mVSi/A2I9/iWfqjynX/Yyy00Ecie9c1KkJdQH4J/+q8TMTGDm6HEoML
Lzm/sKVZFVcL0aBnCrdPFKF2H9L6Oscrr3GJONiE5LZcSPkvlllrHurgamZGZBTt/1yYKAg23aCl
Lz8f6WweCuEQMao0gGhARA5FnrzEG8OJbOHy+OUGKXHEwwlwwsrSDpe0eKBbY9cRUsmjNPv4uibH
/ChP8JKqVtcwfL6b7IIPDbGKBiPnNyIyxbBOcDCNDj3EGvuO36KkAHbnaJkLYByaJGBqWjatBFvk
1Y35+JZhK8XVbd90y4JJqvmsLpLlk8GV5l6NMsiEbWb64PqX/oPHAKPJ6+SQ/LoyA04zqDo3pILz
gZjm1K1mKlaW/EHOSITIigMubQxwx+q5sPpti/ygiDYOPKihStS8da5mXAvuTyo9kgzNV3q3b/Qg
/q93UV8lkhTvU/LTbJAoiIuv69ugQ1epaSg5nXIvt1asBawfi7KN78i5w4S1ZlX8J1C+wtsccCNj
T6+DP43Y80Dpx3wXPax+Uuia9bcJFWhMeFZGTZ4qdQ1y/jD04kStij7R0ImPPDE7Laoo5IJbKrdG
zVMEbjqmLcTxKQbmKYQccZyB3oaNMaVqO9DDeqfgA3inqx8ox3cIeT46Jy2PmUOCD7bFw/WKO4a4
2xXwrPoeqrvmahHEaXvn+PmdDmCrBBQNSrFxkHg1M+YJNGkSNFJFEnp4IUd9PYU3+uOKFRW9F1N/
zRnnNl76GIKHtutIb5v/ruGwcbTh0fJpG/YgDyF/AFc6NL7Q8CkACv6LLjHDRsm1vuB5yBSCKQlE
9gxA4BcMlzboTzrzQuOOM4MeScj+SkPDvaQB/a4kHPeaa9JxQJCmjklqRM3CmBWM/7010hRy9kvM
hCdpyp2UeK91ELugRtZrEyQtAVvcjFlL1oaKw9NlvQTkPQiE+Pglo7D2QMVD0/trlOCmIrZg9cAS
w9Ejyk2EjHuNxX5XpAJeFfUQTlxCBD+Hv6uc2g0rGxzpQnSiYRGAktp4ZbfTqim8RtIkM3wFfUKc
AR1fYcg0T8LNngTX1tHt7FfU46TJ7FVjWBtT4WeWBtdhAttPLQ9Rc7maH2kZJm3sGVWyyHRk3xvG
nfuBTI/HYuN9BzNTInyXADtBnl4AiFoLlUoXJ1Jap+bsdlOWSyOVJtuy/wvUQik1A/IHwT+wakYx
Qfeaq4dzfb6BwihR6GY77ceoYmo8hq0YhdY2UU1jBjSxvDwQJH5Z4fhggph1M+jTCfjZkHldquF1
WRjFdauVR7a6eQLxq89UXPLVdhc6zRxO0YG5Vj7Qz9VntqqlmSVTxSd1vlPIXPEp7NJ7JZ1afNYg
VT53xvsCHqD0ObhEz03g2z5GSoZnwELT3zGznbdtyPzY/fTpEB1/xHfNcxtgfawJIJ0IpRpzDlQr
ERlDXxe7VMmhiC1FbNZhHjSagyeoxf/ZgHWry+ZEqw/OqOA65221zBVB22wSjRM5lN152HznOHeM
adKW1wSaNq37se1H7rQx5LzMOOdTy9PXl/Wcs1B7uR3i8QGst8vgqK1soG0B4QkAXerVQIrfsQzS
L7hhQRLl0S2CiaUYQ7ca2Ms1QCrp8BrsRlxpXKaMr1j2VU81Ki6kecBzUpKkFvwyYNjeQkI4YGYI
hkLAOZIwfhh5YmFdMxjk833SPpvlenvaP0u2Bhg+q9wVSsNokhHBLXEqjBIzurMKBhz9EM9pS1CZ
FfzF+iD4v3LUMecbL6p/dGgSBKngsRutx957IPcz9+VTYV42v1Grz0iF43GHbgD3BTWDZAKkkeF7
whDPT/j3NmvaX01n2nBjLiai/JYT9GVDtMeAESsPEXxNeOE3Hbg8kx464f+v9GILPbwKXp0HEt8v
ukifAM2hpgxg3TSLRRgU7M7EMyQuqejU3m7NBTNPLH1pAkkEURzZ4AaMezyqpuxyaKbO+xMAyS3R
m0xgy3xK5PcnsJIhscwrBJqbm9ew9nM3myBfRJTlO9FdRccQv8/hRhHGNQKNyr4tf1ODlAtkGpAB
XH6t2pNgXXyhRXcuzFEsnMTMz4MOdHK2tM9dBijcANHbxL1FYFDE2AJdjI1h/f4HmQ+8+cCdc8X9
DNwQ1Exx3HQSyRPyPTUoFz4cbbIN696zjvlHXGPD39CVkUNUb0nsF5+RLy1BFOlAbmvlSiaOD6uI
3HFv9D/jAI32IOFYWZ41li9Aklyo4Ac3tPB/OK6Owfbdm3xAaDdsObIkMBRBRZV50+CSVZPPDnBg
PozxEnHtMf97GTaz8+O2YKmUpd829TCw/tKWYDw5B+knWlpCMlVvVbYb1qYgLCgaahb4JbFr82HD
m7vwhZjyKbyLd6IOcohd6+m4oGdqJCcQgaytpHAia6OePPtKfLCmsFyI4ngf7J264OkSjAHx4uII
Br0/NfTv+5KJemYpMc76S1BD7pnWGI3r+QyT4oP/z3tdMZe3EvCWApqTqCqJDGPykTtYLw+wEUJu
O+5Sm0IC4IFXeefRKBd1NeH4vp58VcwzV8iLPCRJjGAQ3dJGTi88tTcXuod+dE57P3ynwJXGelai
Uk3JYr4tWMgSXKmbj7k831lxM47hd5PLTYkJ34cL7eOhxrrgZmSt8nK41T3Y9chwC9t1S84OyLWg
rY+V5ert88e0bf7H+cTkBcu8VRo+H5p14cE/GbI95XjnUL9rYjnRlwXFUofms8ZiKrbVnDVjJchW
HNERQxBQ+krfpW+YVq0eLf8SVN56TfNt/3KzDdsxNADr+wFmreqFeTe8dpwWU8PoRiVNbS7wyLpp
G3+NaEx115ys5Ickx0baxYjrQnilD3x4ENLgD+AY5iaEpiAfMo4e99fGY2iJEN8fd07UvwvLr7+1
H6LyYtcsV2H57Lh2lZnyX0xcAHVsOryvui9nfj8i14j1PUqVrZq9wUjBLJl7IVH9Gc2+snXBJ6lC
z3G1cVrPuCaIiF7GH3qSSx+EtUkCfQ1UJjtGPbwn+Rosgl3gZh3NEdxfZOAYAZ0WX3pMjq5S38rG
E9A/CtRyxbG+tfstCcZ57f74rm7VmvNsBY+QicVUBY6un/pV//MnM0MKS9njYA8/d/9IK7VbDEqb
xmAVrPqt/HheI76HjH3FJboHlKb8GQOib0AWpk3wYiPL/SyLBUOijVfJxRBeGOArrCpPrnH7CQU/
ICTKBfzi1X6CKzhthIYOZHK9j80Z9CWb7ftl6QsgUk4wE89b14M5E+ZuniVMy+2s9ZmW55vN1FF5
zMFs4Jl63Gx77qv/0ce89lYHN1Nv31QKF/7gIkI8lJk65KdMb5F22AiZfXJK2miUumgGnFVhDz+X
00Twk3ZbY+/76AHTHWFyU4rUM9TIB/YudgAdWY+k/upyulesmQq+HcKwVMHb23UN+ixEdnY1bs1q
J2Mr2Qix95bLop+ZOvCXKFyHjvYsxEFt2asQzVNl44WpxVaBmesH0oi7R7sIZfdu0m4A9YSU9+C4
slXpH9nUPo3HS/62d+rk0lBaANBZg8jfvXUJVS5JmJgMdkRcYRhiFZizqcKPqK5xmIkaIMkYjG7w
AJHmC4ew35JNqtiaiSpnEsmsgY+IqHth3ZgDYxizU2iKIX7mU8jWV+f9zG5DOXldygGKaMFmnRra
puU2w6iD+cw16WhjcQtY450JBnpymmuUn6jsbZ5afbTKVY03owedQngDbTMynH7dkx0jKHjyvrVJ
JwI+ToTUbCOOnHc2SS11uUhGRP3qC1Y0nOjww49dOoml+/p8mXtEW9xYHtDjt/eYvlJg1W9AB5Pa
ZZPx39dI9ELzMJb2XfvviEoQF8l/5Fd1WP5L95Cgw1heDKAQatrK7DC+o7uh7Z88sUTXNSDlMf9c
Je4K+e6DItP8/yxIwyqj2ISCZA4N4mIM4g5kinloSage4oTG9jaWls8i5LuhFEPnq7lonPojsDH0
xIgwhn3/lxZvhQz2TWNcYMSujtmPalwhvRhzRj2RyQbOADpNPQ1tWioio1KW+xgYlJhjXKQRG3lj
x+n7WX/7FUmAYI4bdEMUuOkVdQm7TLpLw9wL1iFKwV0FQfW3HBALHoh3xoHj0XtmZqlRoFZ7e55h
Dy1uSubdX4QatMX3AMcoRqeEfrEI5yTA31iBWQujPPeflsPPha2Zy9wIES/gr+fuPimo/QkF9rZP
wPvuN+dJSP7fl6CqyJzMPNgf5I6v6kc6KsjWJlvjrhCMGTrSLBskX7mUTiiqS7l2vNX6MmG6f+h6
QeGYf5AzPnFSFwRcS0WrHdt/PoGczeLNwVAwLIgROqj40RbXR0vL4Wl6qGoLJL10PQx7DIULZjzO
5O/g6KT2mwbdvNWRPh38oJuMspSiEkVu9o2+4b6Q4MQ5mhMGxJ5nH/5YsxiznQuPlw6mo9qMgmJr
JB9Dk8hViI1UGapnvYO19V2sb2cDDYTAEYGwQ1G5qZbEKXKKXwQzPqEuTq5i6ePpJyySfHatKHn+
I0CXahTcNOGdjuwwe4pHcEOh4F+GYJ1+ko4F+yZZGGaUHGaBt0tfbz8AFadvql5qEnb+hxfDKqCM
qZTFif4vESWAaI7eLr+CSodJ5SbvLaKVT2v10PB1hTgU6OYs0WecySKru4kJ6gx3/sWDXEps0DBv
u6T/DnGf/7YlJ90MZUUIrBm2U9bBcOV4Yr5GFmy/rWFuQUctaNnG+g3bJ5q+BIursB2sY3VTUNOv
wMOYE5pvzVEdBuwdsqItHEuLNvK+vt0EP0MeAedSXV61R1Vm/zDz0xUkp8F1iOgiqGWdSTC890sx
rJ64DtB7yDj38nSiasC9UfiLtBN7W29MsB3l7aufxZOPkQ9yJ23b6+IlzAd3NcJQSrZ/tYH+a/CH
vPxjnlR721+rG6SWOhMap6nKind0etjiQHzMld7klIRS7pnYMvIgU3eGKJycm79LD0HtzkN2XwNk
xgKaLqZ9KKQqH5WRqLgzqvLN1kCZplLsr9YQXkV3QgciMhyzkvS7f7Mye33+yyTLOl9u8zUH1cxK
+9agG/+bW14/aw7aDHDYPZXLZI1okSyZx+n2J60S6XAc5ZPYJQGYHBMur3RrJyJ2NANzU0fqJT8P
cUzA5tXd9Jt9J2WA86shnGaFG/i99X3xf72o831AHW1fb/b3x9uQxhGb8U0Lr7gCAj/WdO08vodP
OHFn91kF1qJjsxjAs7Zzv4Ii1mPOX+j5Yrk1xHjz8FDMArxzvlRh9E1aIpdUafRZLXYtbKiC+JeZ
rTLiT2OKewwOfi34OuITmk6+UwMAshJ4CdUNYzbw+xpr8jMup4kahGCAwzM4OHOf7Bm2tTCtNC31
5Y3iIvq6vKVJISuRdc+FI90UcJv9Y4MwesYvHzwDNfwNEIe/CoZuASHsynabiNqIVeJGcaK578j7
ATjTaTF4FRdq8zmDKBJ0yrOcpv/0zSTtPzYJqCJAiInZkIq+S0FmrV8aY34/myWjppobIT8Za6aO
5RVvgFQrA06SmmGYuodIlVcRGAeKzBZnQTxVWrMh6ARwwWHIvF0JugHglk7K8fj7QPwO5ZwYSd0o
eLNo6xI6+BOPSHBinrEHvG0XzmvBcWwiMuSgbup8dXyK7OJa9Wckh+avzGE2vxE5+HEUYeaDc7uT
IA6fkW5MBQa5MXJSyYCNq7TWyj9vkYaB8NM2Ig4F3cw+6c81V2iRjhPaO8YPpG1bE+uwtmMyE7Gs
TicJj8fdcqJ+Aolgv/uojDJLWBusNq4inJfX+gLdBePyjv+KlFJ6SKf45jljPlBBnspYritwsywy
S9ZhlfzC8leK4g57kQb9WbMW/OvEx0Ux6X1y69ebpuzBJe1tEMSe1Md8QSZz4SrI6eOQpC4osfuv
3gHPEoMYEktMh1rojHpPwJNM1N8DQKjDf31bq7R3p/OMgLq40pg6SEvqs2ReUIE7CrbKJRjDroM0
gEzYEagXWWTjONqEFhZqFlb8Il8YuWb/8PEnpfbkyyzqEeAf472UjE4dp00V+Zkwf6GPhnrr5+4C
deq0t4/2gUBOwxhLvAhDoKpQN2tUEo3kHRgTBioysmwCK1cz9sN2nX8aRGtsgif9YqLQNvPCsl1/
T/x6va16HgUjKEk0kOEL+507ThusUu0VdP1PtVVPNDvFpPGx7T0U4NBuKyJRmGprZLyx7Z4T1vnz
ECdYilYAwokG7/0nZZKeZOcZdgrDCuPZAZkeUMeI4VEGCtaNGviZMA0SHQJ5guuEUMewGf3R0YWJ
1egyzH3YQDvlM1hKFAmizYp+m5B9qaTbhA5An6zVll9k36fTgVYvokrGPsuXy3KUSi8iuBbGTK3P
jw1HPNXASRj6HekQN5f0vCGIPT/+KdOkJ9PEs3nk7I+X1niNgFGLWmcmBL2uUU25TCU8I6NYDgc1
RQr+O/tQAwlhHLTtS4LyEf7YuGinP1PucE4j9C2B9V3+GHIsD/Fayxrdrif1kjw7zaFIv4HE2qv5
wJceBiUA4w64m97iNxZ8MVYp5njjXC1god3lY2ReLndBg96XSwPTw3j90UKEftrCOFCPdlBUTXat
Fyr3BcA+ljO6zkeAE1fqtBj51ieaiPdm0S8x0RqQsIwsRpM1GavNOFHn+xksmf6nvHNNFBxkOvaJ
PrJSM5r0akyQpywTZIqwNtBPY8BTu+cI2Jy9I4+J6LHvO4hdtXwpJxZgxL9OqYhaaIckx/B5pkrS
5gb6nJE5VAEXVILtJyfI6cn6Nwfl+JCR5D1Tx+cOpYV12wK2AcoMBU/zGWbOw+JWBF+RZ5NJD4tn
7mRLZ3Fo8OXfBsOULpZnL1Lr4OvpVMkzNtstcg3Tjn+8DO+KvBCwj9KRSzsyzPT6BcTkiCy11LJd
GwXyLvNe8W4m3CqsxFM4GbbHUV7I7xifg1qRZuUpnblMVnUWadC3oW+nEgUCoe4XzczFKDxCwqPX
w0WlGGKuWIma0MSoi/HfWSkfiySGNCVP1BBGTW5hyKtM6Lxws1AkHYX0lT+YaBHYYzDHymShIpx0
9Q8ZwCibksUQSjswRp5HP9Ga3Qxytv2lEY4T1IhLgPF3ifgQJjL480xUQTxgMb2HlqVfLpJEYEbo
vkbiQOZsx6PvYkuWrV7FRrHD58j9u3xWlBJ/MTcvOxDN7yX/5Q6Es4ereQrJL+STXBORuFZqu4hW
YwAuVTTvOz7VgFd/m8HqYW4ik3tlCpmoIWp4NpBPltj+4gnGScZikrpxaPG0PlTPR8Pe+pfs5gbt
j5is54SqfPq5uCmVizVG3arFmK9k84qXhWuzu/1uJcF9sU68idSQu8oMdyCUKAiMHaXRNy6Qioz+
VO0K1bWoeqy5uojkKr2GGG1HOOlX+X4XxYd50li8kOHXnadOW79mD35z6tcVGlZyO3RWPT4YWURM
dZ8cMggSUa5XBZnYtL3TPyxw1UwVvez/xS6r1//SY5TYMuqlIMhPWQUOqyO0i04zFyLAgsLaq+7z
N/r2faSECOzksxz/35YnMcRyx6b4lU5GXIMCPbsrvbW0PnXxyXpdDBbnj4XNIRdk2iRa29011zlo
4YjxOo3OuO0hyzd3JkLekQQFVf074qbEtj1AltJnGXBT1VSupuCJr24uDmAcseXr2IUnEsQ8myLu
S9NnI+yt8loiHwhI0t3BLZzhMeZkBL32vYJprUyWT/WSuZDDzJxcA+jQ1FReQOcLlHleno3D9vaD
CQVCqNEbETZ5dXvyrf32DWnOpq2dpikLjW4X0ehm+I/ZeE5RmC2FAAHe/M7GYNIwhi55nSWHDbly
dvBvSvAHB+xNRMUGzVCjTPVNbM4J5qD5zSH7whbe1ChGtrv/qA455qNkDxCUfy/jCeOttJQIUJCT
WMZ1CWZ132mkKnRcUAAC6HdzIrkJAWJa1XYrGamc9lYD+Hy2qTyPFORl8jgbTYV2oC5xcvCbnxi3
GGih2HL0tXmIwC/Psy5uIY2Y0FNxAgtAyhgfJUWkXVexgB3kaOXdsRGw9HZI0Qp15k0o/yeXiia9
J31nBIf4b1En2LcZLaLjPmCHyUwq1EVwE7h41MsSMMdFbCl6MQaHvtDeFThlSbCIVrwELUaX+cLO
xvYn0ebakjslf0XmlaBCpNIKh4vcs7xSBuWOAq8XCG0hfIS8+4ixNY5o9AFsttOXgoxIncHFT4n8
9j5Wu2tn34T8hSsWV1pVS3koH6zskOp541xvJ/jwFDNX/5KUoDarzBtio3tXtoojE256m0lgNL2C
bCR3n+G/wu/ijWKm0/FFKc+iYXH3Kf9kXcDt7hqLb+fiEWjDa4BKmScumI/uzTYleWtNWdky2r0F
uBcMrbC2AxgqWVOv/O44DzjCubM2Kb63q7mcpN1+v4LoR7b+hTFaCclKgUWBkYrKs/zLkpdowNUI
5hMyUr88mpI/zOKy11j8je91hPqgPuVrIpAlG5kvYFwd00ljMcUJk0PaPJDFR/cGJhsiLA15GDnc
vulVH4CoI62TVBCraNXCGYBI0lApzbT0bU18dMHDGI4LEhlIEI/WIOpXcOtVZdLiAFNCOFMTf+5y
pMPxE5+zOGcvCGLHIVImicjnIz1u16hz6zNftxc5hvXpu106BuiMAOX9Qp4p1uing+2euLgV6wun
rw1y42P0o4QMLyI8YU40U8t3rWsrBBt+wEBPr+Aow5vs4cC8dikQ0hy6ZzsPFvFLXqu+2FyRQ9NG
AJOrICa8/uotDesud7u7Xp412DSyCC+/OzfG8F2ckWheV/w5rMbPvFjOuidMxkokSMSQSq4oEtL5
h8D0qKxD3kHg6EUlw+sKJZRvINKpImqc5kvDqxEFxdzKILz8LW1m0Y3mm/fkeC2aHrRbfOrLNdkw
BlsEAUNbg29N2ZDWc5pszzs7NLG631MllyCV9RSdD5eVxbgM8tGXyP+riORx31BUm05jrtPphmrB
AulHYmczHI1j5/6nOqv1kzoTXo8pHU+PUf9bQL59UHiLxOtKPvVDATeegFGe9PcOw5ce5OXFK4av
x0hiB9wCT8WqlsPfDIAwLboFHDiEAmN9RsiMrDezo9qYC7vknnIf7rFSlfkTrLhJW4T4/99dERQ4
IjmOBdpc5VdKjMSJMS2Ev10K3mf8R6PrLGaG68f/Q8Lp5140FKMcgQyP4Sw0eIjXqfqaRVHmisOH
8AOf1kphUMkrH+Vp9X7+txFgF/C+kebvRhOUhDXDAcgyF0WbfV0sdKgyEV2dUKhJBa7qvbDAzrTN
9mVK4nB/7eN8h+zhC4gVz8DjZQysDqjUdfKqqW3s6PQioRlrGgD8IxGONymoTEBJN0gbIU3+kVqg
//P4E6PhDGW9t3VNnsr+OA8MV3XOQNdobsxT6IU/VmPHb0MbCTAHLTnLR1ns9KCqWoww4a0jwPKw
QYPSrizwtYZdvxSX+AVONyf6nkdDO9Zry6nLS+YKqeaCHA5WIK9HZEEjr4zgGn690mrNAZn/zbk9
sYK/70pI/UTXv5/XGdSnnTc27iMLiYO9zjpzXUgJXGbqARJPPi0+BqE4/l/zPnNGwYjbUMHUjcXN
tfJRPn2PBkqIJR4W7eK8CywqOWrUWjUZgRVUyVZrQUyXwsxaubH1oklgYUekjRvobZS70hXZiXpR
+W+u+mjiOXJbJun8m5r5ZEpN0n+LYteiX/s6RQC6IRDQ0TgzDJAFSOY+8i9kpAyuVPG1D5WgqgXC
vWIfWsFohK8aPogeKd4yCk/kg9uiXq9pIdM6rrLmkm+DyIDwcZT8HUMqPaZ80bYOny1aOaVNrB6T
Z8qRy8yfvV8y9thMLvr9Qxd8sIKF6UkUj7BpIT46LaGgL5BSc0PWiJ8ZNlCE51OQ4dR/C0yY9JZe
/V32LwMJCV1E3l5DpTO6hU4AaYsW8SM1ierD6BEqJAwFDhUTP2FtR6/GOAIR6vKTrdiPg31Ns4tY
pOAZBKG011mUW7w7/XPVwZ9nOyWHdGapdKBVCHd/mbDOzhQ4yk7O3Ui10+fUkkNX+tYyDsK4inrO
YYFkCwMYwozTBHot0xOYJdddBG+T+p8+HYC8Iz5D3K7mq9blat3A+P/ID7bqsWdpjJ7gu/ArQog1
+aplE1bz7kKFnciYBrJflmVLr4srXukxEsoPtFzif81jNYNR8MfDVi/WDntWclbyjJ+bzgKLa5Te
WPSRoxufs3xY7zBfw4YlsNMFtm57QAq9Vp+Ptvrlq8vEBOKHXZTXG+quoHDLGVV6mW4S3KiBm0BO
EOnDr+L5+8MJPqSGhpy8aIvwnJxDJA5AznZzaHrt151QPAHp6e1ibf0ocylQLzfiYIxAK2Z6nhPu
Q/9bOnx1snT/Pr29d6Lwyq6oPAZA/57wox6mTw9g+IyMNh/qms+dVx6ELAO0Cte3QxReMrQHkGhF
VPcXEWne4rACq86U4vCxeQ2Jko8AlEl9j75qKqxN8PycZFpK6c1XCp2F5S/+WrqDjuksyw9CVye7
4Y9fAV17xNf040n2dXRtt3ZH603bWc3xx/SZl6wb4u/eyA9FMhPE3YcYNsTYsgJQxYzKE3Pw5sh7
3T9wDx//qEKkPMYzWNURV1ilyWQBLCIQC3kJVc0x65k9UOYbrLhhHN3zHmul3tUAV/vzmwX2hC96
/AjWnjw167e3uRrWV+0b75/ku4nt/jkwgf1XnP2rwbgJ5yU8Au1E0uzDEM3Gu1dqAzzEb+sGz3F1
7o8RyG8XTQ/+6p3mfT9BuLHbjoyGnpyE7ouYt40xUePZBhXTPNcjzbpm7cocOPNDMt7Kb5sL6wBt
EDpUEN0ICw51alXH9ddbrmKceXF7awljBNqeQfyoeZrYj+r2G6rme5Lp2ZPluZP9QtX5SpolqHyr
kjpkjKwDOkfHL9PJ/MtDLTcHRNysXFUbxC/mny10rL353/4dIxRhuR3RsplMBejL+oSevEsegfyG
FvdlD2bwNEFKw+P37e3eXwXxvlzS0mDGttLK/Iki65DfMaxlnoXQdFpVyYc5R2QZcY4DKWXEp27n
kFrqW23/04LOF6xUdEtdP9fxsUspKiTsbbYxW3Sw85HdzKcc1UhJYYeoYTonZ5qyC1jYyvpFneKA
vqyb4HSpXnGuBHUbUXAVU6bf0PsXzziQDVgmO3pLr2lXNv7kmq4YbPKHKrSqXEa/y2Ww9t2R3crN
kp+KZ37sCPb0q1GbNHSRTZe4E5YJj5TDRYG9QWz85Lbr44U4C4jZlQygMlI2WYoOKEOIAgtCr0Ci
M+9EZwJUudP6DedxXKy6ExxjkuXFUgUbpyguJvgevJKpe7Ga2s1RjUUVl5ZSdJRbtghDzChR0DXf
N93WudkEMZzac2j6THjfsctS/EztCP/HeQpN6FYBMtrdaMi7Ki6mhy3LXqGckcd+6d6AYr2hIfJJ
G5U55raG+wykCF6qJEp4c5s04o8Uw5tyoUJSrdahlrdrMe3iBx1mIK1u4urJSwWhgAZ7aLvvIuyR
64I/qeOdvVetdbJlFCZ2Y67svOyICkHRkUjNSp8ER+zvb7ixYFrEXO1oW49VqD6GO6D5UTSPrrEx
f/a5LrtxVhJcN3uB8iOzOizcrqPiymtluwP/e5ztx4n2Tc1ZEStw+rjN22EPLzf/ks3M9v/S7CWM
F9HRJdMQonQSg0rzt1hGa9oGDy4U1ePBVyf2fIuboDBktUFQ/2dwQyjVHZiwiIkuP1Fw3EUJscan
dlWN/kGG4h7ximC3tJHrp7UqHeHSpM9jcEwl3NCdIEJyDEmYEJFT2EXX9RrTAoEV3qlW3rhXv4Ej
8p2AA84kX42ElP/t0nCXl0Hepk5fzHqGNr8EUKWCDm0FMswP7N+EseM16Zfo5fgF5yxD4f4kwv4y
vNJjkNK3PeuLuKg13D9LmqLB/uaRmeqKEqO3TJvBQjBU8szmpxijhHgYuoTkuvmzwnIOUo0B+1d/
lKU5IN2kif007pCi8g+zlt8xOfsZVSGU70pOAwKFJglxd+DWa/6IvVqvn4f9NwxOhMN4f8NIU3VJ
Opsbwu0+JLOHj+SgDliaPAlAKegiS1VDs0J80uvgvldvCqvxwyDH9FKM1rOAH4lpwojsnnO2TC8n
Ko635VjCIZZdjfhJF0Y7bBRhLPcIwgmOFfLiqyMDG0eRLW1X2VXohWnvMsLMyjVr5J2hPwX++ifN
jHGdRHtvsHlFAYco/uFAepq7s8BK9897xmdhs0I3jKWwj5iYB0PL4aO4pwYEf+6jyLtPyOsHo4pJ
3PDlDaq5N4lF4k3Ci941rpFSwkt/OSRljIj8j0CDZZ1dELGZl+xfatxyPlxYs8DhRmL12Sclrh6O
2v7gPR3JNtwC+/YFEklUZe/epRIHMk7Cy9NLAilaz9FpWJai7r4xAY7cDZCINN2dSfXlfVDDuXKn
05eyIIQTs7EZ2uYSbVbqwVnvPYfPLuAcZ//b0MWitfrJKAwRHng+EbG7egU5XbH1FWG9RXI8jApl
0qYxD4Z+kdEo8McEYH9ojG2uS3W8y6zlA32cuHAbFGWBMpng3V0ZwtJVp0Wto1ChvHiCcbW+fovi
ghGY+n91Jw2/JwrrDAYKMLrvFUM/73B84gr0B05AG98E/dl6Y4IHu8EwNfV3KD4vw6jEjSp+mZQG
g5pZ8n/+MjUwiMd/hmkham807pXGrr88ONa9BUFC3l99vkGHaNvDGoLrLzqMyJtDo7x7e3Bq6YKU
zZ1Wup8IPSR2W4dHwJS8EEzzp0UXUpHHPRXUPtTgNll1oQHPxiueM06gzOmAm+eSVfTiRWpRV72G
tiocJtvtebjSFYIEkpFCS4vbDl1WiugGmPZXbkh/Y9OWbkBDjnEf+A9XJCO1JvDbfopjInoPGqoG
iInRttn7BTM6KhykgmTsz42UwNOWl0BTe+N3cRUTYUho+/ApJRkpfczHc7y/qk2lc79hcPtxTw5R
ZRYjNaT7NcgkfV8mh0vOtKFg88HILTOe82Hv2CF+UfSixGUK8rpHEOVfFzAzk5D+axNhBZlUOMly
CxZehvrFLXcctdGNFtusBf6YG0wvEz6OGGAk/1of3YOYtjB/tzOG0tP2qo/PXi7hUF4fdZdA2I/B
84MYsp4F9faINXjiP6I+AdYvQKZeYCHIKDMHLN1KQBJl/YXnrMKES4Ena2MJilDhndbhdSB5kIv6
rMmpYPHjDNp29ICw6T9DZr/wrzDcQ9IL6Sgf1qPBr7Yxjy6O2qxkWZuJjOTQw1hFmdPS4oamx4pE
5yIOzEQq5yrb6ouLOzWwxyYtEkKJswdPJL39ALQL8Ib5QfwQixbjY3kLZiN13SxrPs775W4ZgTGN
QJoNwssMVPRaq6rfS0RoYG1NE1HnubxmIOo83YKsUTIbvyYNSaZSx9gV3VECyVxQEKzJ9PZdCxHT
2ndtKU7toDmFjA0pHRdTXJYcn5ie6wwU3v31DA46zZ39Bjlwhl1+G4NLPdaxWaSOXHNTwSOEff2o
r5vFpfEEyoekHbdwYArXcZw/AolQUd4OhoDT4HJqMThtKOzzjQFGM25YOap2Xa91OpGScQEbjDDW
KsWpE1W67u5WBfnHizQoUzQZqRSKweOLwvZowVnUA4xzdX0Dq6wfyU8TMj3zWg/AmOdn4juTB0Db
OHNdPmQFuEOIGbDDAmjA1AasBkgOjhSVY5cvrOIm5XT2Q+pr5wlMqu2wvN7FbZzS2JYsABI4obGq
yHQ9A1RWBwf53FfTEbWrktF36racMH4qkVAOloSeUQw8JUn6WtCXg2d5CYbaS4V9dwix+xb6lAjD
0iliakPwFYW0TFuzEeZh0cBzsc61KU4tAu1ILaOYmEVAVviwAqdN2xxXJC4359uqG8S7XmnPS9ws
2gOl0qdqNuBpKS4qc9/acjEaFCCV38U5Sv/6fcVw1x35MbFovLUT/jzMHY1R07GzQximqMdSJ6RW
7v9BD0uEtIbIxZ2wh9qSkL1vvi4QlMvhsxIagrrtomDS4t52FCkdVxgEQRKSVqDQsWL1Xqeiaa3D
1y8ZKPbhSpmbf6NxE9ZxayxsDkBKQVpeOlB2jb2LjALiuol3zZkjV1lCagv3MWEU5GGLy/cnZzFG
J7p2KKzemrjN3BIBx006L+QjZLSmN4tmAahvmvb73TJX2XXKdYEonruiy2kmIbIXJJxUrpWQc3Ak
NwYNcqcSBxPnW9oqxoAYhvGPjs092rGFDD/sSb0iilRLla4UXTXT9GO/8lJCx9MCXQp5Qe/PgH/q
AzIHdC8mPxjPRb6njo+5xDxnQNThBXPDirqbwj1oGxde9ef8HIj8T8xtGEw8uHLsoIBzCpH2F+kA
QG3A+uaWpElAt/xvrwJxvUoHMmAL/KKbux1C4AUKAiOWLvytYjUxw/qmbrcpJt58sfYwE1yHXCx2
YyPBKM6W1Sl36TWWhrJ6ml3hiU56/czblIGSSz7RmeaXU/ZQ9wa2oVY0thqosN7top3MZqNYAldH
fLtpB2zR3S6qk/BOp9VlzZrqFKG/JKo4e8XI/TC6zpBQxRSyU1r2M1f3yErwBDJ/Co5IVLiGY1+0
Od1Syj3cG414gH69enabnV07mQBUdK+Nj/6/fL4k2gMdTi8nYlrMmo6XsYfqlqNIbYj9jKXj8xyE
vCDhRTIG+J3fCQH6hUqX/sam3C+bkreGrTMjSpQOTHtPtTE8E085ExhC4AA8LzyCB0vzY1ozbnPv
wHRtiJYiuZIec8nhEi6Az2VzN4MQBQVMT8GvSBSxAw96VSjDQArCiO9FW+peF0/Sb1NjHVxhk4W6
gj9ohWJPboYKkABChSbayAZFP56PY5tIyodbD3yrcXaAqn/EqNaxOoDzfFpAmfA2/n3aAVLlxo2y
J+ysruptjtzfukBRqpvgxRWdC6IStn4CbAOLIm1Aw/nR2NhQ8P10IskuEh9h1nazARnnTViiFhcx
GPUAJA4pfCkYS2evVV1J2UwqVUUgFu3V5mcdiADbR5s0ZaNcbvvhprxUBXFPTTHcXfl3pfAJL1pG
1bFhHOFByibO8b1LF4B5yrIDkgCOvOlILQVPfli7u2w4LSjE8GEF4QtCu8DxvBIoULN43llusF5b
+m8SRaXTQ5oB7tOWkAus8QpKwISFPBcvb8yAXdqCvuAL7vKvKKcUAuMXR1xJFy7bv35BpOCmJ+oz
HLEpv/M8KzWeruxOhRrq769OMzFwJxxd7+AQGdU5y0VXqS4dWNJbkY5guNS8oj6jgGd9Gue7LtsJ
fMoR2XhZBBhsAwUvNd86ipBkaAFiUXP/sIRHGxMqFDWJ7ZefvE0dAy7uODOq2oj7J7WIlnRTOVYQ
mik385KODxKFPAmietbiwuaqpmju0j4hYUhW7DJiW4Rz+0HjDXVFshl+ZZKVg/cJ6c/Z/RwE3yZ3
2kx26nS8c1D2+KWuPBq0dyr4OAf7vNzF0nF+FmMa6UdiV0fUEaLaUSVrJhMrxsqmow73RW2gnO5f
Ri/+XFlhBoeyMh1fSUEZVpqw6pTEoVoDQML7tLjGnOGikxQ5sB27HjSX11vWO5pf9nEs7MlwFG3E
VVffP+1+UOnVFqEHQq3tAnhlQEi0bYCbhzjlGZY8uw1lSeD7mPqNjDTe/Ux86pj24gH8T8ncbiud
DQ9xsPFBplV/5y1opgoN3sxRG/rR6sFfl7we534LYEk43k+nPUKDRBiiM6gRAu8cdM+38qH8HOZn
WL3XTEpu0GsnP+yiGgg81ogqzWE9LtwFPZ2iBtOYNhhSBwIMGsOGeqE2xDdJxdQyNL78W/Vdy1SV
W/SSS06ozZjLcksuYs0KibKYCBKtr8ZHwB8cCwagPsI1E4VAJWcyWwnUx6rs9rOHxm/OcGHhb0Ax
dltc0wty5JT2vYXgwKdjfwzkWRdc5DPnvD+kTqoZrpH0vlnohvbUVTsBtYRzwRDPOQk14kSuArtd
+FoJsazn85KHaNMJa/vfYznKT929GtTwqnYnVBDYeNAFTbeCV141WU7f+9pu7oqSA4KoZ6pcHgUt
plc1dY5eUXOYWAgdp13VoDROOEPiDKmTVkBnFEW9fUeYY4Ws8UMdk9G4FPEUgqk5lrMxqJCxLwwE
k3UC0m7WvNTmxk1UuPsRozOF93dRNnYwTGdkJAYnP5pX3GPFC1kNdd0/LOCLVqF9bY9gH9V8XyvZ
gm0/0kI6yszzcmfH8gmBrABEk+nSDctPkllkv0w6fD2HzoZqIDK0j1ukIvGEtex/IdTyfiKBgPNN
eTlFQs5FRun4/dbiHIT0HAw5gKCAVXRfAGj3AwbYEO6ZSOUFKt8nVl1dJq0GRypyD6GoTHkOmor/
emC0iFUZSb66d6BK7NmdLBI8afjqalWXSAfxgI9ELZfHqEtyVrC+ol50qVBqcfZv7ArCbDOZUUjj
gAmdSl2A2eeKOuxPSkd2zaD2BJJcyk6BrtpUqtHfqZeC+3vP1A3ybl+j9fyJLc8Uf4imGvkbmURV
3Yz4P1hxdvD/BegTPzPc4lECL4fYiKmdpUPxIAoiKxV1MIuYEBgunn67bFFbRFynU/VIjDb6GWbj
gIBhiBuFZQePvAJ6lnlH0e41NMVV1kKj7orJ0LuNGvmNu49/A+4a5roPDQjPzciHwKjt7PF+ekiZ
b2EoAgk0EqgtgUzdGPF+Eam79UumNtazZeHSlh99qKpC/iSNSLyJnEfR0rESFht3qbOgTDE/ZzcU
q0zfEtqqDDI6d0xrGBSs5sRkdADZy6YHYipJK2laZAE+/UBG5iKBrRii0A9DqDUeFZdDhkWynMvp
yqbN9mBIyxr6hP1qAO3g1Qz3+fqAbg0uZTLC9QlWRLyijQvPN2XSQJSaiD8xx7Ok5JrOr992g1wp
5fR8OMvNn+5LcU3C7X8fKWkjjkkxLH4hhkhIKJSW3W4uw3O2zWjcubxmreie1Nlj5K5nh3o7+06d
6hSlS0c6EBYGBivahBDfaTZt2Ma41C6RZsrvpg9q2oakR5YutXaDLu2eTpR/ArUIp+OLgFdEuJCm
8969uABjdyvMug3uZ1YpVLOZyO1heNbIxK9cPegPxeGSgmCgdrJ9JyjZeLLZVjz5rHicPPPcKuiP
WLHc/LVpR4TYhJbNSgf4lhF93XybRsyr5WZ+fNR9NdcTv6af5ExXy+VG1l4k1LcPpCkAG6Sb9rVB
MLDNhmCw9EMJM5dynZuWBuazpEzWa8FZwgqtL9Q9k1eAyIXKHvapN5p+FBzze7+E86NghtkVzD5+
xCTMRuS8hwe25rPQdxeXdOuIj4QZMrzE/aYkQRst5GV6f1eOT7YKbjjuOaKdYEnZQo3UXg5/rJym
fpmokaSV8vHXm9q9H1jf/hpY06eZQ8w/yG8U6ztjnBlAFOZHLVEJZDeeGkgUPna5v/CUKyS24eeF
lS4AOOHgRUp8e1Z0K/fYFOBkZrjRLVyhMEZR+AYYWB+AcBCY/az3nsBPW8BDTTftPOhLyzSj22ZH
fLpbQ6nQktUTu1l+VNsHrywZJupR64MhqEp9Ar3ayRH8knsvrVLZOB/EzFYiASNL9El981oCJ3qN
yfv0fC/VOERM3lwhPIpUls+rn4wyBa0OIavnGTXK2a4RojxJEA/nSIW1JFxlxChuvNYFlqVBIhkE
JZ6tpCaxg5BnWDRW3V2dLTzbxv0S+onEhIficSkvHQXC4sf2uWJD9yXJEWrNIXtp5FOHe7bp3ede
VtRf8ajDrpJB9RVxi+MQHgpj2an9PGPVvNe8oCivck+wbUulYRVZVPR9hdFEIBnMWQWwxGk2eeyc
FvwosYBbZefu6511ThrLlsGJdvSgeG0SsDbMLddTwVqVYbZoBd6qYZsku9Py1EZip0qGuZmZvrI2
BcaRud8riMdjhlvfkfQ1LgBMp8ZphGM2bFpnuRIO5+FI42AZh3vhyx2FcQmNE+xn7xaga1zAMFvW
C52XG1Z7cUkTfHlAW1efn+wppf3X5yihZtYnjZ0KsfuC6U8dlWRUXQK9D8fiqiXHu/KgV0g+yh8e
vABwPMCFmcN/iP4lCW190xa9oIHNNAof35RwKGZtXr1pa7TUKTKAfy6YKNryycY8b/nJfMQVOYLq
SyD6uZmS/HRfVP7+E+7CDr5Ia0ReuQivOiSTBgVkEtW5ns5hcTAv0AE0sQX/z0b1JMzmOYWosKDP
nTgPM1EySt5rv8TAojlAdAiC+rfP4WNAc4LHiL7q8vkM9S6m44mCa8r4NfReSfuaiCSDGIIxSD9O
4PPdPgPUPKK8zR/1ZeLiqlCjz+0LkjrGWPhUftw2zHMn6Sbg+/79qn+/khN5HSIH/UtAT6R6cMd3
Gc6XtyzD9HYcSIDyQQTb7hFfl2h19ulnTbarc3uX5uDwwAqDbxP7xP5sMTnfD4pJdGhUNLg8QlL+
o9wkIwg/sDXu4S4yfoQMzjSq04sZI7bTGUIINZEgmWbuO0pAFg+fMXNklP4uArgSUk/qmWCh2/cd
l6V3Ar+XE8GJQUl6ZocKXYHX5QBSV/J3ufl4xCGf8eEJ/flzaz5SfBm6Dvo6XOK1UZBVkCYBenU8
nOC7ewJQGOp8d+GKClhe8pbFQU7KcaRbOLrYvi4gcff7C5R46x8leYOeS7+qoV2/NsBVmZoU9Q3p
FvJVSb7vqw6i+8M2tvt6YWBTjNAnWQcETRRIb01bPBwLHqqm+PQotpEMa1Nbwnoe7wW/wK+xRGl0
5VzviYjBjlNMZhytP9G/5WoAcF6eMnMkx10/svwYH4XeHdee1qJAY1Tj5bVmqsubTebUOuUeRI3X
WlI/dwMLUD5HP5l839qNy/DyOOV8tgUfQuIJkZoUvpKc3chRAAZ70Wv0by+D2PnJB2/ZIuIvXQOI
IDRVGmDXTbM9HN8iQdQQ+bubwiKdvsNFLe4t6TGDsNG5bEqbwZomP8V30vqTkCDNilYgPYWp2H4L
9HrzURgoXWXgBeMgWobR28GWeBZKfIFlfbedVqpie51YuYIVd6nALXi1nCP3FNCyYSWWoLfHZ1Rp
IHjM5eM8x2Jp4+Irzrx7j6+2EMGCWjJ16yPAKDIqea4MeyZXrhGsGO9izNr5tmU38ZON4dICVF9/
B6oVOE2Zn+qbLMzHQOwOL/mP6yLv5LnRffCx2IzfYHA3LowMoylOgr4v0oPn4lJZIRzjkZcaWFl/
55SQRW5053zTxY58Sbb4fna++qGy4S8/oE5ZUo36sdj53xaeGYG0kXi2lsx8lvnFOuq5NbFbw4lb
8u36JlZFHNbPXoKt+vjpO2jZtj1OuMqAFzZF76NY2GcXH7hIymJYav786BH/6VxHP+xKYytHtSFT
h8pSwVI7BOHKFbB1DHIiye0MLBUniU0PRUGsNKjHLVz4w5g35TrKP/WReUf7RQUa20PAYjLUH8gv
xw1EhqZFpXeFSUZPGGJ8XrjYClVT6Ok9OPtKX7Nlt2hjGB49V524AavM5ezHRLh5Ywo0Ph7SgoAI
Wt+6JzkJizQRW5/CKKKBbicOZW1mF7QUjykkKFxNlCGAEpAyrhrZdrCY3LgQM/SXp3AYXMBP+qYJ
gbg0uWtGEIxnkC94uly9gknHX7t4pBhVkH50Jj7zk0JBc19SA38yNSb+i1m4lHARqKideObuUULB
E9RPceQKqpJwfCgEvKy3F5Z+qsOIrNLAime0DHEvw7K3Bzlesvm4WVdSryKfpACFFG7+AcoWMYXm
6UidGwMI0rR+VOQpPBEXlJGpWC6dyAxbyafiZgkx53p48BB5ybmOa1MGQ7ZU9o+73X5BFGQmJjj8
Ww5umEoaijM2kwBiTx+jVO2Eexlo9BuRVbxL+OQhn1TkHXKuZImu8+TpEGEvcCGZm0h/uG3fVFMi
tNGETKxSKCz297kr1YvoFNpbJkUgQ1X8Og9FlY/aIFeIlROziKscaoE7kJedtWySQdivM1MkhqoD
icbWNzdv4Kkv3Jts0Bp8wYXIJ4F3SWPQZ2MtnNcKtk0nEyEQ6q0Rpm2OlR8Qp6Et/4kzQ7TZkL8c
6w1Q1w7FAogKZ3SrU7vrl1W29OGqPJ1H6FiQ7o6hnc40ypLXd+Fj6KNE0Mqvhx2W899OpUNa/qyv
RymFbXIDubAAJsO0XiZbD0R9g+0ktm+4NEMODC9Cs8vOdYtGPhNCIFkmv+hBCsWmenCHQaebSdo5
YJbU4PMdXbTXbOazQ/N0fzuZrVpbrgl2rHEqb91x4N6m9ao/hKc77Ln5e1i4WCBNQ4r8cigWcc4N
ZYCcfNAFozVyvkg53eas62KeAZN4OBknaq9LUMjsO+01xO8qNNYiiqtCve3entSay4BF1LILksrs
KPiFGXQLLIxM0s745ZosVLQB+r09hj1P/j5u8RBFHYqwjGpztgv9OTQ0CBZ3wvZnc5jeYXvgSTFh
jnSzCJ+4U81NISzlHB8xbQs/s4gzVDUfTC9SrHgnI4UTO4okYSSiLohHwfeWGq8SuBqEqX29WB7k
2BsgAnGHDZHJ9ejhLBQiZYi3qgn1/apR8AF5G5D6HsPBrUtr3Gx9ZShQ9gmZo1m1OlUCxvf1iSiF
RnXjoWUI9GcNidAuZrVZVI5805LCGNR+QFdHJT8cRdBWSYMkyqiDU8Xuo60MZG8kHKN5XozX4j0v
e2s2e7NzFTND8P0TghdujCEwG8peuKmaeaWMq600YQ1NQmEIbka+J/IbMreUUUHfh5FwJNaKFXnJ
MJiN2fRxGGmHDHCxG8z20JEvqfgqUNJ5zniS7Vhv1Mzo3a/3PYZ55uyMDexrGCQ2pA+3ZwgsXuQ/
PZiBcVel4W7aTOxZ3zfDORyocLWUZIXRdRoK9ahCBDHLjVh1XjroVI+JJ5JRFxbT3xIiGTaOx5p9
16iceybKFLNL/AyKMGkHCb5MCx8iuA5+6Q74MEwIxmjd7DXCt26zU0uwHS3yi6TM0+Wu9Cuf/VQQ
ywqczW29RQUr8ChnLpMiquLoTibgyjvXk09vPGdTBgHFBtMd2BXeL9/t/Z9OKjcHw7fjwiCqe1lQ
z9dKhzzxdgv3TwkiUu6hJ7gBEpJKDtD6qFabO+2Vy4+9LC/3kf0E65W4dxa5r7JhVQAYqfJLqetG
FrD3/4rM4gwhuxQdwwsiL5bVDC0y2otQGmQ5OFjIeqzPZBIUdDoFoEQLRbcBrhphRRKW3CUjSQ8P
gIAGmvVXP8pZ2zN/e8D6kzCTvavFz2n65JYrEspBhB2PSAd7rrOkX190d5dkF6oJDC9NW9/RadI2
oO0NLKXGZ6dBi6sFMcyE6kNI9IxtypjFP7372ZJt25RngRtzJs1DNt2UHS54t8wtL0Gx/bmtPPgL
1DYWjmJz6ucTZ3+GmbUF63o47fbHycjqdFgcazNOMS60GO5DSgOf6zNSAXVod1It+JQR85OFN2IK
koOe1znfsviO8PRkd19HIQYppq5NxrjwIeeOJTXRrWbcqU40K9PdX4SsSyU5QfLXJfF7Hbl4Ip3I
f8X6sK4OJGdmy+VuFMIHbKroyMzZ2eYRAjMz/dok9y0Pwgp7lqpbhYkZ2FHIADgrh1vd7YQOeQcn
7j28fMz6IK6qHOydMAaJI7m1pakaiw4dhBf0brYLV0pnoNWCFaskgtw3knyml7W5PhDUWpo+m89D
XbCXZ1VTsWXI2UZU8xn/70QO4rAzyvjXq7kvBJFipGF1ppjb88IoF/HGHdptmwZ+oGBcT9dyk/VS
AB9Do9E1K2lQ46/fMumf/ok2AypyRw4U35iRPuUmSSFD9PP927wB3xIIOVFc1GS7gJMJnzEGx+RR
MYkHo0rExQvvFNJSY7TU2qXa+lR50xuNj3J8iWDqqVkLshZjd/amTzQfhhipM67gVvuptQ6oK0tY
mkmpOZMpeqKt/e22DUm3cNIkfK0PdVUz2kLvyLY4E4vfTUt+DCgcymzSyto6OzIcmcjhGQ3+1sJq
yVqRPhOemrAFULSb3n/pDULNBjBHGUHlIeruUPP6oV/FI2KHOR9HSennXOTL3YN5JvujInuvwKKn
Jvui/OIGBbS4KByRxaWvux59akGwA0jNhiRS775oicPq5MM/wJSXsJBHmYy/oDDL2DVy0tzEUZje
ubXgevx3saOkZK7EGM8TMZ8iHAfuVn1dgwhDZbJD16zMdZCdvGJ8owG0qWoikyCdnZpBvYkuvUNW
RFmWLD5CjiwtP5Wlv/ZVgoYPZbfJCk1TzDL3SdPg/CTosrTGachxUWQBuzXtk63AfPqKmpGYQqrZ
XXYpJwjRoAL1zpSU02ND61uUV5PKrq+qHUIra9WCLIXzVhmNtckZz+qJ7PjiAL7CEh7AQ3KAP0w1
w4llqRsMhdC4ULXqbPa0FTNNw9vIkaTghuvRagv8b0p9gad8YVZWxb93fERGpdeplNTqJR2jvlDz
oPC2KaqYaS1uPuUvDjyh30vJ8oBro56ZfLSS4B55lYehWdHoT7Hk0CJYMOVuUsSjcfGHnFQu2FnF
BgAiHSzjR4F1z3ZXEOkFd+N/9lXv8lEXrOJ6TFR5QhcAQp+ItkgwaxXyO7xk43jqBESeIPccOML1
7xY86xgGYi+KATYYO6Zn8Ju3CNiQ8IFPs078R4BcpSKykCSzlgZPQgKHWdLwpLUBm5+w3XlvXjCD
5lnn2+6mFpMAiS1si7aN2P++0snaUSBX4NsIzx4vS0+h7UwSnJlhX4lVQZxvZi0Jdn6/WyoYyf4y
IyNIG/T3BmqdHdq842A8l5CsWC/8Ti1Lj54gq0aTCVZqtAoEMl3hKDt8QXp0YvK8VyxpkghcRpzO
w5bi57068PaZvAGMuKchrzUp4HXHpeWM1pPCckJ9gkxgrqrUiyGrZDsEreKtMn+83EdIEDIlDkln
hGurq4Icv+6glzK62o+tf5XKTmUHEmqPbA+730cvaaAHSHBWdhYN9oLRJgfTu+lGPqqac1nsBwrf
3giB3aBf+Gj35T1qOpsTchMM1xKC+zV5q7lZbNpr48UW8a0FocdwWQ1BKfpcNXKAL9VgE/53kJMb
OcnfgAOtDziLX1qI/RuySJc5Duvl/d7CJ6VICJVp/ZJ0N18O5jL2STilbJk3Spo+Lf0udiMQEV0M
fHntSCFC321nBD9dAdx7bZh2upxOySK1vnOPFyk9B4SSWh7Z7DX3jfOYzb8QxjqAU8LZFzTuq6w1
jBZ2SDBdF+JOCtsQ0j1KAhlID3dZGCxls4K5NlfWlls5ONQy3p2xMVSygOBQO9fs3Z8M9SmUi6WJ
oYmBFB35RFcOzRK44AnYtbLaQlMXYkLvPguSXg9Ql9JED7BWYx7/SWQegL/sRUaQMljgUEKw1bJZ
PxNTxlMRxMGTTEseGmZIOnfd5vgPdNcXbGu/GtVq+U2M7FZ1GykKrgiUhlDBjO6lZrNl7petCivB
fqRCi042P5fopg3iGFdkPMM/YoO9OftD687Fv0GnYl9r9ZQiAK5rI3GQkXAtYvXrxXygxPpTB3W7
aiN7cAzjR3q//9LubFsklXG/mBN/gWlM/gR2RMA3Om5yWC3m1Y+MhupHGZ0cJIB9VBt5RoHvEaA+
LSZShIkn6m3qFTuAMPb/uo6Pg2wAM362VCsmtvWC9TXO+Ix/sFqyuhzeQOV/i5iE5ArO8Tdrt7tF
Kqsf0/ndFejXxrMVcCgU5kDvgkELOLpilkGe3x3jkQufDhsCKdsDrbHZbJAkehAagiPP+k4+iYjL
jT7ALHsR6RUCstLFcIMO8tki19a2xzkXYV8/jHZFXdySFaysUR6yzj8taln1VKNJ0pDLtpeSyatn
oTd6VlBndTrr9Kdm17VV5gaac1o0wpb5dC+8lkjg0uIjgD7a2A620XItQsxymvHO5v/P4qrCcag9
miwgcFp6vuk2LxyOGNKm0v/sgKSaEPAsFHL7Z1zzPh9jKEC6RMJhZI2idNhe3N1m7CYS2MwXY++/
RlBXmbMoLhcyoFTk1uWWA+Xtu8lkiQ0xOBZBRI+HG2vI0Aru9k89pVRkfFodyCJSik6V2KxYJGik
b3xCHhhDLV0kXwp/V8GIuSNX5C3O+Vj9gKLsWdgoDEI6mtGP6UourIYuQSPOJzGPy0VHRD86xIrh
vUGE/Ua0qqK6dvyGDaWJDYC2bxCKuwXEt3Nfe7vMgb9nGlImu5khoXz9D1WPovBK71oS3UyrSgNp
t1XkPk9tUA8OfHh2ZEk0FXMIcypQUsEU2MP4wkGZgtKA5vAcgnXWDWawQ0lz3FOqw5I+tYPh/w6/
J57RGZK/nYDrqJzIR+7M/uEdkCYxbnedH1Nca/Fp/O8RlShMNE1MqatkcthBo1c9azfYKaD3bq4g
OI+d9xLoGp6i2mZykbsRfKtDb2V76QuxooX2Tddi4FSLDHt+yY7riU7fItdSHoDLvxze1mYPnHiz
eDT8hadyHEoQC/rtYcvvx7NplYXQMWHc8eQpxVfsopGhumMsZ+mLSOzUBLQZ98F+x/FGsV0zox4B
XMGpi06PKDdSjliZEuShZGYh735oig/mUklJGFa2VC62qfec5upAP8doF+s/QfS7c1gh6E//sFqF
ZcVk6e5+hEb8sc4wIZdBV+OBVFZmccOeXlnoV7f1/0lZTzoK3sVDG4Fc1aoeev4HsjRYoanK6RAr
iiBJWi+WDYk7kur6/DNJIAlqp9C52cUPPA4HJNn9OtgoBfmAWHA/1sprZzwyus96/ZzTRBTOS39l
AVUk7yCRbpBKpgpedWEH3wrLVc4hNQF9XYkzWi0GfvPSyLtRMoLOoEON0KwZn/FkOLDkHZst2iU2
LMt/FDw7O/n87YWiczMSxVE7vJkY3/zsCL3NWTm/vofRao1Lvln973fQMTHLwXYrl9+SmSkt6mCa
SGyVrLb+B3pPqhFYSdIptLVZVk2dPqo6Y3gQtVX4dyTM5MNftqx/uTPgJdT3gLkAvU1SGVSJeWNM
1K/VrRNAqt4bLIiqJdfV2AwP4UZhxQjUGjT8arqaM/qBCbpwH2vk6tGBZa4GyDbEdcwBFk6QX2T+
o8tJCkLIMNSPfn9jE/IhvK+9jCQuG1j1lqLReVGnKzIvZYgNCvmY3OgI8odKncWvHxeygkJHNetb
7LTZaeqy8WQZlm2xAkF15uWtVera2LexX4tCyPgi0SZxurAsTpxl7KWNya9p7ocbq+R7PABC6H4Y
wNlguvwzdUSkKSRQ/MeuHhPkGWRPTYRT7Xlb0s52ZUnPVOB/yPT3bEkFmzcnOpEWmHGBQx2D/G8M
U0lfDfr7Cj7IhpxEiKI5hbE0ICEjRumHlCoS3Ej+/xL5pZ3A/CT6eoBDVSfHFgm8Wl3mG3cXrHdj
02TOBxr6ZaD4qnYXfs94MkFq6bj6hZ99glcR1JdKpa47jg0vudATnqF3Hv9V6wX7acPdXNjnYRjr
29FvBei+vplu1MPkHQvdjp69Wmb1hvFiDnSaqnS8Xq9Q//FEeVGu6vLOH7RiMXjQ2QRxfCC8DjF6
RqDN7ZKzKxh9WZ3D1oagZRwbMa8zT0tQO0PHEOOwgN9fOEpAB3zctE5V3q3sIplapYYFjKjIPz8I
Cm2v3l+7puksC865uDhgGG8yVyXnGC8fnLO83h1FLLJJbT+2WfxOiN7ZzKglxYijrKW+D2p4Z+lE
PNZgkApdp81Pk3cc3xNtDVKcY5ckH2I349scCwGGZt9CWvBkPkBAjmqY+Ek2P/bXFJ50zPBByP7c
NvOXc8V13PKbE9CfdZvxwNXNMm2+JQUnJZhH0aads88RqoFnxhqobqNkvpLdsWxj2kKalzJUZgOf
SyVLkiBaBQa3x9+jQXBoA/gKC0rgP4WB+/bkkYWx39W9TKQ9sv8yjEmklnktEM/9VEBFX0TOgUa0
ueIpQ0uNUZ7qL1grhcHo0j817vPLwjrGnhPRhmUOsNxP00yXC5+j9N/tgPKpW8u3bMxmIyHzmfiG
8wj9f9DzemBSq8d8luTECJDWmarzQAifYeRHPEI5qB7uLeIM9TdhC947lkPwsj+DzYEhfANDXlE+
Vm8DshMCxYcWNiqKnW0Dm0zQrmuozOHyT2/Aup8WiCquect5yLZsw6Dv2qnxsr8jAQLRSOIT08vw
vNJ/baz9LbQiauyKqfDG84P1xoVZGwRQLkdCab+/f2elf8AoTTPP+HcAyz8h/v0GWUabyUdBOKnI
S/+bofcCG1v7rbXoIlxuja6PrIppfUM3cJ/lflwuvfGmBevpYAtICrvDHaqMJd8XHaCT2W1cyowj
V+4HkDZmlmYVjaDTxetk85SDJ2ZgCo3I4bNBFtI+soSgMkPUKYUJEPfXYM8hY03PFx+kd1jQeR4R
njgiLAsEjmI/JAs5gE6ur+5pG6yqgxrlKgz1qQRvP/oAD2+GmWWTdvSfO5QSb3TPNxJK2B9VxjRx
I7miUTZO0nUw4EUVVcdwWKF8FRB311sWVLp0+mjRh/qa8y94l2lbriYDrdk+qIiEcJc+rPQkOaDj
ubsYmkaY7az2rbYddx0UyKgPKtIToVzD2IPU3+0MLLmzIlTChiLZdao8+jYt+Nh57oZP+nGos4Zn
OCFkkc8zYRWu+uBURPDeTL0HAiLzCs8BT52l114lRoyqKhClVKSMTQPcOWauxLYERFc9ZLW/hey9
k4C4u/LNQZ6bEOTKICA0RSc6ZOXrPZ9aYON8LI8kkfd78Un7nZrRJ0Ym6ZDCdnhUTODgAw4um5AH
fidfGQme5P4LTap596+SlJhqsIXxEUkqwXx+8u3Mno64Don3jjJ08DUSFQHjAjnjQxeRujLc8QxR
XkdxLiUrtyWgrdKopSqrw6GkjgiF8M5UB8yL0dYuh0XsRTc27u768Igj4DPmywTb1pnC2ia0bXf3
tNOqifuKVA0IpZjMn0suQB/aZqy+BhI2FfrRrwDCSJwQySvGgZbcqf0Lo2xxeNlxMIGlON942g+5
n/dMNBRbkCfXgpXGd8Tq3RkadrxjhsYrufROfa2L1RDSYRANOMjkAf9Af4BQ6s7G8dcxSVbooM46
JAURQuHmfqdevSzBL6IfuYTuJSLGGUJYS88vWXlFGCfL3dgIL0DKF1TZDkLFP3mfNfB9t+t7Q/16
V1jGYwDS015SS28F78qRn7ofswfYgSA3p43K3cfglxCw1jmmviQNE3fG9O/Xrr9Y/nMNQfX927uL
L/zUlQzsELKVSvjiytNuW9NEShVHu2RPUk1AhOCY8LxWJUzuiqq2LelWbrb9CQzM0TcJDex5ggyU
Ixo8tnd/E0rFV4jh/L1CaRpaflGBXlvHa6xAzIOqbpeV+CMs4DFb11fTIAhYUwKArS4jdi5/o16a
m3Y4O0hF6YQ5k388R6+soJciEw2R1ew0M4tFFhskIgqfFVvPpKzdul0wVqbh4KPVBTx4IFdJpy79
gHGiSEDUFtv/oQ7KbHedhHxFhxlYK5033YfZ6/y1CagSiaiPI8Jv+WHi2VkpMIOXj8BpFtpU0T6S
ZIpkK/2qg3KUJlLfaQL6u9Wjtt96q+t3rgq5+aGsdIsDjKJSVrTd7zY0AC0dN03LPyQvgCWVD+1W
h5S19oahmZhbx4GifTf8TM0k5lwF7sday441oLDttQIKnM/o8yE753Xb9dexulkocdRifsvcVWR+
tztwXEN4RBs5MBU5effDSvLtSciUAk9VpAJQTCNN2oiuxK/jGh/zMBDjJDtUumrZyE+SBb1Pg1J3
v2/K4BbvD+uwIqwUa+lDVgFUg2GaKAOfI/lZ4KS3jg4tUWTsxKPPoeWcuR1gislQuvqTiOJuOCSV
FVmBUVFlEaifCPwZxW5i4kAr+uVb8m/DbrbAlpLmf2HcKmHdgB1eEZ+qpGzw8bf+yHsqq12dP/W6
cFPUL5TluAsZDoT1dIm5Gvlugf3BK61sAEuasAYBPUwZAebPh5ByurRy3LW/rkRx1Q/a3Oux/8Mh
/o4WtcJGfIQOfb81NFxs0dPg0tymBU6p31wq6Uw9iEogsUd2aOHo3J07kMlijQfhAYIaNY4zZpTo
6cD0ecI/5Gdw471Ct2JZx7i2mCoAhQ5YTxbzdskQd8ybjivl4Omc196PItjqqVuLNJ0ZHhIVK3Gp
frzfJIvZWcTcmYW0nqLY40Sil5NGzZjjjBRXf2UG+BwtzC2TBpzJymOq/xTvqduPGyuibNF/mu1S
0F1a3s6r53n5v9vJhMhuPHnOd/Mj7pXvecFe7Jv09v6lmxL2amUX3NN7DBKD7GtDW7vBxLPiGtQk
DuPatqdTIrTriwXU/KYQ/HCyEYCMPeJn1XgKKfHFb/TGD8+iODQWTtfSCz+fHz3PIVt2hnIC2HMc
Y0WkRleoSm+hXHo3E7QqnTJ5/LEMiigLLd1StbpELKbH//HJWPKdQ0FSrsZeyJ/3YwpVS+1NXFhn
D4EJrBDbQWwNpLUeTZbZsbviDcgEp7n/9DPBysw4KbHKs1FzlujWO318JRc3sfbSDY32PdclUDds
D+g/HpJdGrZofCzJJW1gH4YbreSDgCKKJer5pyYQWm063UcokBL09dzHWhaew8SeWjF8NiM49mgV
r4pdzmogA5nPYw8F6R02N1gleyThIPc6smZZAE/Zel6c/CO2yGPNIX83UT3hsf3NAnKxz6/A6X2X
MrbkQ5V2IdZIUV4uQREIyxbkKRm5/JqaIpi7hsW5weW7gxKGJ+ONlZy72odpebHNXdHCFVs10jlu
4vmUDCVwbTOHw1zIiPGBxHvVXr1Q78jVCuQUhGuWB2XyLupT/tmXiK1QjNiMH55Mo+/i+uOiCAvu
rzboTCIpPab3SKMEeU+iY4kHRY2YS0OWb3yBK7TnrSdoUvoyPDHeBO9YuYFFrGahiS4TW/4n/df1
YSi1I76dy+R4DknudB2Hjl+Zls4hQsLOCO61SsAeBAEbw3rzAWtc3ODF273hK7FHrQNmpxOAxn02
uCnpwcfwPHrvLlKC2XY41QA2cudwKuMcpxvYbvMBh0gxDjtQ/VLt/ceysWPwSwjA+4F1lBGuS6qp
/62Tjnj3IxfO0YtvSEHpxt/8H7RlD1nOn9Rt0vvHziP9Ql/DriOR91LL1hTNZpCILyybI9zvKH1m
1EuYBCH+NA+de/lcagIRQNN3f1kxd/1T3ywTa1w+A5asAPEZXNzkYNWMi6dBKQ4ei/FstTsC9iN4
c7NRpwM8dH+FX3SwXc+Oh07oxd5MXOGOab0fWuc8BzDLZLH/kbTGmBiAlJXdXJT4U7JASyd0rHXS
H3skk9FOLzBfHJeOiItmHAZ3alWxgy5SzLiQcOXWaINkFEF9TRqoNS0dLdjJqmiQRq6ZuInPyW9b
1x6tL/t1NDym1Za/3F+CO4uddK6Sjok6eqlXdfrLX2z3H5I9aFawGDDNcLnYY6UPr8GtL8xKIW+G
oIR+s0ToSlZh48+uz9IEIGaXMpEotL34GQ24wztrwCOMXhTl42aOrd6EZJskgYDpKHEOluf4+ABJ
wFg+jKTKuuqW7C+BCH9+XOfsQHQ8+ManpYjlWMBcrGU+4s1nue/X7xrq2hZhnzrSSRAzaPM993rg
i0f4L4TmvVANy5s93NUHkhMDCrRebHSC6whGbF/2uhXhs6vD89f2ugMAUPgQsKGJuHNYqSB26FhK
zHPw5httj+NE/GdlpVU9JJp3xFaepCaPU/xj1XqtEZAF34lf21dnvgNJJJK6H2AuVWkXTJ50iy8Z
7RSqayFAE2nS1CvvVrDTQR0vUbGuMPjvVDWzMc9ExCGLAoptJ5t3ic7gHJ4Qg+/AjsRp67gG69jM
TNGcQMByuoQQxhGOzqtcha0J2XQR94TBgMfBDtX+jal9G5oCM0P+AF6/rgVboRaR+I39mWmBhsow
E5qwWwZV33qEqQwQ7/7AK+9bX4n6qrwCNsmbgZ1D7mbUzCZqq02+ZVDaLYpJStHjSfbKDprJG3wi
AcXzp1adYBSNbl9AqvRuSVub7LMPyXmENSV36C5V3Chdm43hPDA1tUYpwYpJYn+dj26L2dGN1+RD
8Uu2HbiU/bDYAkw2HfHQKC+In1eiKg0RJjvfLkcO+HF9eoJaVdPltC9EEqOSD2fkcUlrqT/TTmtp
9H9br53Le/lS7wMzDb5pRN2NcUmXgHcTMQ52itP1S2YMKVRFmSVeS1p5NDpdp3HynxHCjc8P3PAg
+PLLs/0FomeO4lUHPWVAW1n7nFjsuHbaaneUeJZMkD+H2gzD3A4aRGZVxKLd+rx8VFL7b+qFBPdG
5mYjScFU7D5X0iGo/fRsLo0f8J02PcDt82jE1fxGOmErEuaQM/Yg5fx5hQcTigTcoO+4cyY6qmeV
ZTyd9flO+RudQKq1Wxe+/enW+mdJdl0HTHj+n9+Am/n0J0yZtlOz0aPIIypLZiGjr/g8aOjkpd/2
vxFt/Yin7nkjSq0Bq9QJgpFjCi/zeKPFW1u4Y6mUBcEwso/Jn7/UFccMioZhaolQOABAOqQU7GYQ
McHMR3xK5c9HxmNUvQc+HAPfpiccf5u8qJVp8sIEAUx3b2CnoRdyNMK5ofzY/YzQkwDruBZZUfBI
wWATlhQ44dltMtgK7NXxlJhL6U5WMRKu5kVIz+M5KmukGgnLUcKK996BjRJhVEGexFKKz6kYhHK+
4bDNTb8Dm2MOg1aWCuPPbGe5e2hPbVezT0XzOhN9KBBvids7UAToiBp/NiPk71w3Waxqg37PCz9c
YaUVl/RNwNL3vuGmFD1kvqPKgVap1KalYdANwNr1ZELQWfH9LkomkBk4bdHawCMzPouWozs0eTpr
V9Sg53a1n6RoogAQFlD5JtOpsb6W4zUMPNx279M7SQwV7RvKvjrcUO5YNA3jWMGwoMD583Yo4T0+
KxtPf6aprwd94KQtxTrx8KilzMVpcwqfki5lQMQ7fyE2Q4felCG39BmXoXOZbq5iL2+T+NhqdFeY
32kKCO3zmYbtMUghl23fyXW07R8obEy/yRcofQOvSZD5mwjFjxNwIz+HkFKEqtIzPXWBO2JXFwon
prdzZTyidebaugxhBXpWD0jyi/1olg5uBHKzlydwQKu6YNP49DfggRbuk0szfxivjCY9ddF5C263
GcX/OXKOtgqa/gNS66GmlPM4R1x1K7DC5GxzZ9y/bN2ohRgHRyY60rqsPARCJ/6339brAFgPwLFs
uNKYGPI0IWZdYhXY7Dkc6eNvdsKYHY9R+AcBygo/0GnWKnBKcCFQP6yVJ6MUZhRIVzY61GgDrJ27
3lum7WEzXop5303So8xFtkd3x4XQuTM1fHKaiz/PMnpZajFZlTaAKjbDlueNfl2/Msx8zjuTuTXW
8Wfw6rr/Khm4CrcfL0apKsP/FGzHk2t4JNm3ig3J8BgoMWFETmce8RCi9iNVP9AXa4emX4wR0cdJ
WjyZsbMqPjsfD7FytAXAiWLHci7dUbhezfr2v2czzU402Vm7C5bqurx0neHKyxA/F440ZoihguOG
fYjl7nUnB54SvSbdTa38wxZp+CdDk3meSQrGpo1fwwJnKvTjRWeCa7k3A02z2roC1OaIFCQ4EA7g
2ow8zYdBC+gXjd/mbN7nHtBISuk/GdNVXNTjbyIPw5BVBCXY6tBqaQHVsmVLOJTOKQIi52VXr9YH
w59sPn3hcpOE24XkHi0DW8Xk8gr8BS76Bof8AYQ8BRSwGyhdYGaNjiTyhHBAHmoiNzJijDG/aHo5
qm5o1iXfWazKmmz1V9NPuDm6Q2WGpvbIZzzXpQldlc8PP1LfnSm4BPCGYssX3CqacGRNEsfrzT6B
A1zzM14VR2/m27C2slybxgBQ4+tF+s76z2zvdgsRvNUJ5IEgWy9InxBoiWvFyaVZt0HFSPkj8ybO
54WIVqg6OQfdVTPSePQcQmP5X2O423vXFbemwiajRPInlz+lx77/ZnE49oXZMO5wVA9+Cn2zl1gJ
F2pDzf3jTF9MPcu0kTUmjLv+wdljnP5KheLlnDQWTv8OClmbNUy8qwZ4eJwi6RrWxZx1pLt24Xxu
N6lE/KRggNfmS7twJJ8CLOu5EAYQfvJXgeE0Zn5W+ZuBG6jZ2Mc3kplKC0dSqD39s+g8n/dbtQLC
SrLYP+HBIZNbMnfKDJ3X3ET+Xulj5QANEJoC4tz0NFGowu9l10+zc45MrFeTSBFV074yzWd/O2gS
Klg7bdjdm6FMT7e61ZGtbFRLF+w/xRvRdUlqpOqvBOO/4j/pVUC63Kuwr6rOoSkr8vFCbQ/2Fe7b
NsWnQUKZfCEo/AjCqd2aW4x5H+d8rV9QYIkyurFPDPQLBaAakKVId8wdbJfzBHIbuw7pwCKUhBsd
0HbzP7TLDt7RmK2acfaVycdpAj65JHVcL2DYj6w6rUJQRtMLCpF7yepg6yezdz5qVsUlKu0V8HWo
Mj8FNHlPcPn7oxEoepmjEfP1GsERdmwQHVQ1yhhBDEjvHMm3l1JK9dXV42XZBfeiV+1B2t7s07Pq
fXCMiKVa8QXchm+iFu4BiIsBf4XC7/f9x14FQyT0u6GK8usHRvZiqXGXqh8gD4TQgErtn+XFuh/U
P3ej0rZyi+4289ojpcTidk+TAtZ39Cq6BsdWeBJNcPkbinmrIrG+RKZ17S3qyogkj0sdq8qGq0CT
hNUrs2L9ranGlkd2weNkVj8bKsyggKQVfoLab3G5uMnioOf8wiVMh/evtruSCqpqwz7fAq5RcwOH
/B0lJaLy0K+9y0IZgD/H21whoQs2Sx076KvzE6he7HSs1d6el7H4oqJIYm/BhOM/fSC6w9m2qInD
Wq9eu1Zc91V8F8SPPwz4rYD7XdqiTus0Hs7pgGjTLna8wUGpF0aZEVUqAwjCVyywqz7z+fss8O3S
gb5ikHfTghFGSk8803f128ZTlR8X/ZQODEfPBcGpf3KbhnrUp6dZKiGJjwoo6NnH3VYQ3yOAhTk+
RzBrLcQeEtsmOK+BM0vD2R7+FMI0XAgaWEx2iiInyLW8nCLX+voVKQOLWXydCZnnZJK48wj94Rlg
lc7iZHapsG+wps1gvERaZ7YdAhqxsj+s+KuTqxpj5OhqvRQVo8OpcBmBZLwelD9m1WU0/ZCeW7tg
1s1oM21pxOeUSIKyYQNoHWUFvxCIJBZvjuXANSd3Roadq4Nw5RZQtvyDxmuQcezNOgYLPR+RVlUQ
qaJ0dbIYNLHr/cEC4GybkV4Q+bSTcYlRVZ79X0M3/xYd0IPL9Ow+nclRu51ZV1fp1Z9SG5fGKWQb
bNYFOZnXTInvjosP1WZ2SALU+xzPCcN3tmcAEUtWnYzIHUbTI9hbFAnEOizEI9fyaxU7yG+l8I/F
UYYF7WBgxAeScZoxkQeVZeOrAHtxigY+hQeUFtio/vhwxJgKjf91m+2tJKePR59CY0ntxWgxxytG
TKV8tsKik1cJGke4gS4NEqPBdyG0T7VR1d67cMoeAovJdYEdgPdWYEY2+k7bDRKxEkoSrRgL4DAg
OlVbYA9NjawLTPqrpGotoqZX8/+qfTysjOPInOwR/areCqXVxS93LTcViRRm+qV8ROy6GUXIW5CY
9WSPed6ecJRpzfsT2nMzX3VPqeq18DssDSF+lpeubg951ojBRe8LctH+UFR7he68sj0Wy1Sdf6+d
SPxpj8+L7XLcwJWaTCC7gcRd8H/bv+GUt9DjFujP1fFTyNXcWUzK45db1ROqL4bdeRd62/lP+SSD
NpouPfwOBXBX6mJq0tkPL2/AqJ/WtLSfxGaiVErbhRJkz4MSwG8Ih3uN5euaIuX+ytwPWvS1nhPO
6Jm3/Uh1JwnDjwn2+vq2bd8Trkf/QC1R4lCap5s9jISCtqSdSXKjBWp4zirvogisUyCx4aKGIAbv
9ik6hgVd9ZMVUQ9i6gS/lRbW/tZ52G15DQGG23s0nK/RaZ+IL73K7BgVurvQHzsmG+1cPVkKJt/2
EmxJQss3huUk5r3Cy7EtG4Xsjn2MtDxHmY26khccRQdmbSu/mLo+xOYK6G3lzMp8hHTGRXE0M6gg
od52AGrtqjgH90ePJajIwoQwBbGQOgKAYjIgB+WZgmejcBHqvy5BJkckOgXxnJksHjuzRt/YuApL
56llnG2jjNBvJ2czMjx82oNPGMgj7cFOqxlpOZFLye1e7aPmFOYgz19pxXLSpAV02A0FuKUW9TMS
abEi6Oi4KqWqFpYi4PD/zEXnSvM3hl0MnEo9Lls7PxS6EPMbvFmf9sNozJX1AR+DIL9FKyENCPVL
oxRhf7yV+16Q7QvTCJuLrk+h9Q9TG4EjbB2oyepb1vlA/df3ihrpNf28Iqhve40/T5rnD6S8EXJ8
0g2EjgdIuEk0fu4AO/rHGyngEdZmNc+nTQvN7uO7Z8wBwXASm+TjgR8TU0WauQbBksSieY9utLRj
eEY90k1VZWo+jY69N2Bby+8pyLdzGOgesbxMqtw2mScp7FWw8LJQPoUz1CGz6pOhl+CpGsFHBXdW
ScDaqQudRYsfS+qn5ly0fb9vMXMlMhYTAmGWIl0YfKcFWOx8atVxR54SRpF/5pyW3a8IGkAa1w8M
X+AQtq/KS71Bl/IfveH/iZ697hq0MO0F0/2mQduoK8RRve8w1AE0Ah2R4EQK9jelD4jaRKaXyJsL
/cyQJYCawFeYtkn7nnMdDxg/ZAhXyZnCCFwpLNuYC1qZkdufGQybOLiaK/J5QezxvyZKR/FGVSXJ
bSdE5wX8GcIvcgKWrv2P+neiULI5mZYJq/10CrTqoQxi4KEZJ6CusxVu7/wFqCVdP1rRByZnuiln
qPkR77SOJGWSmU3vWs1qhGYHbMAXiLZ9ZkaAPa4Knv1R+FJ/8JGUHSIpwaR53TkErQho0YD2UtRT
2l/D2triyPg/NgBY+X7GY67LPYvnrQS++AssTWvRuuZStBpSS3mxlCil7ZQtCdc538usokK+4tY6
XT9zG9Wl7/jGZb0L3IM2cXG5xH1c2cG1oBo6ILoMd9TXH+/F+dIi1JiE3mEjQfwLRhBUh/vIGFvv
pjTBG2d7KfuGPTsBlzoQG5i/LBY0RbMz5lae+MXNFZ7/dkPJxWO6SX6Jh+QOlRhCIPfr1BlwbpUl
MbWU2cYTJIsHISkurDsh2lldSI185fbp1sH9od+dLgNq6df3bOtutGfyxFU0tERGqr9CG2DRjZK8
GCW1TbWRpv0EFkIMztY5KUbetHsXb/M2r+A7Qg9TQZayH7AUj8HPr0dpJRhayBVkP33u9Sq1kvpQ
Z7W4ZFSddX9WCw4MsjdsQ5wGFCX8xDrOF3dBEgBypVIaM/Cj/RFXKaw3SXilhHvpitmLI06WohLC
s3R0TdFW6CMmnTk+IgxkntXrttBtZtSyFmqJIsBmpWLjkJAKkx4V+n55SXtzeEc9QiYk12WTSiJ1
38i+uiWnvFdlfHo6AULMSr/F2FcI6pAEmlZ2WOFKMSZM6mkJUdQPjlgj5YCr/7TuPRe5K0wtbRC/
Iz3k2TJyeyMbgabiFzF2Opv6Wd2Y9Ebkkeq4C+jczw4yidyYbRYYCxzR8BRTQXbiPqWzFVhBazHF
VNMG7EmJ+cd4YSMb5/2awVy/WBV5YZrDWHFSuqEgFFvsy0q5rh3+MNNA0E6e/beUMQeTVbfApbdx
d+yEwP6sFMO+EipqnEglNED1eWNOnPOteWvmCRshIPcTS2MiFQhkO0eqSbDtt+cNItl2p+mr8DXT
pQ2QF1/4qSrQyUTztADGZVYlx2SLmLpxilsehTjt1VMPVjAJ4ZDpcwOLyMf4FmWJVKKk1XUmpkf9
nGrH7AS/vQJDYwZQT6m3wAdN4fKmEtrYYaNDwRhkw5EusSxnpmRKtnZD0EbdRBQrjErA3uBoiFM4
SJAbLxKKVU4QjBvl1ByBW4uR5N35mSkjnPUwioyXBQfRQ344hY/cFADycVC9Qr3pzRufli9OYJJW
aYqsM8nm3zOtT/8bzYg2F6VggW4LQmUR9e9KrPBoWQv3b/lcIa5BWKkwASQL9PYiK/rdDRQAhscj
RI4wFiFGDiOEXpyXszWGp0S2vxqyODdaeKmMocg34awsN6MjR87GB6csG8X7R2wDw2r2Ud1D97k4
vrCrnfiAa9baaoDjhtN6Cb5/abfn7zu8QLyCFo9IhAMmr3CUknSmScGOlwwqkHD9fR2YccRI1nyC
UsTnuiJT1kL+asWADuRYigufmxz70R5bwkjBBNJjKTM0FtodsJ+ak5dAWbDo5TUXFG7pxm4Hyn1n
LQPWQ5rhImvQT4JYraZnQl9gbDI0WRF4tTrnYm3aM/j/Z38cHMzPkCgIU7AHRYiJ4x1KqrLDLL8P
5DB8QhBvzZHBRT5O9OcZxJumEliLZCG3fIt7y2VjTioJEbnLT7Saa3s/IsGWfOCI0Gm/IL7e19Zz
CXQs4q9mDBXDu67xdmmSFXN/o6QKHRXNcgfTZdrCqmDGz+gjp3t5OwEmBEfdUSeRQfUw3lh5fLi/
OGYSWMO7fwLeN1BW7wKAkiVwW2Jvkojv4ihT8GE8SLtaHdMA7w7GpXfkgm6JsUVuSihpBVG234A5
9DLNE6b4tF/I4jYW5A95rfP4BM7q7XHGjAxiapY3xD/fIo5BwX1AR07sfZHv/IUxjzkriSvROCxq
YDCt7qq2gqjz40Gk
`protect end_protected

