

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mZM+QkmBmYCY7NPgF4QadIitw8Eo+SIwG/ZLPzQSVo/+iaeH+D5UcymUJegYkWcUJho8I/Ca6tC9
BcrWLzqiSg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m+fC7UnOc3lEJdF6HAD+AO/yeZSz11oLyDHA0Df3kGgHhj+RwbK/SnWf9v1KZrS0pMJJUO6XV6v4
HlgXy4/LyWr9xInVKpipB37EutWXywoqz+1z6QQnBeEc/bFgaYnjfNVfmCe7b/uvzsznRxv4g49x
IbbwmYVPlJlM7RiIIUw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rDbHS5sy994Wefoo6l/eUEpHx+Zo4hK7RxI32sncxdT1Bdk5aKjGY4UEdTJnrzZnlUNeiA7lqAY4
kbOZOXFRZQqL/9cE+Eexju7i3W9oXfaETCK004ve+Hh7ccj0BXqFm2Y4k07Ne/CtUJNcyH0Yqqti
gCrOLCDDO0bLrxPHhJABOIcLDs6XdASBzfQSOIX13iKktynuDQy9P0UWcx60e6rMtbpwLXUBSYUv
U+Hu1UEMOHnc/WTTxxmY85cP1KeGPYOpLlkIokpXZ8YevtDSE+cd5cn78Pj1A84QhZfP0eyUXT58
QBazbLlAIfh5YqSZshCArhNLzWy46i+D9nhtnA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kDAueH+1IfJtZIC4dXJ0KOFeEyMeE64ROjlOQFn0YA50L5K3mjbOqsUNUOYQ3AQv/MDoPnhQAw24
ncqGrSzr22Eo3qkCBevBDcKaOXbJKeuuWwa2BL9gVLd8x1CGNKRCY9HgRWTaFP3bFE8IC6Wb1MQM
lh1aab6Hc1hCVUoaMZovDfA7pahwN+Ofes0F7tNeWWHBJ9HqmXjdNSIc0fhiL4oCkFYFKxAj7VYV
fvJk1Lt8t3eAqqFmX1wv/GZUSXH/T4wH/dtyGB4+Z9HiVEhbPwshofy5qPAJ1GyWuU9knKZ7oXwF
y0rW1H9CueC082UO0KJfTB5adMlR6IAxdDst6A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fc/3ZbRoeSBESwxq84FLKKHw5JiDREh8UGnn2Rzjhu2zXqMwcnjmmkcDnHaxqko+FpcFl3MSrQyA
N7dj5tbbO6LV2Gvp9gQHdOMqgogI5ZSA2MrQM1xkEs7og+WXFDOW2DzaoVNBBPY30Fxo2z2EdGkK
82BQlO03GRrZB8bBN/1ndJVAqKmb6I2LgcJOsV4HvHc5rgPq6Q89NS7JvmN3YI/cw4uWXXLkso+g
80AfqZjAXMw5OY4cWZscectXNx5vGHWy9fcKNH0p3fS7FRh1M2zsRrVvSEP/ygtXR3Jrf+/xqhv1
fZSqKqzI0Q17bh68ZGd39RDw/TGEUIOZg8lY1w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K3Ao/bH4OtPU9lcf8MKmR5SH3AU/XNzFMyvYN1Cvi8TkAqVSjsRpmiA6psdHUxQ6ChxDL+ifIZmx
XmGdelYbBZX2cseyC7F4SArU6gFMESx2kqccYUXXKgud9VEcW/cLeAiU54NEeoRjHzxfyykkXDVi
5FoCcUIuf1d/5LfCh6E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g8trO3AM2GKk54eXi8fG+FquVAmu50gIUwVjw4ul+0+xnhvRbginNickq5wikk4ZtP1HiuGxz/PB
o3q4N1Lj+w+QS4/JvRo4wuezx5vzkWzfGJh4N4eME2ziyNHCuxLEobWs8KEG+ilhltk1c2hvgkMz
JXhUTpJ6l1apI5+sSCHAcYvC7VVjjiCJQhk8YXIbnWX5GNaeHmM9sXw6q6MXafVhmkI7KkLrNLFO
9p/t2fdUw33+h4NQB/TdcR/Eksd0542M6+Y06QqjDbTR7KIjnhxELKh1JRW3t+rXEJOoLqsFjP7I
26tNqlayy5YjSzF90FiIpUUwtrOsZ1lXamVFzQ==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QwE2AalCFRTpm3aOoXgseW8MLMWLVbSa89zNSHS9I26fnur8dp1ecu4nBhbmdCiT6xN9K+Y9LOqy
eZa8uQGcMgejXddOOIOoRBcM4/c8NEJcAIpN5sedKHupwvRA+1Ok8SjcQdRLHuJbTnYBRLvaK5QS
6SSXFkiXv2R3xlZ4ji1w0O9Ta+AzNh+ntvJ1Hd68xxmunKOL1y/YY43obHssJp/KBybMaCqwZpej
yYEz8Lz8oeoYFaK3poBxJSPhygpk0gKOHf5FNHmJu4tB4+EqhHpANOMIxzKELrB4cS1HL/3VPJv/
uryTtzko/3vhXdbwZl23slwjYt2mW1vcnIXTyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99984)
`protect data_block
AglXNuCU3Lx27DJq5Ae/2soJZYou/aM2r2Z0qJ5hST8Bwbn1oqIMoXPNzcTyys0uUtNVQsWbg2qI
FBBLqu/4dUK55wgy2GtTm13sabjuxy3qaTojnltwMDuLNCybOq81pbiRV8T1peMUyw+FvAXtr1QJ
wyYH1RPtkNMgd1ozaC/3pT7rjIgNybO+v9cFY5aEfpNxc38fpKgVCTOs6wGyzKi0CcKfSeb6yGfQ
+7NiiZP3EdN6K4GgjqKWrToPEuaxuRg1E3S3kAI+XgLI0DPQ2mmoNijh9Vx42Zrwx4jva2gCIOty
NuT9T0OATlKMEYY1DCBgEdD3It+h9crZe6twQaayFQdSq8YALihKL4//VsA5bzJHuADlLZN+HwIq
M/be4Uv6o5k17Yjh6c2aD3iKh9JME60JU1BJfwjy/tdp5o8DuVbNKpTwjkon/Dun2FURNJsh+O1l
xMDvwx8bNjilQrAMXD+yrQFrtxetDvW4wQtAypoENEbj7OfH7K8AW4qlTzls3hYpBTGJA5wSfoHw
fpFVolkIVIHI3JS3DdXEBQn4g98qTNuO4jKqSaH13smfh6I3HOlw4rVwS61RJGdMLOSRYEP0RKM7
MDlm/6DLkncZxCiYx/4EqTQOgIjWl28RnT1ql2qGy3jkvTkzU+zW+JsNZep0G+qGPZdADMCOXRmo
HJnXvzil+tEL/46/rHL/YLhUgVlDX8ELfM5B73hAB3J8G+h2kYTPTbmTX1xW16BUDuSaIihHCQ73
ThArlJVFDxeyMax3gw6M3D50TcWyxyrKw+bNsH4yhofepzco4ijn+pn6F209SvN+G87LTmCdT7G5
pABzf6hNImr39WmYWYQgiXsfKn+xgj7xduSrOvXj3lmbYRCh/OSKDtku9B4RDKyA7GAWnkDPy+UE
uEQYJF0yNz0S9UrRX3CocC5xEy5PDjFPv3aHKPXmktQvLG8MIDQzNP2wiNBYLLQ5DqUZokoKEhoz
l6Mq5vdDPV9AFPrddvNgMEvbWBj9QetgKkbYGyuQioIl5bkVvnCOm05pbZxbjcu8lNk7ESxyivYM
pyF/Hvgx1rNNVm7JgtJs4XxSnKmp5CiGVOzkhy3KiEz5sstXOSVDF2umMvlIsHQI8xFaY9RGZFg3
SaQb+hxxTVfG1P1+nsp9FiZSSCov0vVmk8pqZwS1DtofzsNSdtT/NI4YDFb3tiRUnrXif2TRRhCr
HXIerTlA01BR8EbnbBpslS9+BOun+rmKRVy2FwE1D7fRmIwjJL9NTD16uzQJqItU7ZRkz0uC44HK
WAYbDb4Ra7APvH2RBr7BaSlIP80W47Kl5O+mQHaggLCn91vXd0USbZPaKtc3n9ScO/vw22yVXV19
DO9i+A1AQp1+YPMlK5QYIGFA4Dd8lrMDpI8qgO9juSS74B6E8wbbCrGmUERIf9zArmrX1H9BqABi
x4i68jUCU2Mzi1Y6FMFotH1a/ofqx4HwHIXP9tCcJWfdQ12vwSkKSQ23I1qDp8fso/zDe0fyCt0C
LIJz/UWU/3/6gj20917rN+k5s5ciI2g19HoYH/GdrrHtFHaLw0Vy7HeS2SmpoJ9X+SsvHVEEx4nO
TG8abs6t+j8+BGjKb3a0R/g+IQYK2SPonJ5iP1+ITnyS3ciekr0krydphp2ZuqVFV8BOp41EZIBh
saHpNoZiFC3ZeUFCljgbdzrExt9vIJ12XJBwaM/8BEQrCBpu06toxfrQl+6MaUIpeTfNY9vtPaLV
2JiSrTCrk3hDaZs20GMQyYRcO3Kfqcwc8S9yuHL5OAnUDUTWMVR6ob/Ata8YzKGp5DMGd4qAOPJ2
DFjmR6wMI+jLH/Evs5feNmy3tH2h/g9QM8XbE/Z80JSsch0ryXSE2whbSzbVAN39QmSLEQh1rwqC
UDjpEKcBCmrExblypPYkJZJ5A+phWAl4iiWqheRFTGspdS7o7x45miSucUaO3WX9G9A1HKkvnxpy
HGvAAU4Q43pwS23/eRkH39NUx7au3AtkhGjOTxBRgYJH06u48QeRX0eePiIStO7CBeriHCt0WXl1
QN/wL5cvO2AUoXYO6bZHQz/g6E5LQoJsMM61PlYUqWiATR7vnKPveKsZrexIR2oZ2/pr+gFNprDV
liEOjEKf3RoC6i5PZYPlps/jrSJczH6EP4QItR4yr4lmt6coB6CWu5KRrmFjZvkgNGoUZjJWDNqq
cJi0qJHmucuRBlMzioqt4yMI7tnHFnIg+gFLeWponEOkLDp6vBG5Kg78FmK1XjU/+fMQ3caGG/5R
vN4H05QY2iGoqDnuvAb0yVgSbA0TleZBZ+6IwtBhlniuNL7QKUItcnBNzx7GI8IrpGoROI5Zl5g8
+us+W8CguRaXYbyWM5M7SUTrFSNBYU5hjUqIULGvD8pRnlf2NqUemYPVyuuI1+rrYe9adLMfYN8F
jWWwK/xarT3RsmyWWbYojbdjAuwYFs4K1LauZN/BiDRKfQc9ZgVzilWToUHuejhoHuoRxkGJDMim
EF3GU2xAmEto7Zu842evh2rK2XJzjO+SOxUfRIu1k6bHGy0cFWHB0xR2rIHq5VTZgHfhckEvc1nT
DyXDVZpM2euVj1nW92LLg16/F+BgejcVSxgKKYFsjlHqUGNm4og7yBQkyWmwQfwDkgh7eQwjNWW+
JNBCuhHQi22NQtun/Y6b3CvZ9ewMxX5/UtCnT5hnWb8Ugt7/e9nbnMtNTGoc0pVbSDEs4bcgozUT
Frz4jlXUN1PZJoN/tpOt1LNYeiAtla8Dfio/wui59at3S1WG8L3FQe62PrgrXbJm6JR4u7YIUWwP
cpkDt8r/fZ06+pSxyeD0BYkEj9pYmvBCX+OUu5xDmSxv1dGTWK0fc7PWIHZYHR6OOC1GxleZys8p
7TbAbCHz1mo74EiUlkAHLnOX8yNbKqzwUsCEsKwDT9d/D4BfYpRLHkYJo7xmlzD4lDLUTBv+7gem
P7fFE2RzdrW7jm77NtcuLVxThrWzAFTXAOriNQZkbRM3KZbDo9qDmwndj6xvERzrT/VgLK8SXT0U
VNYtsYG9Beo3QHVxKq/JnTZnQkisJtRD/9dzxkj3Lix6tQT90WzvtmOX0RO9IlEbH0x0InQwAQl+
jGM/2f2ScdkywF2753dxvVal03uwZ3AZx7I4akwCn6d/GYPaCbM7hxrtIrtRaQ/EFLaGUgkTGfjx
HcUf4J27hLzDvz2Kb27ktMj9tJODep0udSQy0qWI/fticf6NTIK/4NN9yi91DNcEGPKX8Bwj0Ikx
QgLbTcCyVFW+/QC1+5QyvANQQk29otjpnAqR2sCC4lWPq6nrqWIhn6yNuRZRI9d0PFdliCXyM8ge
65tfCi89EfHF0QXlxUHQBvHj/6G+gxYshB2n0gKZ0ws6xWWTUXUkkIkfdnaGZva0lgLfqiL78ly9
kqLcM9i86EzC8QvVe1NFlNg24DOvazilgiBVmn0drrDrAdn39NGBZnBPPdqEeOh1VbsXmmKhl/he
Ww9HX/sN75v/jzXJVKOG5L6I+h5TD5M80oHdbIIq/LUaCSRbMPUFixGFqBw0NBSlc5j7ozPio5gk
oPGxEjwUrysAHzIam8gx+47nY0NSY0qRASE4uAf0BoxCMTxTtnkvE3xSIJy5TgY0xgZpyD4xvxbt
VJiJahC3PmJhoxpjGIgjD2Yg6m9mvpHouuCYAv05+YFjOUEyiFZSkpSC+Oj6BxSBmGqhjNPKuJpD
/tGzuudc430ePgP/gtT279cjIdhPLfx5WguWHQ94vi5+ztLRT8ppqiAbPgRXQv3kxGfucxXgFmTw
wpcg4VwLRU+vo6vgRMER5GjxfTMwvHjIPAS4HCiI7sJLV3URRWjKKsojWltSXEmeCEpAmgrzvSqE
9h+cwwpyKHrqzjpo0Gotk5DX+PRMCquOKVC6WhiPDkryAZ04YqGHM3BbZDR5UALJwN9er4sd9HnB
9oE+9+j+zR0i2Re16siRlWI7MQGLGJVWyJqoxnI0IUUHhg7Z5XubSNjOGvI90hFjVCBfcSffq4Pw
7AJ052ULV54P1+PXgdndmy7mar3Lzyn2H92Ff4C0HuAHZU8v3MObb7UaetnXztadrEclgjsYlVXb
AnZnc27PLk4AysIKtKUwBydH9O+gNWdzD68BDmGHezusOp4I1xjTLpYdmwqv0ZA5gkAJPhCxhC5x
6kJgIvUS9wvONWreBVMRasTl+Lctm7010pMuT5Ufwo8X05CtT3Wt/kb4U6kPznjaTysf/no6lHuX
y29XV902C5rYXpmDWjC2OAX5uaGk9L02bBH6E/j0Af9oJFGjj0EzyyZRnHdW9TPhjkVnt6BdsQBP
kENz4sOu4lxS1Ct8rABjPayVxmT9FICQnMKbA1A2j125f+fFJRqc9jdAnu8b6jy6KdaQlhpHMUMg
s6XfLeXl+FKlf+UJdaMifZoLLy8r8PNsXvaC0seRdjqqbZbUox4dgRdl+NlXqZzynWg+e2EQ0Nom
PmSSm3fNPmok6gW+VaPc+j3vZ47gHwidPDy8jfMtn2eFeaLrqWSFbBCu8t2HF34hTQesHF9lAU/V
yCVcAG/zpWf1rwa3/Y+bywEQ05+uIQIEvdFJyfI3UsUv9cRzO8liN6Vp+p82l8VJ8eutoCaqDlWR
eUTJhZwbHMRB5YO9e9ZsW+6OLCa6KNUM7q96da12k9q0O6+AUKbZPYJRz1jMctk9vNCKvpPPoAl6
l+Eo16lsScfQqL/zx1+7OLdRCKr1QtOcFlCnhF3zkjxVB98sui52Z9PHvDtltTRfDrL5sZBDDFjq
EoetH9SUj2wqfTUuYB9Vc1rk+QlKUhBnDOrzOfRwu4kFIcj3G4HdKv54H7fIpxHf5rTC0+lD89ko
fCMzBYowIYbWTXGhjLtpptq6/XpBcODDYjWAfr8aq4qG4f62+GDlTgzqohpVlJ5pcCbZcE0Sjf8b
RN3hy00k47O62FreYM3h088F84BnJgXngDDBEp4AjYqi6eRBJ7Osy5BWb7esdhE4GwyKn0AuHWhg
Bx4mODiofIRAMd+gg4QeUG6n5+M7teai+s3zFTKGLWrZ8u0JkSlUZpgAP9lTeIYsnBUqR2QcDfJQ
zXcT69QBOQBdicFmu8fQJCGkErsPXopW4GgSj1ItdB3fI8Z+YvPw2xg3ztQGXqbAKs92AJgUwt4y
PjX3eT5QoEOsSOkjz377x0+qXUQ2M8hya0+vG/3Qsrzke2Zc/L9KmJHaBTcAZzInkwIRp5tMRcbu
cTLK/IRRK+/hh5ZEAS+wLlpHhprHT/8G/Cwv9FUlwcjWRMtrofTylasHksdKCREU0gp+zt9rLOZg
iOi4mSesBtpRcs/+q+6hzoY49QPWCgZTZu9p9OcQ/4lo4UGYJ+52BC8s8Yc/mO+61gi2ws567I7o
xuUIjRGzUyvnvYrR8YMH23JdkN5vSx4PmYuosWVCzdbAV0RF9DVX8oOHrx87N6HIP3ESabA4+i62
dEolwsMsHAuGHNddlgiiCLaA7YEdY4CQkvXlJzK5EYneCwhz47gtZpVXc9Uf7owZOYKq72ZrRepi
o4Rq6CjLaatWKiHbRjz4cCQ+hYE7vBMDtby9+cN09OIjoPyZa3WpRW+0ZNASGi5l6T2vLB55Cb9e
IcSB+yk6xCsbVk9eOSt6XPTspjBlOb9jGaMFQBkVdlp5bRQvw8GiCWUl7vzpze0K72ZKeFYa9uoa
t8N1MRNZ4uj0srMhyVsbWhTefaY6B3cvF5M5JdC2bGVZ3voclBIGMteD+UQF6j7gFq6dAZgxrWJx
ArDGa4PYf52b5cIMdYaaVKeFhCk+MTYtGDJLxhJ9bGL+PG/QSZlt/01e80+/ZP0bOq2oLO0/BBF4
WtNaoY8+U30Efp5wmtG70xOIQpfBB21DSa5uKqCRk1MNyzqwybifF6kWMvFlzyn8DYLyx4Al6VAk
wbzTLEFG6sTl13O410y6FQJaKiKYzUfgGDcJ3J+I6fBXp0WT6bdxaT8JmK8235LIvlfmVo+gPzWH
b/qa0gCulWxqsuDxx5s3b8Y+odSXcH5HGc4W8uGc6dQSQACWzUGm/1GMigyMlZCBfxN74qEHCc+M
8NtBFlodscaBP0NAo8dsSTWXA2Dsj3kJgc+ozEh+S2ZS++nBtjzQJp8t1Tf/b8WEZLz/jEQkAVSS
VPm48IhsxwtckGsoeyOZhmeYJB/Sz7mHoqk3yO8u7NB9jyoGB6mQZbjDUw2aXgSu02fiJD3iJ2Vx
j/rie8outnXpi5QsLNc/GpIDpyIQTUJHU8bZ0ynAF5DsG97o/SiljCoIuonz6hBe2LuqQl5Dar/J
GGaP2OL8HcI4B4LdOARuExlV/lNBfgafswQbc8TN6VNTlzm61UMUjRQsvUjlJJ0Y7F0fGeGP1rDC
jEWBEF7Y+4ALSRGT47tZyK8jfWsNVh62fPr8DNiuCMRR1EVmVgQQKLpKmvplVe4BlULcVGZ+TlBC
CK/t80avRv7w8/3MxhwYUJfjAV3p53TZASf0YlT1WyL7gJi0YT/dnSfU0vItcn8QJNKwOwRcIm+9
s6BrgKYtxXYMX9Yr3SluUoFlpkh+WGjLUb3WbXBLqCgQdloke2DTLAK5RuNGvPek03fnbwSWPnJr
EW87nnjVabpeJY7FHSKz387tE+jfXNM1CeJprugOJkb7C/mLEkiCQZ2c5wiUHdaa9WEYvaG2ChTl
Rp6y6m9RPD0F4qJU8BEdpM/Mn70CRYUH/tUoAWY94zsU56o6AjH83MGMYol4QkdwxP6iDr1VAKzM
1STpPAHzcwiMYAFR3oOpTMEKBLxXkOAsrS6BSDavALYt3SGVyJkSgRJf7fuKoksZqg10HhPxPpZl
UGbliFXqObMjEO0i9OzdfGnfxn07uEQGYuyw4qtmsqIInSCJ280+YHWKgJ6uYpkaZMyJ1GT+DAAw
+rNRCcJI0fZ4BnwfbjUiwFgtCw5YoTnQTseuDsVm26TUKZVdSOxKo9vIuxQo86nwQyFi/+dTuoAT
ETlKdNxSWWS2B7pAB5vbomXlZ9Wkj8Bupq63otwWPHlvta3ehNNLzr4qqsaLA2U9gKZ+C2bHBb7D
n7yqO1qtKlkLFQBWf/xxAR55hBldbjbN92h6YlDxn7IqY5E5PztUWFXfwskakZ3SSA7cTafFWeYZ
+Is8tmNShpWM9gOnxItz+G4QtsRIh9KaFh255HMjVWUfba27cwTsupHY9+y12qKH11VFpGQxuboJ
jGSRDR8T+eWpJCTe+SdFYv/UT6j4jX8Kh5w4TTg9LHYKbSQSpuOHRK+O6qlrvibOJ8NsbKawl/AC
VrWPLaD8IYWNKQqkxjP7Z/UNpyV1+FxbQYBmwtLYL2/Ejty6HzSDuiYKByzCMgxyGy3OIa/Gyp34
pixpxlONjmHJAE8fFwu8YGjAxGGisXPkCkFjr8unpXLHHImz+vLLlkB87961Y+PL1cxLno1fXbHU
dB2Fr6kX2bCRr4Gunwgw7Te/moSfcDZpmNISopV6ys0HR7BYn37N1DSrq6Z12PpfsOrJ0Ugcas82
BL/kvuVGQtK1UCFKoE5FvPACSJJXHAfFJKIEbBjbkquvbP091tPeQQuKJ2tci64GXei4+QVHEum6
AA4aAVGSf9TVD7XRU4Z5AcTTFSynrff1YRll3ePw791ubtZzXFDZtnm7XyP0HFgyzl/MqhGTQZ3v
sI1a27yDpvbfkf2vJlO387vbV8iXfEQamFUp4BRQZTYMDFIh6GElfXr2jnv21B/iKtQ1dQZ5lK5q
i7Y8QVW7XlX+fD+av+X217Fv6IdJ7/rMZvc1ECoVK9yqUDkqysB3hXIjy2+zmSLuNTQ+Nqz4Ju/Z
1FOzW99JWyhI1Zh3HeWlDQzB2i30L7kjobMNd+sAfscL13LcFBdmePU4KKOrUurpjAB3LicwQF8V
CYzfIVsObOBrFX6CcNPwo84wQ+I0TPP8gSVRTo4j3FDyrc0T2X8zfAkTnAwxXFwDPSrmKtGmncI3
rUGLLvYcgft62XZhzNoJrk852d0Z3Jtqe6A7VPPc2612hZFgupG6Riwqi5cI5QCMwJCZ6Tmdt6Y5
PvCgsMInULZZ4oqn8eLQbIypeNv/Elgb7XzSNEgEBYvH/wVb/bX9AdPEas9BPDlULatd+2T0Pawq
aIDK/A1bVi7/uWa+2FlOstZs2OZchPqTPfjJmtLGhxrWKwRmxrCOo7jr4cYDDHEdK0Fdk2oasrL4
5uIPvYeuETeO0/0Kndecq5uqyET0B80k3SSPVYtEvM73oNIqECFwiAv64PHvtNM0Qzznspti7gf3
vdFAZeykgBh7pewJfPOOICzCkzHwWqkS8JWRdmGO/zGcKxZWL6mmGds0/HPxgS+Wv8R1dCk9hBeL
NaDSQt3S8nzar+v7MnoPukvXatrO+KMmaBSWEJ0pwf4Ng/oP7QeV/aUQIfKSVrS/PQ1/WRtwJtLT
mllFLHh4MVRssImC9NYyVwwD320Vx3PokQMs5TklbG2tn76/CHHbML7g3eNXxtj+HV0LPkMesa+h
/9AK2fhOi3w21CW65GbKSL7UNP8ipsj/sUV4tRsDJhJX5Hr9wpGrrq/7U7AHPiXtGrZxpVV1T2bS
ydHXb4YHZeql23oTWk/i1B8+4Lg5ybjTFikQUFSDaqsEADMfvPeM6NqvXjiJxRLoNrFbCx1n4jKh
tEqKMaE/zJ46KbbX7drWA421flAF6I2Mrl+yA36/Yiggy093hnmijnmltFq7dsJbwfJs9KEUsQ/2
LUiIvq98+umPPGSc5P0j729hk9sNphzjpG4TVRuorUIzjTK3t7NRMhrehgS2Zy1rzJkLjN/Bjf7N
Q7+YPS65LpDlxOcXonOh6gAEpl2WlxWq4pyZbPMiffQyyc+GAK2dtpJQ42LjDKqiAwL1K+2z895U
ga6bZllutfIcAPcqTf81mcaDdQo+Qz754m+synQnlPWPQdc348fErVzawmbzMX/sK9V9PSVfEStL
3qEBKxDWFSOCWWSSdQ4rmnXGfyjlmigr6QTjKcSSb8M8SU6NQNJA1gA6V/n8H3IJJNlM44RhahYv
GVHnfRO9tZVyA2rD+yNLKUfTsVwLJhE+y+lPFNUZi8F2j95w8ocBfOq4zZd55D/kT+zf59Bz7oft
f/PqcYviIDi7N/8aiVnZXOcH84y4ugcgChCTjLda4jjlM/WOQjnNcbB1YiCaz6u2PjXPVr3TLl91
gtDTdmoE1eGv1hbsWcg2z+DcH5NMjIGJDAC1k7gmJ488m5PWUpiBeAO1wrI/u6b8Oc78OkVnGWkU
FraohLqYlb5GsmtoaRFigidr5mEveIUMblopsTogwkTkwuLpAvUlnSRE3zIVbYCy4FGq5jmfqH/T
Lro9M/U6pu+tfaiAoeTurME4FNcRt/QInTua2xeEq/Kmq3MLZO93dClv6mHhrR1JzTnl/oHL+kCN
ZnZ8Nec0eIZPoMcgQi/V8nBJsaqt78CTImOZ6xp6iZmpqYRpWm9GU75wgCJCXhZn2YUjsX+vVSE/
f00NUglGAtxQVG5t3TMOhUPqAFmWupvXw8rFWcKsMTZnlbqmLHS88V+D+pTw0RL2ca11EsvKj+Rq
uckQqEYMVjEzS7/pifoVJ08ztlxoaExgBS6544HDY8A6pRoSr6Xl4AZaeoV32j/ARit7ts++uGbd
VIgwZDhIZ8MYvWsTOlJWlMEK7ozEAM9zj2ltD5f8cupzDSHbKjilkGQK0136G1/DJO9qE7VI2Ffp
1R0kn+iqXJEP5/u9JxHChgZR7pIUes8EuLKRCU1VgetkOuYbWZeWzhbD2/vdxppUabTcRVRCQAfk
/J4X4hw2TVVSXU01UeXXJf8YNXlevhY0Pu0zXlqyJUEPNHDhsIeiDUQdB5aycoEAXCVabbbYx6CK
0EuTc4f3Ycmw4FmQXNkKH/Tvb+hk/z7RRu2O6D6gh2k3PvihrJKPUPSVd/RkHrCjKGDJDS945AeI
RjKwAPPZdyw7b8N5DLYVJUei6FNDTVpFGjQdCWPgtpShzA6MlOvmnwRNOuUgCBDRSvdEeefYcm6S
J/z8CnC64wlhLIAZ/lyDj4d2V5rbOurKyxlVs7fur0q8aL2uX3Y0wa2CppZBJWg17sALL9GEJkj3
kH7W4CniyA6jZji2HSpYPbERuAJ5qOD0HH9RdXcBqcFRHG5weuXzmSXTnexbEH75536c7ZHv7TDp
pGN39w7C8ld8jYvlGhgq6WYHM11HDNMlU5m5rtbhq3wrFuY/BfArsvSnC+W4i44NSPtKj1eo9EhR
1Al5syRPMo/qG46w/xXoXTOZIs9y2NOZVVMnUauUNsYv2IO0h38Ox9nQtG4szXyFI4IDnIHYNTxc
G08TkuaI3yYYYDqZspVBEgREli0O3GpcSISrBrdlf9LRZnwbI4Nt5pgF/1OyCMPVg28x9lC1SpQ8
5hnPb5RhpsOKnMMDrdGRW2XSySWzkl7ZwEeEpU96yyylU62BvdcSChLxXPCqc0XBxIKx0pMgpMTD
JeQQej7jTBCkx+agUDUIfESI9vRp3MnvNlsovz9jEXvGyejT1SmQWynWRtIH3MUzb/KZ9vTowVuM
wbVI1xwV+YTEhVDRl7/GzeMdp9W6M9JYo+mUAlfmdwd3MpagSKQH9Foz8zT4CZh87ieKP54CVS5p
kY7aJtLkulBFkcnjHV46i7DBBNWdc7tyo094rJKnNCAVsVu1NhdwfS/RpzUgZtc7e7Fiv/8WZCNX
E8B0J196beGWGh+sWA2Q69bkz5JdSfxdi7cqOFPPddAMp8PKUVwZHSDau3fNNLX7NaKDG/gbeVoi
Q2kxVreu2iUotyiU4E+on6X4GOT4oH9Sp949dfjun2doRT66h/KjgFGOHf8W/9Zpj1E7yYXOfFDr
u4Elr059QieMoXtBqjt9s8X8bDLJwXWq+ydPE8at/ytddzW/ltNZwSk5Od4rGGMe8/6PPnLxXpXL
klfG0N3YSRuSTwvE2l8Hcqa6SG+os9UQyy+dbW94T3BZvogHX7eFvYLoeiHDT8AePakn3DyGBP8B
0rdd50Blfvma8/7yr4wv0xWCcAhZrivqzmtP3shMKNB+/ZyFbsh/0dfkHmNFxQtk5KGntYWIR1IN
utRM3b0vebfz+R0F6sOAPGaObT4v0f47bRBjcwtrLvWDaCrkMRrqF+5M0/zYee6JLNg4zlBdzqrD
5/indawM2oCLOdgBjtpZR0JX+ynqc4aTFBVoFAflJTS4v3zygV3Kha6jCAMXnf+Ll6jWYSyk0AUI
t6eKjL8PgFlODiMzzb7Jyq7o1OOPrBh7mt45lSZ0Rkncf1+bOWAOrbcTBt49E1dFKSSHSHOBxxhl
HeOOYlZVWSmiA+KqJNKir/5oaaEQP9HvEWiCRAwrdDHnmEPDWBz+RKSefzNZ8IXJ9uKCd8KZzU5a
u0oYddFmXbSKSms63TqPHs0yKqgS+r6Jzg9uZX3rMI46hyXDaAkPw68mt31hiIHTNiT6TFafhzeL
DXT8losoMbAIrv/K46MwQQO357s+7P8dtpLc1l3meSta1FhVnEYACzBA5oDWm9WhRA9Wiz9UrRSg
8Nq2nxaw2y8Y2rN06NEcDLbw8w5E81HOm9/rXARf1KZYmfK8o2mMpd09nWyppkbLVyGZZLi7yi/Q
QqVZCb8MRtOR5cBjYMIK3pHOhRT4CGxQQZwHUSWqfyeQXEP/xfB7UxeMzQthGjDifoeQuD5td7IG
neXAfBHgxVaAlqfSuR/+yCQ/VrrmlOxaOKTrLVMZI1+7ubOFTcbeJ+GBQRWPC4aJ+LBCinvjAYVo
DPPwDCh2f+nyI9AGqt2LVKz+3hM9Qk+j2l1cNxLynkqdtv6PPNApEGWxcHbrWKYqwzDJiK9zjVxE
RVy9D4roYh92LY3tGKKYygoVIYNNAhjxSQbAL/LiMsBNGIpTEMh/NjqLslfofnEkTNFe6Rhlkgm2
LpZ0F4mGOtH/l4lSj2Ze4gKTBePCd1Q9aqQna15P9853cdPc5e+RCFxnR8NgGszaph+wvjYg1/cv
e9Sn9eBLchR4LCP7cuHffjY1yI9BvKz1CjdJHb5Xq8Y+c7jFsTYAUiq5PzCWPKMEHZC8FGH8pU/x
+p3VSnsp5m4DQRUDTW+cMHO5ehT0hLrTLa9Tn7ciZNbEKOE73NGBhrCzeygBb+dKPOTXEpKRJR9N
pVJUfAzHMc8KnOL6WjSnncLI3xMWu19JJRdblNuu/X5C7hfT7888OwCUp2Q78Ps7ZI3cN5Af5Te1
P3V80m5fC9bAje8VF/6fpYPBDGYd5HCKqxgVDVFoqbdos1iUYy5/H4CaNHK9L0Jtx7WoQzAimWTd
G6y1trJ7R1/20D225GhM+67N3G9RaSuvqp9XQy8wHx0XMTRPIl/MbGd8K2+3L9oyz5PFzOn7NRoG
MGCCNkQ3Gy/Xf5CqtfrahpL/M+xNRBuRwm3EfXA/+4URc7bKzOUI8lZXd/FE9KYGrfHsV7rOuEO0
40/A1PJmH6PfV9+pq2EI1M/nUeohPMsnrUP4OGlMa7bxT4rMVKW3OuzU2YHsj58XQy7FRd+SvaS4
VahvCsi9/7IY3fXKFXppS4e+9hzOMIym2MxegQg1KRZoHa60AD2bJZJqqAl31ceduwWe5PnQlf1M
WDrHFql9LBYa1iKZfWdyHhQHqJBF1w4RQKLooRndZ0wV53Kuu68VZteoveH6jq+cOMNHhg5f0A7h
yTG+3SE39eYwr7OFlzbxFdcP90FYcrJY0Flwqpn8Mz7dTiyKLCVa2KivWoPTblSVd/387npC3fGP
k3YACP1JRlSMcI5FJx2MhGd7EroYW/LfNCsivo0slYd9IEGLkU7C1Ide8NkFN2ojL8xb9rN9WDq3
HE+fA6Pfgi67eaHmB0dVDyE0Wy9IeiBuLM08QRrPGIN5FMuTGK/vykLTR9gFc/HkdHd3uB//L5IA
0z0amh7Lo0SCV86b35gFSeyXBGUi/cQfkDwCuw6qx1zriWZylRZgNe4B8loH165Hk2MbGIm4Eo3J
z9MQSsNjhQW0DUxQ1iKTrMGxK8ur5aNwPchCvRPh6lmaMTWYeczU9+CDW16E0GyVuDLxoxH2uxNK
NIx9S1NcazpBZHnhAUf2ckivAHdjMkOKFUm1X/rj7K5O+1vOVPyC4jRon7JM0WHM0ATMobP4XDdi
irsu6QywL721TJa38eG0cAVZkmMeYizWyhfDSlAa36ppimqqthiX2SI8tRiAPN5VlT9h2ysZV4kA
A+CgZ8+uzpkF8oZBxx0I//oLqf7DT8Tj5x2WcV3PL9fkXoX5SaI4i8M6yB27RbLPuTorHnjJNyVM
mUVLjUaLfHqBMKBY21lxspU3Ge09QHF1SBjB6tVRSqSJZJXp1OuYxAwBgO8ZgqAhfpOAbywpViRq
DGGbkGN0MMn0zHzYYSDSNN5kDBMtkzsjuB7+N4znHq7RD0D3ZeQJALpD2CPKO5UzKiSqFJgq7yS+
AFTYVxnfDH5D4lJonJzv++EiXo+HYgy/ieuj8gWB2J445gekdTEAEWWFhrbukUCQaIL6Cth9lNDh
2bAbPDQ8QH/CAgGa89ikIwHpX821d5bcgocFymOklh3WRNh5n9UJdm8X6SGoq1C7QWtCbdqNDj/V
dqF6cjNzA7ikIqakG9G/w8SNHyTKCp+AEN6Tdl2HFeEPYV+l6ubL6Qz+bZ9pcOUvVZHcRwzY8zEB
TFfE9sYdOdVqHzaaeHOmRmzNHxOXypKMReIzJTYZRBHNww+ApuPAC8n53BSjxxk1UAqaDplLUxNi
cDA++7N/nWtwrNJQSYPRdunf//wPlzMY2sXpQsm82IoIqxxWw6Gsg4fW0JEZSE7LQLrAEeO0hxaJ
Do1dpkDXi/3MrVD5uFiKBo+axPWJyBmwxddnd5KvEnSoEjU6A5byPooDEX8DyoZiKidn6w5b2+iL
8oZHZeBa2nWX0L6J37NAgZGup1xaC2XBWBLZw6LFVa86N2CLdB6k9EGmZqauepVLXU1UzGQn97Zd
o2YqGIELIUR3xYKtVAK+06FcADm+JLcK6AFZbPfLqc5NVMOgn+haRugS04KRMEjFwsBmiImf93OM
qqYlowndPwnCanCV1piOOJ+FUusK9Konof0PyOxvuI6V+LuJ0ntgNmuxnDIyHNYUjNhE03cF5BmN
7mevULOVNaJGBKw8Qae07J5c5tKnulRy80Z9AEWHJ8rXi+ehUndlFGOlqWWGcNnVF6XqZcrOKVw5
FBV1px9tf9gy+WhmCzs/KSBesRGhLR2bfNK4byFLHjDEjjBMmMP8YK2t4UQ8mS3T52BMx0Mm7Z9u
FLZuROyaDRHZq/VnRWcaNbSTVi0g6RTGqfPwYqxpoI/+28mo49XzH/HGNI7njmz7LobWBD+cjyKo
iCb8F+B1FHVeGZSG03WB4vJFl9gDmSUrGDaAhO4Qal529/CX9pF8cpGB0aaeDc9s922Q6bQqL3e2
8utVaqmevUGNKckEJTpVxZgDUBeTONxu8upbvlONCoucK1sIUuNrs//tR0ytZtFyo/dXm6gRUcW/
qUOnzs9gNTAXhrQN9m+oeNMGQlvs9PyKG+A+C7p14WM4Yv/b2Uh90YZgXNm4UsN9RIq51u72Gl6X
DFe8qzK3afe8athnfaWgBXxVWe6DpF9lNxZ6YbrFQGPY7s/Dh3nTNngdKdKSLDkpBSGKqw2EajgS
D2xLbHlGGfzhM/ctZYo+uE2IGFdf3n0kKUMK4idbvSWPOQ+1TIGGR7sQV0o8aBC2nxlvvZjEWL+U
1lZQu6bJ0txzxqIYOny8NnqbaUiklIO0THfQKsauhGZio6VlMcnABZSmIkNqGkpvjXl9tLJ/oi/z
mMpyumHNmiGZT1ZNczFCbzl+WogNCHbv2FkdL7ljkwUHnFXxyHNU3rC1TSCUVTo0ZXjxBZHqdz5c
KADi1oq5i1qW/ASH6IMQiLmFtQaDwmHVgejM2BpRrMsZBF/Wl6mTiihfnBJEK0n5nSZ7qI1oeqNC
MhLQPg/1QvgzxIRT0Nzm25efNdMnH4922dd2k8xtGY+96k9qn0QS1myLpBbYZk6b0LLma533B6Qa
1J7U65Ui4eZkdB53xdDLsBB28xGvEMCdiw2UY69qJSs+nedN8qYmB/HerBh4XEQwHCsGQ+lzziWn
VWWFXAjCqEwFO/42ZyLIKMCerw1FEe5R/PhORjS74NpBvGH39T7YmtIRNgvRpS7sT+Ttk4lFQtqB
YOaLhNpg0Z/2zFWJRI3IpU4PP5rnFtiR9FPBd5KgkkPVsWolBrZ9/324GCRDogt1pTORcGY9gG+E
wGKydMZ1SMMo9bktMYzxFpag7iPv2b8IVF4rvJkoC9Gtl0qzLlIWoC+ZUC5B/2LOt5lhAJJF8IZf
LnDDTHagabN9sAA+aY3Rnh7IfZKHlh5cw56n+NpWUHJQUdHSe0raDBv7aPYwZ61+ZAWmyO9KYCzf
osMMGB4Kd+rRJIgyUrW0N5qaOBmicC88tjEkppW9BoreKmcy9P+nra9X+fTgPVQg5hkCogbvx+vv
NyUTZfK6824B+vrW3KrSa2AmVjZ7V3mHXatvRp2ZVcLyhBWz6wfu3kpQyusQjeP/WXyPPuqWeKQH
4cC67U7QBCJsLY9COldTCgay+wuPLrVJAC0zKfSmDqHtVaiYOQX+QPEATEmt5Rc9fZgcdxr13LqW
mOanas8LzBSW7CsGrbURuiMzMTBmlE/Sf05aZ4yrr9UdScK/cHWj5ZRRTT53XvAWhNpUrp5QFuEC
lJBEVnQjVLGmuqkBv2X7KsplxGrD2KTV2/hg1wyJl+Ue5joT0zMgUD5xkiZ1g8YaLh6ChtvYyons
LZ56OK6iK4hgFWu3lK1WeNB3rCTx9KFTx20aYz3a85eR2Zen/QRi37lOC6JPZUC0AohCwOH8kQDo
qT0Qp0FO2Dog8IGENj96u2Frfa3T3i+PirNQy8VELQ87olyr8fjFGWvYkv3XuKA2DRgxQULjJPNr
VJH/dIRpj8yIFriRZEZ6h7O79RytkRnDHu93ouoxkFyvQZqQSCaeuADLCuV1Q/Sfdo4ReqzDlBQn
hyTt9J0qAPxqQIqgYsaO+zACcAM4+oY55ZhX4+ieYYDi7NfvLPc89tkwMMnpzvg24tI//6zMLiI7
ChbfNChbNXg4WhuXYo34yOcHNzQAkpvPA0LZKGdn3yIcysPiExZ8B7uhmC9n6KNnGmsnUVOoRbCQ
/oc2StZDhypuzgmgC7YmJOsxWfhXL8howUv2r5KyHPRAp5SaUz6FuZwCl53eBgwLx5U6Zu61IaL7
iOU56dvAUpRxBtA24klWsSoOvRtr3NAZWG2edY0RRW01tzwMj+xdmeDNOgLMv4AKgZf/hQILzDcR
6XU+AKdH2KrkihVWnnI0kQoVaX3EN6OXgsatkRIup2YnPecSDYi9IOg9WkIKvwTobF9bCPKWUEWN
AqgnrtFbuOqvw4iCUj25q99VDSonxXJ1qXKeWOvnl9RTNQdGmv6A4Ah7/us9iQdD/18H25+j0wzJ
ye8ErMN0zYWmCFupE0OCeuQmcxWHItwCNFvGVv3MWC9v5fQexjC9ltIZbKdcMOVc3E02zDFVwJ7I
08ziA2hgyXMbuN7O+AqhZJZ7iT/ZTVDt1zhzwNKFfJ3jTNH03pW2wb49Ebdn5gjG1wz5ky9l7quM
ejtVEb3CJu2tK3V4xI/eGZB7DqI0tSa6eFHA52bjLD9lIH/E19YFbEkZIyiKnzzBL4T0jXtJXrWQ
qm3MLCatAhFN8LJDv2OzE+Ba/gsn/jmjbr5dl106ttVxgohanASPMMSWZ3QeRCGnjx6ihD4MdgsG
mtBt1XP6Un4/oPxLD9CVYc0c+oaScpAC2b7IztGSTVI8VUjiRGAeQrnfwwuxhBZ3DiMh//I3RtW5
9SJ90iEFiROYIEJvqe7DbptgTbaqPCvk+e//0Gqs24LGIfG2D/JXFCqiDfxmgNYdQwb5ky1FIbjY
UVKxlknxgXEnZM3IDuocR2uX4bQO6HdkRM8jYu8LQwpCL0Tz/nr8NjLYkkeHj582jupUxOWyi1KD
ZNYE5XRZxc2HCa0pcmdTDsOb/Sl2uvZjtWka/bIzOWkUmQyWtwVyD1CWj11ZICrNyE7NXoRZB1Si
24/QTaaICVMk1BQnxaam+SENmyTJY4debG++fj2NdfWrN+Vwdjv0ZYCYGJjtDNDEFDiUC9kv2e2v
ujIANObpGmeJ4dk8fvtqhuPaLHYru1BzohRtk31XiDKc1FdDl8x8xh9lo5qxJ/qpRQuRxeBtzs05
I7OX2x6LMkogkYXyaZJXrCPVr0/aE63IQp5z9jMa9tyQ+zm+sXKLw0F7r9fqQUSIU7dsbHLGpPK6
162J5tkLxyEpqQgl4aJ4J7vgonyXDdQwzN4zirYJg9NjPS5PcoFKZUja+F9n+Tk77ngFyyNvgJ0b
9ODcJrpNYxa+uWBwJ7cYdTUwgOMx3LS9Z1lx0UMVUgrzd8lX1sMdRxAXHhQh35s2rW38jA4TYmob
YWx6c7H3unjVxUmw2OBADDC9KS+P5ouRF/bVuILmxZMLxHJL7WXSuzwoOF3uqewCw5kDoxXkzOPd
tu3aFly+ZYjRXzThps1MfvE5+oSuwYo8hkcS74G+qlsg9q02vfihMErAPJ8e3I3S7vLoHw2B6LiX
6qqBiujemSmO8z8kSvPU/HfqWfKTMgU/lBK4X8b1vU412/tcPC1kwWwF5Sw5qqdYsDCTONgQR2po
eKCRbWL/NVTCveYOp4m54PF5Ud7ZKo59IdjuYbzmkkXxe67L0gLD2lecPU5jZ5Pvjc/5SNT4M/fm
A8sEtjqgViYixFIHJkwqMRNalh8y2pUclYKO8NHHNJkT5hv6ajUp0Zz8/VCaTL3N4qgDo5zdisoy
w51yKaPJuTNk5M3unHFSR7CctZ5gQ3w+nVe3WN1YQdyL6JfBYmd+fKOKt7rFd534mqZ/WWuh9jxM
AKHys/TVqwJhH3r3B+c8V5d94x5z6Xss+GAxoAT7Yc9mrsOroE9oX+m7Gdzr/l83jef/SMv37iqn
OBQ+pKiwUOy/wO/6FdA5HbxT+yLpipouWgOyGSyfBYJ0USLonCaaoT+b0jqXRZx4oUio/WBm6bY/
QH7O2QoUa2PB5b1r+Lzf4Psof7Uprh72HKVBVFCkUB25ipkEpUxNTucpA+14waTOvFI0jRQoP9Aw
hiFIu+wlZEoyMWQsLkr2RIsgz++SGFqp1TBtHZG2Pm5fvKApIukgJGN0kwcNT7qWn/n0nVFMelsA
ym1ofh++bUtvGqcmFBZIhzmxHrqOpnsmr/PHxbgycaDZqUzU6FMgN3BM7QAx8dM6ZNPx93boXsaO
e/VnapRIVqCQyzFRjwaabhc8+H8/TqdhNbTbPB2X1rYtMUnVUnMQRBQbz42b9inCunb2fKBQFgzn
jSgv5crdHvYr0NGEbZDQgzMC5kLR9FRWRxmVJVnpFriGqvST9lJWOx8bq4jEhbCPTQPIRBL7EfW8
l1pmQYW9Afixh0Nh2pODoFuL8C9iuoMs56RKRsc0m86724WT6XMi3qkA/Js5aSnHwmeTWQnnRsYJ
SbmriJCAquB8gnxLQTkeUnOHOK5yUJIJn42qSS0HkxN+N3xgKQTFwHiBCImeqsCGp+LLSxuuLEdz
6ag35HvM/3OuiQnvC/0K9QNDF8b8oxaBbGcPyHaNLATlo15vdZ+GSPr0SBooG6+Qj3pldTMIuR2z
1uf5StYO5R8Rgx0H4qx5HvZnw9wDVVpvjoUiqTTy+mfAmbKcw4wUT7hHS6ALOBRgG4j2RcapkWVx
cpTB8Yl6pLKSRc346o2EbnmqYwkgYWK2bTJYv3ArEVmJtDVn6qbNZR1enTBEje5yB05xdY2L11oS
ZdnP2GUdJPVJ2peX49q+W/Us6URAX26vkN02JdB0Z8aW5M45By4Te3I9+w734s+D/v0omVr7nPDC
HEPXEJmAXZy12VcRJn+rS2e6NPPwDwMiZM50UC7Py8W9YXcNObbV8f1EBNv6swK5gl1zJMgkUDsz
xWgtr06Ohqr3MMqbcAt8Cm2+IxTdcFSAT9Bxcpv3zrvf3GKkKQOLJq/tx/AqRRHB5bLZiWBGdUzM
OODZBPPb9rcr4Hz2taxRw7F/FKrM7evuLHJRBGj0NMXGJrgGbyca6ObPfttzlW/k4dDJ2xZQ5kw8
q12pKwNv9TaxGNuK9ddA9sQ5IA0KXheKTCLsK4jwGA5LixgUU0W9EXsUdWOenT8E27FdbotFgpVa
sX5zt5zoL/bDn2wBr/cz6y8W77+qLxm14oUogDRsYK+GbdA2cF9asw73IEOPLdy3htY/3YH7He8g
dBPb0Gw+lu8ypWVbppZeL/YNdybdsJqr5cS3WLr28zv5CPoP+PBNFLTDssIhmsu2Lm2Ile6Fplv0
twluxmmJcOHDZF3Au7SSpqNZ3PRfC4DCy17XSaNDUEDN04uhOhZyUxtOnBuGX+ghLA8sfTJQiBiX
UVEffP0andjmmOmQPCbWLpmpr81IIrqRm+rZBGVby5u1LnQPdS/JLpLPWDNghFFGXvk3n+WoCUQz
YOF+HPgV3tOBXp6vKrOtRpAQov3WCkd5Q2UwNFbeqbdn6D/rhRuRQbZ+npFFYJDUBHGO5sWV36WK
t3JeGIalN/eLsfCpKySEVzhNItj4XPLoopjxOJ8Fijo1PecMc3ItIbeK5Iv7fF0rXALloeKxIpZh
0qdJxiPJvlCA9phXez/A9nJoHAEnCsrDSu6/4VfYg1Zobw/WYZ3kMm5TZF4BVFaH0SgxUwa3dR+W
3evgbJC2W8IpT9BkFLD/d5Gc+X4hPEEbOpYbkjKuS+A3ucBqwgMrkqAL1UYamnblbeJale/bNmrz
xZMua3YrsFFm+JKmD6TSRNJ0I0bFjV/teD9BxJYYe5JqAdDCeEVCad5A3o786wJbe/aCjZoK5ido
VgaNojf+O7fb2hYf/x4BHLTu4r8ob89bQ7alORIci2YMhM93pBhcL+1dYIOepJfNV83d8zkd/tlx
WtWGlsM099fMLbrEdkad6AMLDVUsfqYTSSxrPLvyFe+DRoq5tyrLwFX7+1N9svXtO7BxDf8rZJKd
BS5xvGLwTlI0WgTXPT55sbIqobh44hdCR3ZBrSqshLrkk51ZDwF8tCSrJ/MQ49oY4WTcfW4KbNVD
EVBaCJlfPD+7CzrCKjPddRMGgdoSEuMGy0kqbJFE5NNHtH6/8+KZyIOoKqpN4eKZL3NRXueti9gL
73YbSyIiVcrBHWSpYQp5PgNF56Fg8tfO9p6r2xowqvv5mTttjra/mE1FJqQ6/V3bo3TTT9DdNQfB
ASHwh68J16VS8YyQJkNlvkacy+gRVc72pxCXXFMAO8D1lWGflO/C5PDtHsVW7dLnugF2rKl7mdrU
AWav/0jTHOf+jrMDxA9+kdBZnrzzzJDENqCptcAeDpULOA8YTCcv+qdl4XVRTV9f8KgSWv8wjSyv
dtfdXCQyrva5MtlAqAE2IKHVD4M24zElfAmvD5tg4tYcw0135vmoHXktXprw7q1c83pYgAdnn/qt
4oCB6e7oY5pSe5Ien9MlMU23ReQ1g6m32i2pTwRpdBx1nMXgoprQTjTs5S2FqVdd2naTyYnvvg/Q
mi5LveG6dHiOsCLwiYrUfOkgqlUjP9TxAvK5/IDLy1S5f74OD3+BaSVEoCJHqMnibqzz9o45ngTv
oWkopDW5Jr6Vuz4FaILv1A6/AMcsoOJ1yiEQEj4gxzGhHTjbIlptOuCA7GNPN8LI66NEbVIC2qD2
dPEH3ajvdOkteFlbfdvbtHWzB2Vz8B/RBlc+PY2F3btIcCeGTWE8HlV3dQZbonrSHoDhWRpBxQ0H
YqmOJYRsPdDLVV4enpAqEyWhZwMG+Xco8Ms2/59/DgWnyrCyIq8K1EXktAcqFtnqVJZr862BY1dN
g4uRpsBEj1FGybTy2ZVWJS5xwlqxNrBCRnRH7iphKoN5I9CnGCbmz/sJYbhNMhnsCBXG1G9PQG8/
cJB3VA+3iKWW9Ff/opUpI81/81pOaJBiGT9zK10JHvmTeA+eaLYZrtNpQ9PNMZJ/mYg17M9j9fRG
0JzffD++FP47PWjvBB8KxSQEsEugetUpzq8Nm6bKXzTynTb8kmWDcV/ibkPI5HZ/f8Zn/H5TZ3QH
6bqI8tygdfyttujmKLLx8r/806slbcbtnlCxh5wTOrFOQoThWFs+St7JMrniZZVH5acr+Tbg1xJy
uBUvetiYAIS0CnQO3Oe96nzni5D8dWP3GgLki5iM+udR+GwDPaG6i8q6FfBDlWdvwXAqZfDPPP17
FN6hQxO0f9TRdonMkB+atG8/5E+2hTM/rOYpc7yliCcb2f5pspAAtRMCDhbVpseQdq6dJfx2+sx2
4Pc3HRssoAQkTbZQqh3h74iOvtsurmULPcEMFoo+ojrywVBXIT3Bf1NtWO0ocR+zUxRp9jo5Fk9o
IKi4bNI2yMytpyn8K9INNZfS/58+9WTNvVFh1hb0H3tsALHKF0A5jsdQOnfDmc3+QnU3lHZqoqOP
Vyq1fb40DP4K7qVZOqnDvSJg9RgO266E0DGZXyrqfLrxpcEA1BCQFC/uUwCxDaHqyTJvXDmZvgNy
BiI+Yt7y7ULf/DRa9KQlJLKHtgi/A32dy80knmoXkkyZe1HLyqbWhHpXPGFKn/1OfsanTmmvEh8R
J+8dxTlhFdRz7gGIN4NmkG7LKSyFLHYJzNfabU9ltACxc3JBT7iqbUfAKwT+AjlPwXfko+xKS1B0
VUNBs5rJqiWmxcxr2DTzbmpJPZpMbqkFbSQ6fwo511dTEkxxzFhOIoEZaCh8LC162er6zjGYZn1b
/O1dqZufnFCNlruoYe7Q/HahpS0h2P9ZcpF4/pBhXBcqKqn5D1mAlOAplm9VGme1XhgWCiG4I+dz
l/1cLl4Wf/uVISbghm1kBjQJp1pph1eeBjpn/IQY1VpSXP9f5vK1dYRDwTgsr8UqEbY3F6hTG0MJ
yKtedGHO/vTLRq1ntTOp8i4YHd92xuhseYBKuFviZpR/WCGa8UXvLgkZR/mbImDGnNElmR6D1q5U
yZE9TEFMkDvAZF0sTKFgYH91taXDdOwGjwDJfpuxXv5grKvrf9AjZmed2kl3CfzsaS8mUoiOylUh
0tBHky553Z5OFnSXcsXN0O7P/NRoZMY3TiKdgWR3YKhPs0WHXnq9+PDCCWLq5MqrBcpQlDfoT1Qe
tV6iAuaU3VaxxuIAkW7y9E8evs4Z939Fj6Ae5sJ8fq9FsGHCUPfo4tJiuIW2cpjaDVGGLeVGLpvX
lajfhJl4iV/Z2GKRuZTykY5gTQLA8ZE1dyB5meiOspZ1vxlF+hQBzNqEqrtjO4V9PNCqAZIbGtC5
jg2i3KdU5iW+JfOa+1Cn6XcwjrnN3lpaeg15Rbzg39f01Z+UWYVuT82mCIsExBmappF8BhmmYd3u
NmuqSw075IDIPvw8JgvSXRtxr+/7qpkd1PFY6MnLkpxPnMEFzDaCQl523yQkOSue7zKTKvfXRMQs
upfalQHMq3ytuNuepG6R7w6CZ0bWJ8vN1Qqpe9E/xRY2b7xmuEYeGIFm0SkwMEAHlRrwiwQ1I2QC
9TlXFnKCUCtWU7tKblXy8p4f4h/NywFkQ7xzoMDxWo/BE0QlJywoLULF/J+A1aK1c8A8dpalA3Eq
1mHxAGxeejCTJHZtT3KvRqdO3xTvKJRI0YQZZL1XMgoN0YexBEl8bTGge48YZQP3/rX8Fyj4lZ6A
fT0WaUTnxbfPGWgSwAOIVrqVzmcGkObALTTzOxHamWe4g02NV7MlkP5YcmYGmA4jm0e0Apb9hwKR
1kRYFEJO/PCEnp0KIvIHd9WspaEVg4K2UP8KI7pNspAjEhiW/+8JknJuCbdvl7dWqJy3RvNN1Axp
6sMFEz4XFU2f6oV0uDezrE8YmuWahZBtsQrhyivbCbwiNzL5dRkasklNqquh8lMcJXN3wQvOz3zR
ROyCdOe8NRMUfoWoEHgyN5GLcFk0T1Zs4Vra8U50tc9DqARAqwheSZElkRm4pUrA528jM5T06nYm
6ynOm7ZujvhH2kIfg3cM2Ze5Jn+afajqMNW9vdjVyIAubNAfkihALf48uvnx27n6Wm7RtEqcU4Nd
79DfrTdDXfe0KQ6hX9YEN3HIEJ2/E0BVa2vGn9n+D6qhbCeupsrjKNy/gQ165FEeCAxJoCbCpa2r
5RKl6FjIJEqQIcuNDXRGRp8rChQ92ZOqDeMeGuioui+UQRacmVZ4J8O9rS1KZH5R49lA2eIAQuWQ
DOkMFKYwQZLg+7xRJ2h+tqOdiZsjLI/vhnKPGLxyF3Gm0XaFsRW3iw03JH/QAMTw7jIM69mvMjX+
I5pHVC1eBJGQ6G/h55/clyx0GOTBBlIncbdhidxtnPXMHhH0tpioWnSEVHAyT0gjCfxvwTr2ioQy
AET6bJXXfhpdVcaHxhxrZGaj2DiqNNC0qmjIKKUOBmUS+l1yUq+ZwZDv6KBgI5IETiikoedRNABj
lIg+rquaX3VHLXIz8IGJXzdENpi4iubfVT06zaYdm/stUpvPX1hD6KWC3DM3I71F9xNW+nIFqgCh
KMrBQWU9ZLL2k9VFYfmAroiNxHgQh8TLGiLeA8s6I7LWBOwKFx+bdcWKyP2J7OnJwXK/Kz9UwZ/g
MizPC2YF1zgT1kGs/JDy07lpzhZdZQ86KqztgWWRmQxEbrUKmPgvyQR/kzNe0ZG4aFiqxGrOOa2S
WRKTSztMFzGjrfJAb74g2acFlFhYmfa67XIJxRgJVWfCHZrEPOR11o1NF6ZK05EvoH333jGaiSqm
gNFXj1zOnKg81CQKFlrtFBtNsPYY9NbrSOW8tfFxn6d8NiR9JQPRuUAd0GJpVm9rRc55YD4GjNNX
Ra2CBvKNIfK0Dudhl3Wo3gHZ2xrenKTk2d+LxnorI+Va3iKNyqMU6SVPoaKDBuGLJp03rJKdXDBE
Inv9xSrAUUqHy8WouUaRpHYT5O4Ixj6X75eV5cHhd6zU9xQ0jEQZgwMDND5AdDH3DOC7rCG5fzp+
akuBYPWHv9ytIoNdoqkonhChdMpbS0V8LwDfIozXh/1wUitSTHD+BlZTilon45czNf0YOQN+cteN
zh8lbaMuzjZDON38O2qnddJcpweUkm9t/IMm1IhBktO8YfS95Last0QvVfCzCikkd5G/DMLVUx/4
6Q0P6BnykNaiUpBx+44AFhzdQ5OL5gFiXbfZiPn3J2zzCYsVlK4tuhejkCvhCwBJhpSgvAsEgKPY
Cb7xeBCVQl8J8r9TOLlW/yIcXSRVieXoMtmOPd1W4/dfNy2e6/JVafLgPO7s147OwtvjDcsPrUjv
MUPvTpkcQtgxQM3kz0RFBD/H4wPhhP2xLaFkdwQNtHTF/Xu7bbc7tvHXTwZ+Q6UHqg5XkQUjWeVJ
oCxlpFzOpXD/takYXwYzieil5Cl2q7SiE+O54YumfVQ8e9lBcUYMTnYVbW3sG1nq8wGI48NYRaAG
4aPAS0kcOZvJH+qBv9grw6UjHiO0wenPqkmIaj2qpxl5l/n5I6l8GQsJvPEeQgWyLJorMeWhTiiq
EDRR3Ur9LNBcXPTZFC8ZIhOQu1eVGgblyN8ZrA2ytDqzvCoC4v0/EwinjHFeezwBnGRqZ27kJJN3
hMT0xeqgndpZZIwe9oB1e9vWLL/KeA94zBSKFJ8BzAnFNlawiE6Bq9E3uk44CNwTAwVYfcGeWeLo
r3bu9I8nkdb6tSJMSWtjWWLGmt8YSoxzvlcefe2tGTmAp/QlfsuQ2gXM5VN2ptNr+HJ0F3ber0hq
f9d2cybxkK1xNM65nc8FT5ncBrOXSgCtL3igAyS8x4SknEqXnnEry9IPoRzCaMr2LvawHHy7tFUC
uTYGiK73tdoXoqTmiq7VneS6TgxLn4S+bsYYHrHs/APidPxbxj0XF7S078KGDxktPANsBx1MsTWl
XCNM6lLWosEFf4tZgm7GHIa8Tg1bJlSe9eE2wd/Cv45zrN/cSiQOIHrYguzNRWLlbZBSChyeLxaw
OHZWK2mN817uSsGXx1OOW/sE6nLZDJqn2MiztBFwJuayHWDh1mZ6FxHEsttuCnFkntsoP7Z00xym
fPm0h24pdqjFDWtOvooMudVd4UtSTkiTYELct++D6iFjiqcg5Cx6iUSq83upuMwuTsirSLrp0apU
fz16Ut7JBWPbNWinUqJjo5knBCf9DvLzkI8n20v4GBUxZxRcsEy/dY80qIGxj2i5DofdHzlpoea1
fh5c3dpsHyCbveFRUAnXhFKLc1MoCAi5JDAXhb0iZAeZfXJAMx48HbMWBLTYQhvkHPm+5ZtiAG2N
ICkIVBmVZFdUqyEZc4A3aN34D+u0YFk15OnpGzEMPA7YEXVDTilG7LXGloCpbmhYq4yGo2wygHpO
gpKRMI4MLEW3TG8bUflwTxha+5M6vREuGGz8L+5s7if3g/nXL2rB4bnk50McmYQBHhuyfC9+CZiP
VxVUOmi9EnVnjqfnPrLM9Pcfwreq3e4JgGWD9wSE4Vir5jjfR2J/4tgcCj/gO8D+5YPnOaOZkG/b
+ZbWGQEDzGudKMt4+iC0eVl+zKHKrO+JPQWL3tdPRn9ZeTVPrFBJ0Y95WLwt9tkxWNBfYsQD7ZCN
A+mE/Pu0bSew9LTQvVE7uekHKsO4aTFKPqB1LvXqr58H4q+xNcRIUMMzh3zw5/D/5SuAvv0jL+M0
8GDOtRl2BhngjVQWYcHYPXihpGL3kOhRH1R4lQhu0tBa2umI+hlGelYj23gGJBUH7SJ2KyoE8SDL
bmbmYjTRRsdntlip8uhWGrcVOoz2m/TsHKUJ5XGk4buQVew5SPtv8rYMwqYY4/Om289zHObplnLx
eXA4lWkMGUlEMuX2cKiDl/87a4+XI+J+Ii7EoHo8DW41y8Fo4kRSJY2/xzd8ZbhRtd0Nxzw/Rv0C
gQGlQ84Q7uSMzpCZLzS6GZs04sbt9xYO5WkrXrA9jHq2HxF6gvRTiSnRVPmwz7PGsnB9kMod++Cd
KPDpd2WNvuqEjoQ0eZ9n5zIjdBVBlu25Jaef/Tnq1+x1UAGVRg6QjJudDtjsJlcSnmyzKL7FnTTR
kjZ5MFGMRnZbfehGapdWnX/uVsxcdvae0SwrerUWRR8Nl8w3FoYm+92StmOQldmwGZMYBtYEEigF
TN5JXCEJ/mPmZvp2fijb4HkUG+/OmkElG52OaRBj+SNFppK8EadZZCx+aN1ofZI6wG9WplWcreHQ
7Qkuf3CBS6NqFUa8RuNyJvXwoLfXfMJ6Tt+poOw794eWr60d54fAkWxj4OiFX4qT0OkboDyB85bA
bFPtBNk0fZdwS3po9/sC2ts63hGOWV+4yKPp4g8F2UZ80eIV85HNI9oCvbAsiOwwVkyIQhizigFh
M0n0FkXjq4bOumi0Ld0MV+HnF4A3kBcTVdvTXKmawkrIRKaYJf0PJTpOx8ptYHUjxLSmAOuHwxPh
qdYvgCVwvJecqlZDOJbk1mSBagK7qJwY4boz3R27NMuTPLg085498TYJl2qJdHTYnQp4kL9dCkT0
UiP1pRxQd1RHdOWzjP5hbzUqXYIq8h1uaq1MqNph2LBYj9bo7sgJr5Rlxz78X+FS1WIEFTERWbQM
3rBAMn13dnhvzLU8+XbeHSyp0Wnc/1RjIO9eGKiQRZrOF3n0j+89Qbc/bCe3BdCR+mdfzLsdHKp3
dWyaeR20He8X+3/w8sFYdJw2RD6lrtHv4JwoH88UM8ZxlfROcSVBPt9p1eIdRvHUEUV592wvZFlY
/VXV7s7susxFgectS8ppVh3Pu877LEbASQjrepCeqmQe0vMx2JK90pdwc3YYDymi+dnagwswIxMa
5oUJOjZYsqSEF/6+ylVy1OrQn2EXJ7jlCcViv8ZKfp/KN2/6YXxuqk3qwMNYya6t9uPgmmwlgAO1
Ti2BA+BsZBFXkAKscNcuPRNo71TKB7Azrxlm4y4081z7aLdcDD9+NT+iLyAmlS3YILfaXMbAPUhC
nuZavP89zr2mcz5QLV0i0nXv4zbX34/9BjyNFYtrmpBbUH6hMWd2iOB/gj7MG42OWYeQa9/HyG6I
8pJhDP+1AJVaIm1qpuMcf/YNqZ9EbsKa5a2YX/kLuyhEpZI6NkgWTjckwKQvZiKAjKD3QavsoM6s
iVSg2cUx194bA2uecTj5gEwm3A8QDABh5epWowQi/69xWZiIP8cG9K7Jc5Unn/dazQ4lRqZ2ogBI
LXkY+k5MpsERfaxzJNUzflxPX6zd9qlcN4tyxtEIzsTBdx6Q9uxr4P4n1jZrDueqTJQbshuTWDfH
WgljaNyMjPC/MooQ3FcPcn+dVafqW9LUUTdpYi8s/4QlcPWiqteSSIIv8kinCvTiJ8eKhak8o0nl
LKZ6Sia8HA5mDooWlMtHl4IvUs5eBjt7gEUKzt2aF7g1Ji67j3499U04SE//SDW1JQr843MH6t2K
DpadzEG7inroT+Z427dMFF46k1lCr1pHXsSSJrf94die4TxTRM4kc+x6kItzGviwolVATNZTC4ph
eDyc56xxcynjUo1TKW+RJcezs9OO3xNTlYbKHZnCDQgel1OphOJP0YCk0XWkVaKG23swZYEllTlM
Xhg4CzokeaJSwAMEPXXXJS4zyMOPJwCTFIzgpTfiajVZ8hW7Mj5us9k1Xy9oc0Flp9Q19jYzmoZt
t9WfNQhxh24/FMXRkrX9LgTJe/u+FtanHjHeMM9VLbMWVTb4x4eIuneMa/vA/NwEyaB13AB2PfSn
HN5bxDzCWFZfK1bp3fThCLga1KmtI4ipAQ24T78GHEJK6vIxMANkLTZozKnQj7wVt9nc4byKzjC3
kiLRYJT73BEvHCdU6SvyshIXXXq66vE7lNuVQCVRGg9moc7I1OhIAWSA2wTkzCTswg1E6kY9CbjA
HhLuLl7vbAfWEJIcdRak0XPHVoK2RXMH+y9c9+sZPfvLXVb82js8V6p6CFC8BQgajK6kwIn58F5Q
YMVRjbgpg9rO/6kxdJLg3YIIGWD7MMHjmQ12O7uML6lUe/uTD7dwU9rFkHuguSEhtU3IIt5WFYGJ
HMPovbg/Bh4TQilXLxSePIibveye/w99cRis4ds6Ni4MqHQ5eZN4L8Zo9RoHsoiKie5JhMxL30zC
GK7P0ZbyhhcCQw8r5ctWXaKK2ZlYfJFPJHs2z5B1RRAmpkZSKdZlUSP3okVjTjE9nOUCjSOzn/3Y
9H2eS2Up33x3povfrO9O7vA/3TvN6q53U/GeCtD9yyb1SbCqLWkw7Ot0gIHbi4D1cKcslwjd2v7E
7aT9GIbCme3oveCBRV+AvNAjx7yG5W2oTj9wH1hlutWuo70xNfAo4KWsEnxuXKgy0Vhsfprs+vuh
0KwGLZaiJkBxhYT62/3zjWzooDfUYFBC02pmbe9/KCbXFihqpLqddKnCdAm7zSOQVryWEPLohvJ+
Tv9HeCqmGTaDZEFjSJhzpUs6qqQHg1ln2BAZfBvDWqeTqnQkyhyPpl3rvupFPqnyqzk+49JbQNKz
9zEqZeoRk18bQoGl4Nj/btuEzfp8/WFIjXtrbCuEq+/65Ugr/jyXdTYAIpFfuKVYMZn4Nhfru2Sz
NUEIVmC/8BoBTCCwcOtwPy2hvnePNi4wWYLxuMJiYKXsEcm3IAgazQmfJgU71UG18YAnEOQ8Xzj3
fb0J7+dL6YPhKngk0d9dh/8yR4Y1jqI7ElVzOlOREuDJkXg+OstG5P6iA6k+8ojzT6OeFDKZhUYJ
pOc+QGxGOkRI9GBK4ta+wgaPtrUPrOrmsK40cvE4znucq0Aq6X061jLSvbGulk5RF7qUVOtST68D
5gHQSuxQfeihsXLcCKap+Xt9ULJinjRlIZrgGAbPdSXNelFiom+UGiLzomttqfNk75bxtiUwvWzu
DgroKc/IxNLSIbWO4xWHY1dOoKTSpd4mFifUrtYt3TiCz49cUaHQSeBgXFPkLBeTM15owoq17mMN
c/zV4XyCBt3sRBv8j6UYY2wnysPvdfX4+ULlQShnzcwr0VcRJ0CIzJQg9oonWakygU103MUnsvev
jPNuKRHsxuc7VYhDzjAJ5hISLFkMKmacXyVJiE8PVRpRj1ArdwMzDggW+J7DowiuN6jwp6KbRzDz
Gvu9CJK7dSNbFv/J4Hr7nnSfpCcT/tcbJBlmdyxuKSJEBzGq1QVvih8eKi0pw7Y7loy0XaIiXjBs
AEBSdRtLQeNBy67piLKiTnr+xoPg5slcVzpcGPV5cCwpVc4rykVjpmnVplnVnqK6lcoKeIwezAj3
1ygwQpGOMzJzjP+Nuz2Lolw9upqJhnbtH8Mo8UHG4+B3L6pCfJAuhJJneNGti36td/VIADN+j5+U
0v5rUwsg2lw6bRVbK4dHnUnns4kq7nbSKXtRR9bh+0IupQimHX/8jSiaPEZJfmGdu6tnibCXlUHU
8dVLkIz2EuffZF8xVQ/RHen+M1i4XrAzFmL2Y5YsjOrSMRVJq9634EwA25y7faa1j8i7Uixmdt7h
jffy7P1FI+YDCcnw/AFq9gtdvQCuQDgCW/DZc3BgWM+dlj14CsJKK+b3o/5a+wy5T/lV9xJ1dvaE
RaTuwBAjoRa8Jjpt+3vdu7w3hdzwWl4psz1mxA9hpkq3kmQ5jWUCp3lhSQsWX1BeRP9EphAiDBrx
NFpkKmv3eQ5M6K94NGc8BykzElQXNRZCweaP7lJKhyUwGlMxBV3PUq9wXCUiSdeIsJjRQbIppqxH
QYxAZn2fKEhlAkFsn8BXZUCuEMRHfLtjjA8d1lJudZ/kHUICJa4H+IMU8aIhLUwtNc5/MudTD7hi
e7ZH1eNiKRgN5UYNZApxgxAWHM1+t2FD70RSgiXS2LYrcpt2aULYZCuTY+/G0pk+U1O5JCihwWeK
OSFhW7sBqJmLVrBYXSo61m0vf5q2a8b087iMya3eZsww7gyo3Em/wE+FmoujZPnKs7lZSXETcji3
oLhDCL1KLd0AE6AIl4QbjqEHnKDroRTso5H7KV8U/+rUC36Wq0O5qwWUqZ9NrM3zRwnpjBBNiy1A
ec8PQ9dJ0GdQe38H4vBJA2EWAZ8V54xQ5r2+IUYARg9xzWrkMQuW5771Za1BegXbRTv9sRbWSPEk
wcZii4q5NPa0jN47+sJylpoErlIe46IYIYGhtEc3CgYFaDaIX9lwpzFCKdmXDKVbgAJeOlKc5vz7
hBdH7SBYp7b4GCXgJMhXx/4pR2q+k/3MH3XxrHC0bJlBxBBUJekueXyLL1eQ3UIPeSXT9DJc6p2p
cdJL/rwLStMlC4EReN56LPd0659PpI3k/7pZLTBmNfBm/XFFhaSCe0N9zTWMs1DW9nXL81uOgmw9
8onneBnIrZ9GYobScQ1vfzGv2Q6jfSYu4a8vYIYoXFkP44KZ02ZKPM6dJVLM0a4AZnAY/KX6Q9ki
K77OKce+7IzLn9LztpFfUeT3iueAJRWzeimfeUykcQwFm2zaNW/DeuEEvUlNUk2Qekm7Ukf2P0Na
bg8cr0RKI0ZOhvES/xfVsBnXZmtnR+OHEArz0G3FvxpN+7lHJ8f4BryI7eqAckixYqD9dCl2bU7Q
+OaZg2tNJsbOZiqAAX8efPseMKLFs4rfgijjh40dZKz0PotcCuZGWYKCgMV+DeaEA6AO6lNipNH5
8IoR2mCo5h8UCfTTcIvwwDwbTSPx/iNqaO3rvdDiSXDA4Ahsk2kDNW2n8BLl8f1pp4pRzJoNTNRr
8SNByp8+VhRXwNd03STlu75jNdUjX6yYtmNyF5KtIPj/JHhqP2ZAJ8/hc8EOdISTNJSLb8uJkqsN
7ShPfUI0K3pZPm2a6bn20lDBXLYwD7aAn3eONqucnXKZIHNg5uuBXQ7h+fNzoEbNpIhnZ8wmm0T5
PpYhCTTD+n3aib9xXwkGLy8sDlbtrmoJdnbd1knpfEu5uL+ZooZ6FILLGiN34VtTK3e5GbSauRkz
7gpKJVhX65i8PfzEMyHVGOtEtAhbr2oTxuAMTGi7/nnBOpFEwp6wdn44gnXVXtRD4mb5yPF3XCbz
8xEr5IC4fqoIApi8qRWLskrhePeACUDywMBKG4P5bnRK6Zd1pyuQW4wYPUrfPIEhaN+byQpwIfba
gga01tILMxTbk3aiubYx+BPKVSW4+wZPCa2mgj13U0IDhMx1ohFY0LR5Mixy3PoYQBGSwL6SAsOA
qAAuws6ddM5h2EMgMJgMmjgAv5pD3on4wsuCafxaXX0pB1Fo8l0QYLfx5FiNJ5j8cHdMie5z1UcI
BNzObaPYSla1SmAxXwGuqBEb5IH/RfZQ6UElECP9ydz909X0Ou99DSrEfH57wNL9eh7rV15mdfIA
VNaRlQ1UhdRmeMCvdT9U90GJP8h1TlJ+Dc+FknFEwfxR6EVNohfq51Tzr+aB9FLlLjREqXiBZhJl
mL73X2/gz9nkjM8+PYk48A4gfaRYEjp52ZhJQTAEqoCiZTTEJVtGoC7opeXZuaB218xMv0qlCY55
uwxZnXmWf6IU93j/uqn6J3lUWIkb9U81pmtZJsAj3083vle8CjNP1MvAJTTktlNsKC8LUMTHlgVF
X8OnWPhVx29r3Bxo+7tx/s4C1fJovNSVJ42nN9+euV8OPW+qpx2zb8b1AjMIY84sa3MY2TOX2PEQ
XL5vMYCYqMZKIgHsbYAykSiDVWz6Rkb8/Qf9JKo15zZKZMbaW7bQEvEfhxlGnvEbaLmU5zozxck4
R26zofrwS89z3N88R9LPIBpofYcEsh9PgSFDuleZHoh4kjaEA/8wsdgKtJ77ng7n8RwR47DoDaYv
6LRZ6ecXNQl6E7sZhUH2II3IO/mzj/p63DNdbVKO+O8lie9GdF6CisjcEVMzZYAt68v/oQVQebod
3hZwIirOHcQaNOk6eNs8WkCLHZ3Su8NXdmVSRmzHfiehJIWqr2eb22VhjzhS2j7iOLwfyZjzhELg
RQGXZXEHLxJJFYs3hx+vOVljk9c5ZC/EQlPWTJPZVmUga5z4DCnSo5cN4//fjZ9mnaO3BdC0Bsv+
bfTnsXEb0jmYU1k4vQ9oNO86UjQFx7XHBFMFxtXn5khi66u1dqSTdinsdPiJIvdqyLzjYonkXtax
sO1wKolxWd8TtwUy7ri1w0JYl14rkzMpo2zGuJsFa0ufm/1HDbEkCgnA0LAafP2I98+cs4DZ/g87
dow9ElgkR+aHCQ/8nRj60ruGQldb8bdN0imeWbU3jMupGiSRL1xzgNnfPKiU9qZsj3APCnVIUg1s
YFE+jEow7QmXxFjqKumseJlhSZ5Wppny4GlJomBPzhQtEPmaQ3FXDhPFc2Azob9qNjyWIVXcQPZW
FbPhBaVW6DXjHNNcMhQgwaHLuVimPzYDsnf2QVpzMcrzMut3KAkxGAk/JjlUF17vbP3Xwqh4FhMu
QPXtZNnQa4SnNPQYu1hnybpPk4gp2PUVOHXySj3ezUKF4r7DEkt/k4Jg3ThpS5c+P0anmz6hfOBO
pRrqkZtAGrAzG7gCnp8VgCzTb3btbbDrqiKluuhkE1wOUYH2nn15kzG0hqYm1Qlv3/B8qSsp65o1
tQJOr+D95oWcYzPNVfHo1IDxzqsNY3kJz9G1LRl1K04dIX6tl+twh7pQpxp14F45U0bLx1U4LHPI
HhMiM605ws3xkRw6q9N5YHBFFvINC61NdRh2f+qZHGePnQYdrmrAYqOGLWWA8wu13rlMXqAFY1gy
TQ1cFYA9X2cgecrL3r8YUSPNcp9p8Y3cxsV+b0KKq+1QNqUwllJMIA9Vuh7NPJBQ3pyLtQT6oBpB
XBef+2MHq7EjuZI874XK7J6d+jAjfohhjufztlCvOzmP2rw+smj8Uai5TuBc+/a5yljG6R4p95xM
nfvKkrpL8Ium8PJAueclkKyx+4IGWLMlXtgIBRi1g/PP7RFo2uh1A3r89czY4vVNDtIrznuKxL7i
1lUhmNdVgDnHc/yWr583CicZQha0pd/3uqQJy4kQLSY7jOT2fJLULELcTie+x7IYLJmcuZvSaNZv
8bCVfbgkY4tScRUtNC5cXq7/W3h8YZSkuZyP7AKwFZXnJuPsOSk6r12cNKkYz0uWZVWwhkBnunuK
JOHT3ZE2QV8ynhc6FSIX9vYCEXnITe8tJCuSBajjJe3wd94dsK8rh43OjNVgMfhr+sE0LQ5+2RzQ
0U3VhToxVDl5XVus//YLCDNTk0CSMFrEUEKM5JO8AFf+bny15MQgW58zCSmn+bPZxmHt5o2Qepo+
wturdWG27BTy28JG7HZtT4nd7zqsbaRIU2ZYaEIl7cdmFpDQ+DZiTyjLOavD0SvRx6BJpE4GGrln
afQBw2f0INEHIjf6m35AfKOP83961El+8SFGBszsV23216hg0IBi3roueniIEogRnpmOzdGF7IuU
9jdnAMoNVMxUd4qiTFG/RG+fj9ztPryOe4rRMugoEo8vpmfyyEn+acju0J7z/VEEVora1EU9z4p0
tbF7We3t8TguOqLPPqlnNw+Bd7coKXOi+6o6eM1DlAYBOV8Mqo1X6P1UTJmp/cLvvCsWu4g29xuJ
z20NKyQjNwb00Wuh4IkELdjXA7CG6v5Hxu7PXoiDzXXGzET2i0iUhLSevsBaT00xNXIWV9kVqeBX
dNuruyJ/ilo636zbNq5FZ7BM2fXHd19zOj1InNSY5r9Xwtv9gOjpNpP33Y4DFQWZiBmuh02ruiKO
IhwLf9qWH+igATSG69NygC1+ihqWDYVE+LgWArNQhJuyIB+aToEqxwtVWgseck8VtSMd/XX8yr7x
BH+d6L3as7WSkq0LRtP9emO6xn9MyAlyeOpnxgfCs7o4wrjnjuvYLeoYK6lwWW5AVyJxLovFJV7n
pcA9le/FZNmE1w62Uwhd3/7LsfhvYcZ7TVf3mWfSAYK9oXiGZkHTY9/nPFmZo8asalyczB4Vd1F5
QWj8WSezG7ewbnxAT7fby6QBWzAsfFgH6fOqRGSQxftmUkSEvqolU5YA1plQkZXQlPAt201U4jjm
8FNyOWsd6K9DPEbU/BJoCylKdwWg9CrOgjU8yj7Wr2Fwn7sxyMOcLbJhZrToZ3rXSKzJxraZ+VZ+
ZSugHre+iiHaoYMkMiSxsWqomALTqAZpmKzE6YMdaz6ILwzY9M4kMtRytwig7Ivfhk87S+9iuz9d
qTvWrHdLnxNQpFeKIggBaZ8BGxA54G/D+6DRO5HzRMiWSKxrSMujuWYW+nER50cVO25P+DF+SHq7
4oODBuxIKkq6KeSAazoMtyo0lQgYARqQEt3pxJAbt5FraQ0lYOffQvp7aJnDtdAJ8PRbKKyZU5zs
10fAWGz9bVd+DwFTBivkqAdp67JImsfnSnl8Qhb3AdJ6Y0N1N5cZATwyCPybN8/YiCt28Cwh52tl
+eEXwi6A39dp91XmvDUXzX2Zzbj3JxjXHOPQdZB3TD38+r55WYp1VZs6N33VfyRQWcrVBo4+2MI5
QPN/jPbjfKJD/O00Bg/NpdFYUOPWuhHV/rwBwzVwT45XUguCHuW+PS9McyZ1XWZ0a7k1eIyMTtY8
oz5Cpg8jpVODXhYo14ipC7WEMLUaOoNefKmo4UDLOEYLQ4rxmKrVPGfWKdr7T0/VTNJ1eOmc52lt
QlamuRl3bY4l9wLlUWGswjYazztWcF1JVNShVCsg7Xtw51pT3KahSnzjPmjOsKnHNnUVeIQx970V
M8uCXHDdF9EWGnvMJhcWGumUTKZH7fpmk02CyXl8XBfEl4lWgHSMNZHH49dk8yisok0KEsbrMAn5
s7Hk+n37ur8ZG5DrOBMVtJ4fONlYGsSPs6NICJYMAqflFq4mz7eI3NOrnIIp/84hq3kZC5e2nrbJ
QvFrgWCI50siS/ZOi6Gb0Io/TGqe6rAGAbzsFLS/9DMghbkQr44c/ZC8oHw5FwQ0i34AidxHYjT5
SL+dbhrTBaz1/A+rBd6Uf/0AvUleAGqRkzVp4KWc0PDiDdsy1rzceHWLIvtfkXb/mdtkbN67ZNQF
r+zki7QAEtjsfrqzocY0PCbJmqgEvdV9G2ncP5CTJiLqHmAEMx5pMJCxKQdstYDNlW+pDciAcI8c
JZi8adrq6fBvUWXOP11C/eTeh1iGxxj1rb0qvo0cEZX9rnahRXVBbmhg9Hol1iKuZT1ESSa6K3fI
DX5m7BdnTbcERUYB7JuDeE/zDJfQyWKdsWHXZ+MYFlV6krWuaznZopBBMDt0eX+Zjw2u8gyBToVn
ZxS4duHpW/LCo4yTsEExUDEMjkcnOm+3ftJe1wMmJ3dWdHUZh9u421W8KPROkY/GcOrLX1e1hnQG
2J90GPfKa9bPLWDjQNux5AlaxolsZoar2Mnp1fwn9WmKlX2G/qzHXXYr093DhLYluu3xvgcrbPln
SfJT/cLszD7+PX+c5HNtrWGH3TorUsLNHlKFQX/X6VbOdxWOwZL7S0tFF9WFIVMe81ZDWovbtqRD
y3ZqQzHaCMBe3vReDuErzCOTbobWiOrEaGJKImlwwvRNAl6H4bzvvdXw8CJnSfLbEYNZF0T5EJT1
Meuf2MXAJpW2jvNAN3Prk79X6Yj1QX20Wwm04mzyob1T5ygLyTOF5/DsWFtcqtdQAj2IGfXTnd6D
s9TfflgHvoz3tDCemi589K/S2is2ZKnME9Yu0Plp8owT2OVSLHXY06eWJ4YnNilPTBDzWF6LOqQZ
Ig9cTI6h0oCYMlQO6uNVf+f4XGO2i3dRMCmE3s0jAAiKNwyl5wk3axg0fkvLEEjnaKpwghT5KdoX
SbvAFL17+JHmWQNKExhU4o2yvFDYtPwZojzyBB13l7d9xxj+mzufxeu54EpS7Gu8UhWjl7zir3Zq
eW9y3/invZ9m81EpYmjpiqJf7kqewQqLoX3M6XKGCpAQjsve1CIvSjVLv2mrdMefxl4agpGIZlUu
l4Se2RUJQCV1w8DeMqjkzWVDuz5X1KmVgd2eF+yrtx7yXRSBQQqxsg+aCTJmXSLly5Ju1V3TLjvL
v4g9mw9zp/ozJWMYMRYYCvA3nrlU/P4Yl5NCOr4FPIih6IYS6Jr0TeqPqSn+e1WLRGUdrnL8CyJ3
UXhsApMXwTmmmlVKs7ON6GkUrmImwUMc3K7zMbc91fQ3oHAcEjzJODUONEPh0wjj9P/FFk41NVwh
7tiqs+aYqOp/CxRmRGWQ6m7jFz7MzOpxzhIhbN4lzokSJ9VozGciC6/A2cWZDtLdy3cfrr8OVxkN
UkzFYRHEqgWBjtBwBp86AwwdX/IC+H2B+n5LlD3sA8LActlpES450cTpff8cyUAP+C+6HXN9TW09
eLL/k435nz0iyqSy8lFhOCaYI+373Wgs+tGKhD1QhR+lXM3XtkF8euUGJq4SSqpLob1OzSMJSbZk
SUILQoLtySmBUSjpmDc1wTwxE+kU3UxI0VJ+VZ4ZH2jToS/StSQxNEsRdBcJFB30+F/pUx0JMJKO
lB0lnROIdercrixlEe47mxLQ8KX7nj/8p3sK7rOWSdQG8Y69ytedWRqTf5VeJZnPiiA6VH2RCvz7
ANuOllo+Zp4+I+Izc90H0gX/v/RoPe/K3zYX+LqowfelkH7KUBORYAwfryC7giRpJ9qHm+zovXfU
K8wW6SB7CvMKQsVoQVJOhZm+WHwRfPDkK4qqcqSqNS5TVUORvcxSXTj3CgmuZxGtM0VGA1WHIQzr
N82lJBI6cyS9wBPOirG+tV3JPr7K8t1eytxSCppgaNB8KdCU6ictOzvLaVfujd/+q03koVBTEqxn
M5/WhaYK1sPuTElLfGKfTafC3l7tRT7JBNYUJRCaCKBx9JJvOyjOUs8IrR//y5KQYOmcduPpqp7a
LOovoTJpeoxgN1Mz7/AAoHtpiltk32pyhzxP3OMVn9r/WlZRh7GfsH6lhv8IFB9KvEWUVlWol6h5
l/TjjJ09yI7FTT3hUY6C413hJ/h06Pu40orQNAGd3aKgf2LVczOZ1jl/2rdlYIvStBi0Sx+Dc7v1
x6QLbAevgWOQU/uSiA97QBjKb2nZ7GEDYqm2UeFX4+i5aqbdgIi3X5+K4rhMO5kEU8ue20R9CHpM
fKc8ADxmTOsm+jsSVMGlM5E/1hnFH2CR5xdAENY7Pqi3GRVDY8cp9C+XV94S2ZntfGVy9QtbGXJv
pEzcnpNX2TRaJ6p2YjjGmejrk+oy3lc924GzkMETKQnuGiapyEfjmzcMem5Bs5FL4Z1J2F4QLB8z
IMlozdWGFi0dKNa1ONlmosYoLQrPCDZV5YAxxRLjYLVI6LBbQLA5tumprkcDsOrPhS4uRHOT04qh
yANts6Mzw4iuOHee053Xrdp0QhNoi61lOLUcGsqgnxm0OZWxklYvbVcMz0Oeqqext400enUcTD9M
SyqdBy3e3hHLWu/KIlm7MT/u6+lwVPMzukRVkiO16OCqVJdXGd+qrr20A/SYUOpreJnIVMT5ixtt
ycI0JLm7WCeSs62o7OvfBJnuSUeNg8MFHFH+CvEgA628IdCjvMcdF87Na3PJjorjy80pdyjOhIWl
cN9g3LFoW3Vc9zjXV7nMloGrKNSceg8vd0EwQbp6IeDtVpgT3iBRWTvOlQjWHgMK1vkph3CkWRcb
MlY0fMrWDkA7mXoragH6irooSdbp/TpeUrkQ3DPSpm2NQM0HXevin6FNxLpHm0GUAcMibnD0SqnW
4FAoNwLXl+64VcVbEQVxwy+iTAJNtCRGxzePuAKb+WN9b753yWZemPmWQgcNhYgz0xTB9sgXQ/4Z
xuWX0/mXwinEW5t/e3DdSF3Tf3OhsUDVrM4hF+lIiFdx27UiJKBqxdPQa4bNF6SOlHUXUIzSQiR5
n9do9jCX52XI9c8DPy3RWc6VMqt6PCNfMZYeuKATYzkm29MaKymOMhPL4co65in5J6Rv6MbE2r5H
e/pGV2FH8QdIdqx4mcpc0UmBWHJHoUzGDLKZdT8k09wAM3+jdFJKAvOEVpeWjZ8/Qr9IKvFWk881
UplbaPxkgx3VHLz+WPBAefSDxJ9U5iw17zQRsWMPWV/vVlybwLyC4/W0PZ3ZCx3qqldlcAcRxRyv
0Uc5PtxvSWu9hmIOGZvrsNAUaKBJYJlQ6UwWtip/+frQhlVZHaKsm6LeiX3CbAZ07t2f+qBleTev
Iwe9HYJSH5ISps0uNKS+fg1IOwRvfMOyHoBakcH0Ce0NJ4IJheQUn+hcaDINv97h0SqVp/rU3Wc8
p06WDqcJOhWBrNrBDNJBcnnxeJYorSCX0PVuIiHJUu1pBoH3dLg7c8DckeXU0ukug74f40AT9cAA
LnBEfr/f+sDbLM42rHxXIHEtE1FUIs+qKHvsa2g2tOT0Bg5vg5iCItJh5lYbnmfGU6b5Yrbzzny6
K/vzSJcXevBR6VhWBmZi+CW8b2E7Hg8td7MQxCCMxvAagBbgccdCNRqoPq+kX7XA9/B0vW/v6zBP
XoOAWyB8ZYtsv5m5aQ4CxBTCk1ZgVwVYWUBQAmeMGYe3THGtvpX778y+P6T+ce2BMaQqDUOhnEOV
wdorUbbMI+lHGPFz6Tqp2/pV9LzjrKTXylbmr7GgSIuN7BhfbzEFhw7WQhUy3u0fvzhQWWBMA1cs
/wR14VAtWmMBBuDB6q4ZMYkXrClKy8dDvtsib6O9WUuuR1TYEpeWITiu/Lr8o4c1MNXjFbSvf1Cc
EpW3Kbh/GG/YDt5xmc8HpEKAPCpzkj4y8IPQ/cMsooHLcQCWneIRuMMAjZOk48PFMZ0/VQom83kq
pHA+/gGl11wRwgXTXY6RhFLhLQTLNbnDuH8xl4z8Ir6gjt2bGhZIN7BPtXV7Y1x5ckGQHAu235Av
3Iu2GsQVCRfTfbw+fq5AxxvRMZk//TSFwXXb5k0oHTxKzNt/5Hc46O5yTwSis/ieRcsIOVgTTqo7
YnRhXbAr/GI0uz0mV76BXT9dT+Ru0YXMvXOX7/gVFMlAZddfpneWMr3jJ+BrX1e6ISp5gvIkmKh1
YOQwIcRFIeRxb1422q8UfBT+8gVhWGUZ5qnbzPW4uc0+Efo9/puI9vMZdCTo6J/lO3mk2HlGtLbK
41xrH8Jvn3DysqKZyu45YJkC2aIpYo+S3nx7CxLl5ny6Qicy8Env5nsPI+ZsvVAVIMdfb63CPgNq
7Aj7WIuTAcpNXXsDAB2i+ZBkIj3NhsTAKGcaSSYLVAQBqQnBBaq86hqeJTlJ2ZG5jShTeLIqVOoc
t2r+ftc+EdkCssM9GfV19BH5jHceiFTXsz64z8EsyqpC3yJzmLFanvXRZl9qowwAf1WPmZDTZ/0o
EynKjRccMSpeM9SG2210susBgPzwAP2/gmXN8HxMc59VKBcZWyRte/0YdBBiNxY7MAHrzQUsD30g
GJ+uLiwcT31S0C0Zo9x3BJOJEEwM9PyV/Li+jH5PaogepMAqbSs9BMTlNcFMDk1sRAm7G0p2SUfw
drLEJw7LmHTnWmz+gJ4X4jo+IWAFgEuaB3yAUe5CelfoanSzbSsbKFahCHXLnCu/8esxdMGsOVx5
+gcJH2T6qzKyMHfUTpzFw3YclmbG9UDhLNSSYa+2otCt2gB5PSu64XjXfqNetsqHtYS2+KlriU0K
hgDq4kF5K9qTYW3s6CRBP9W7Ya/dMi3+OQdrCG14Y5U32dfwWZzw6iRgOjD4oeju88T/pL7pzRsc
9Z2r5utQhQ7FrqCS0gJ/IdDADj0JBJP8+TZb/XwfoWkyt40kdY3+pRQujNTu1uhZPE1eqX0Kf9zt
f8pq41NYmdkonb1o/4eWglOE+2B8V9x3PnKQpbvABJun/yzCW+IaEvxecVrnDpYXG5qvVO587aYk
CBp4G7LRXWAxBFmAtUqfrlFqDnZSUx+pFktKvqu4A51UnZed+R0RnpK5mKv0PNGOfPEqz3qfva7G
JzWF4OXAHl/i/Xi88XhgB6+IQFq/cYD7B8gbwwbnp9ki9kFD2HjXZHygMGwmuBeDdtaayZIsZmN8
YeuHLR9qxPsXEbCpqMryZbVojrqlOU00H2MGlp7WMRHgmJu5K1N0fZ/HD36MageOAxvjYhiDGSaB
K00H3xyBk5cB8MKzraYLmx7vTdfHLR4B5Nh4pZvjeLAsE2A2yk8G/Lk8yO975nfPynleBbyj7X8H
JneFrlZyWumazPBaTMl7PVKitsqsVCgHi6wXV1N6CfLGNyxktXTrRTG2mualaZbE+FDLq5Nzqjtq
+P0if5mrCW7q7Saqws3p+iImVx2+Vh5g+EVBmXfrxDFZJkBeBzCMixVtRsv/9bcQrGvNm14xTce/
OhOZTNc4UYTXVfePX1fvcmBtPH2VPkN/Gb6/ldAFG9AfnXTBFhAxEY5PLMV81uS5idG+3Qhs4O0C
cElfr3pdeaJXytWNqAXz5eACNUX7g2HKTqsvHK++9Gf40py3CEpZntEN6oE5raztTIRlY/tJdfpJ
p2bIIBhH2s6HdhonqqCW5hIOGMpIpxQT+fSPkDiVsr2XXdaSyvthgnkZErMom+3j3bdO1REcQ9Vf
MtTFaIx6jo/t7auVIhF7AJ9kf4PxpssnU1TR2KjmKkwtN0Izf8omOyj4/fQXSHdt3Kg6xfQ6wLV/
jHl6zGR9EzvDyCySGRim0epTRMCtCnx/ybSiFyt3cjP/A33Ab4bwuiEtRlAt8N96FCSZrba3ZWA4
LCgmcBjkwKj15R/ikLlHxUq+w6lt4mJ44BA4jMOSZ9sZbEyYpRsHSTfcPsl9H4YTdJnfqeb7CUEl
sfCyFe0iWkC0CGfG9FWLqXSPEgQnkOuytvaggCJ5AkwbuBY53DNZdD16l8GjAmyziPetGmnBulje
mGLgknoNrAQsoCxVDwBwTQJqBnl2gtgeS92F3Lcy+4ySk9mB/hy6eVQb8/zdGJR/wKL/ykO/Vhz2
N5hx/bADY4Qztju6g69mYA0Md1wvoabiGR9CEa3y+kKfQnTw6hy9y7ieIq7/uzcA7AFIGTmPzw9M
LG7yTVfKWUf4gDFJTYsrYjcI9N2oyroySarRKGT3wCpPSJzVBu3esDfZJzzGfnrI+SKcIFEW7DGN
8vG8V9z/ihbR6HhJEuWUEUor46mIQwVwehZ80G8iJgpDlcRzjF2t4PHUydoHEWoczxhhKWCZoDb2
xS2UQ2BDRNM0iwNBeA6aVDHGIxLK93INSY31lBJ2qpuany5UYOGr2Vk6zkCz6NPjkVahbTTMNMfg
ckpQcwN7HWJdY0S/WEiAbirUYvVnwgWDg/YsbyxycJatRCWaIdGtD+z0NlZA/O59HqAsSiQyFWJX
e1PZWa15mmv6C8NsgfbAciqWLH/Yf4/9GIDBrnHdFKAZwKPtufqlQBetctHB8q1W0Uh0KXp2nVwX
+b4xtPdXuNdp+dCVGXkhW9mtRuInGVml79txNFrsCkb8Qm8ibyOQ2pxojTR+bZt6PwOZt+A5yPkl
o/o5izKNcuLQCHERNidLy6/Ihvdo9260qKdYdwiQr2wksTtYlqXuP2KMXF9C+wJZCvJZq/u1rvAv
ZG6WGfCMnqwMI2D96XSz11PODAcLmx/NFGD2PGdGfS0fnEA2O6H1YfvcXGOFLzoW+WBEhJwiOkAn
S8ZJbK3EDNJ6JOCmG99frNHikrmII8FZz/lrGRxKl5i7rrV1DJl2VscW7V4Tk930X0u7+izayC+a
ihmK+ktclJ/h3/PfxU1gsTleCCNLYPMG1JRG+p6+kVhagSZfGQI6BqHBmTd2IyFhiC7T/tT75OZN
OJszEKlCFK4ep6a8YE3cdAnKmXVBfrE1TCpXZcc1Z8mvj5ADhn/JBtEtCrNU/VyvkQnLXwT7KCkK
DbF+peHZDD4np55B6zOc57ldhTxO1W2qD3eT7LB5vPOVSIIYDL/oF5067Gnis68jWz8Bhixx6DOh
1eIcNrY3VITRX5tZiC97FcWGn1hl8nZemzCUcLV3ssSqkN+3jvFycU4XVMEOXn8augRn4uMHMqxo
adMuNr4VLOg4CwNnCU+cccJas0ZEnYthmYV7EhE+TwVHRbs76biBoNTr0a+YnLYcF30nay85MkhV
GSSA3sEaryWW4ZGnrEA6EReTylTI1rPwhsQiA0khmpAW1nal1BKle0k7ii19NeP4Y8v4lzUiY0zE
D9Gr20fl0pVdr5xacWETtfhlHNUoi5KlZree6jrs2gToK8VCHqvm+1GozhmBYhfeDYmDTVOkODvl
rRST5YVFvRtJkhsW1T4BazF45vwkTiYpWMK4OcAxol6+ijwKUn+beouS80hhcqHoBcBSc3nslwgB
naMpH77Akgq4YDoAVL6Tz6Ioj9aUIt4ZDdcMiPI/d2x30oJ26NLSSEYajIjIK3VvWEnptY4S43Lk
puu/SmdVuEGijVNxL2jG6tL0a8DSVUTN53Sa/RWrU8umaCl1aewVtO3z3yHJuqtwM3RHiEHkRpgf
v0O+eEg5VNUhKNCNbDR/stZJJO5RZ26+I2Ld71+kjwn0jLff7AxZiZSs6Si/awHMoSWwSznkoAHi
xxmiQNgA9K0F4Rg/rB6eiRCYsx7yAXJ1lEI2HSBa9QLsHsiUG89GVrCym/631a8o8a8T7y6yp5Pi
kLR7bIta9HMZHVSpjx/Cm/KDTsOevgsw720JVzUSLPxq/aUFKbzRvCZdfOjcj8OMCK+XYT8xeoDa
YAX09ku4vy/9Yzi92TXODArfKhrq8d/mlJheyKdyQbqohOUGjxWgZwbaDJkcL8kSQulXC1FUygGU
r1keP9yaKpLipHGHPNZPMagWO5GJdmjZUli6GYsB6Fe1/A8iq9S5oFdYjzc1hrQqh3j08p4yn1lG
/J5YscLxTeQiF7UpZ+2A5+cA9nEhKeLmbYjRLPqkI2zgO4LtGwFmDwtaO4jYVZT0cewGZ2G3JGXC
NSWAfFxyQq9hr1DY0xxI8Mj+qFFlzLuDtpVvaI4zY3jPW+mD5oBjUBjNPLXw86ogJJDh+kk1m+qR
d+qLMruaeATRIQaKpPYac8UYY7lMUac9+QEEj6oGvnu7W67r1Bc5u+7hvAibW8YMT+b5uueWkTy6
vsQJ3g7R1XVzXq2/FTKoVO1AVuU/ZvlRa4Hwho0TWZA3DBgq3Ze3S6DiH5qpxLn4XFQCkpH5S3Bu
RyaATj4gu6MUchf//kklF5WhtmYzu2vB9eOKklBoQmG2taRN/kR2BnGAZoBhECcd513rDJ8b9Mly
QZlfCJ7acOxokca25stOvfDkFuTZ3MzgvDfgPKoz51EdPqU9Ybxg212O1E5FkaUR/YEKaYFNgjrB
2IHyfkM2L984NaBkU+gO/V8HDP1/U3lI/5LH0qYWrL8m1nMlnoFZOAI9BoiNZoWB11dsZagPzQ+h
P8fFn+7nQ+gjwD8zMqOfGQtfOAoXEO5n7v0F3uXc3QqWP5Z+P5k1JLJXvphYXCmRtitV2HjGAYAJ
aVIcETJY1jWW1ScJiINio640tfRPIkPKN4KN+L111MUUEKYkZRD9EgowP1MUJOeasm+zFj9yvfOw
wDZEQlD9rbVHywTkd3VpgGOZl9xk9/xf3u+LKcS6/BexPS24GhmCQYljIC1LRU2ioSolT3pqHN58
xkFaisOyXBMakJ6mFKkvSyN64dOdeW/DGMopNV9ajPV8BsynVBrBHgq7reVhv225aSOSPIRFzP33
GllONFUndVX2INiOU1gSn6vsT+y0UTmtzQLdLBLNf+4GU30AS2RUcPYmgLbezZyl3WZe9iLbyy72
uIFb0FOfsRckMnTYi7n44bczuUpjH3sQRzlENJzhGr8sp8BArUtpniR/hvjhwtRntxsGAwxy2DvD
luJW+hT9RSD0Ox7vBWT0kK7Jgtf4yLzZsHkMKnZMZ3+dyII9Ks2lfW8LhMIVB1kVoK3dpLbzslq7
jKxbFTSSZcxzJ1B/vryWQ/pQQ92d631YI2CsEK189XwAleM3a+jnrDY8rSiN9bUyeKAmDs5RwEXq
syOn7RRMjPZhlXA1l7iBEWtHqe6Qm2Y3oUT/qNR61GcwCdIosLwf8tviOcJR+m6GWlBBDKEkAhic
AmCL805rrbO2ZQaSCXCWzTiR5aVbMTgP+xeTXU1GcGE6KDZZtKXwbY6qSBmb2BuKl4DWzFMpqdYt
3XYvFGoz4Wz0pPMRmq8VZPFWqtFHGhlyhdYsHx06VHYF+yCQNAUw+FHpYyT8rBRjgUm8bs40e1hS
kZC2ZAwPrtT4SiayCtv9DzSOmG0sUISxakwodT59Y/pKEEecPgzTZtMWbz3sZ2tMQYRwaH5Rx598
npkzaVzLt38GoERHz/9BoX14feB68wPj0ufqo4OKNiN2O0ucA/yEEjxc2I50SsqRVBbj2E/QEv0d
6p44wlZW3Ph7Uo2OiOYC8vgJ5eUubMfyNIGY8wB81ExwiDyRnxQ5FAbPt9Khaxey0HDBYpeQe2Et
X/yBBq7sfHE0+ccmu/q95vvlr4y/1xGfNUKjt7BFTOAuEJoLwGJLCR9+b8yCkSnt4UmZKpDQI9d8
PodEP9n3u31tYyyhFvo7/de75F08p3REm49vnkgSRXNOyWK9H/bl/nxGLk7MWML2j29caVo8BliH
mLWCezSHnmNDmT4LHqpS7N7T8+N/eAipTKNG6vtCNa/9EmYkL3n+V/YdYjV8UWL1SoNrW7HehorC
uWue9Lr93BIp+NiZedqjo+4JUK6RRm5Q++RSO3v+l3u9pAe2uwx+YOoyj4JQqpVc5vi8dqulC3Zz
eZhnL+zwmOlYO8Zc2tmp7TFxGe5x8VQYIXkJ6g6LMNO0sbR2vTyuPhyftsOfm13mfd+/82o5ME2O
pxmlhVosOT0IL8g2ayQaBNFTV39/aw5+1ZhI7hblAnBGlAENVIteSPKdDmltZjdwMCIkrIiGkssb
sa4G8XGxfr1issyFemaeJjYw75hWNheKn0fLc64LEtGofjDj9/ghL3BId1UKIntrhLtt4JceMolV
5OdNa3+LJkN6/bzhV728+mvYW5I/fOVLerQ6AVHeo4lWfV0p5L0981+fKTSWalRPl1x8zqdj1fm9
WQRmAFledgGpz+XSUiF1id/Vy5PWByFXUe1Pawrazu73dPf8xhoA7PCfKIrdLqpKPgcfx24BJEaw
7awBfSUZElpzSQXsd05ZSM4MYX1bP9dRzIy9ZWOdVhzzQqRYrK54++ohb0gg30y78vXl/u2N8B68
RlFl5jF/5gb0khIOWadkZefpXuum1RrnW6EpK92eaz7PhcAUQb1Let3UecM6x0o4SMGtegPopXxy
DrAs972TUaqwnK8yUZJdhTX7OfaFd84PA1Vh+MXDfb4flLgJQm5lpNpZUP9iJkTnlnskdg5Hhlbl
CBHdsa5XO/v5GCKhGr2wb2dmZW03/o7yVadMt8jEvquIamYY5Gk51KUGlHFfMpcIa2PZPIGUckoh
kyf82xb0hgi9SJP8yrSMyY9hJBan6JzVnr84j0cYkwYOvNolaLLOi/2iRkNO9nKeQa6rt+J5JxGA
PzkYu8LbO7LC8ZhmIzvWKQCUdkHAzTo5HyTIgcl3/QWO+CeTlqCtL2/xmYBrmNW8uphms6tnXwYk
a42WsNeKjyGWSjuycS1O6J6gIMjTfFV1ssc2BRX7ZAkWYqNbiNOGAkE3CumlXD8laBt21x1db5lH
kNj/w5T3vtiVDNHy1vMYmnUlGTDIIBWPDiGbxV+YgXAB6veTJ8yUqgS5tfjGlpg7Y6bu3p8p9k5A
XSnA13YONBjYlfu6Mc9aXT118W3IFZKoPVGoQOufz8YkR1wU+qXdhnH72s2e5T0ifnBaAr2sTbH1
/Yb7geiUEF6dPU4yJrfHIadFPEFnVu8PA6Uuo4IeIr+U1z1q9QIELETwxvR8GA/q17/l2vjkfaM0
/dwy3e2XTyF3nsKlmuujzLtPFNHif6buMLmddT1vq4mJVYx9e4hzqXI/ULH/wln/Adt1WYZrxA3D
PSIQ7OTqjRNb4VkvS7y8wPIjD+uh2XqMveKqGhp6WVxKsLAiRivcBRZlgam8uvREooNFYpw4tI79
MCWB94hdhMPgplVo72raSJ+K7Dpc0Fi5jG53rbtur4KWLjeFseQLsojSv61yhK3fVkYeSY1yGYf2
Ys6BZsb/FrE8cAjr4K9NC7T/E+eDIjuStd0PlTXNv6606yvdEsG86KOcZh/CXhAvM4/J/2Igu/cX
wsh5ICW0QcimXn3A/IpeP1lww3lwBKQjp5bBc9SztVjEWM01yO1GcRd34tp0yrPH9hYeElhGuIgh
W4rin1vsiOJt9bv/DnAowTWyODt4NqUl8M8yX5bqXwAyvAGOca+Aiym+eLVLBdRNAFkrs8qb4Bdc
frIjKOf2YEhGRixfizBLtinpeplUW89Nh3QBZn56vP+Xbm1I+KoKxAcjjDlO9TBbiTubxpSpIM1u
wLYS17O3FfplsytZkrqHkziI7abn1oF5PmUU1p5DwTxUMK3LgeY0GF6Kg4QufupWdiNPkYnMTXSX
Baq0E5tIanaXNFMWDAtlN9YU5Ye/jaAiVHcsiZb+q9IwKRLtRe3gSaIftUGUFNAPySBbnZtv2cJk
v843catn3gGKivKMsDwydO4Z1E85oW1B/HWN8AEVeBduDdbXlmjmYlgDQl37TzN9rUly3+tesMBB
XA2KbY+kGr8VU1Xyk0nU3tt0+hXp3NaMneE8AsJ37r+iMxG2lVdxJctTyMmBjQQhAFmWk1agqFmz
QpcSQzysJbTAja9oVR9fqjAhoPOwqplMNVeuJXxyKvmyX0brpJecj1WoEW4VLq6HHGUlRz5vYP0T
vswjMkZaQYNAQ67/EnDvpR64pSUHHQ/gV5DwfvM3RzgyhCKuNOezcgJsMeoJX/M245em7MDn5rHO
PVUVkMFhDJW/icTcqs76HHFRM3N2pCTnggL6akWHxk6/POI5qGCpu21fwxjUgsHqxijLtOzfjTbg
+FOMD7e4EXPn6BXrsxroJv/hoZx02Z0mG6VGeBuxktt4pInMmw7O9z+yZpVnxxkUa2AKGVoycA5o
SR886aT0aWLvVGZOEkAb/rIiIPJ0Rjc8sEYVgUvhE5P2MgrJv+TKktsX/jY35NNYZXlEH/8s4BDU
GiGANvwISCZbQwE1Rnsiyi6glWRX9mA6umYjuh7wKWLneLnIxFKxc8xMJUY0GEL+uujLLCFbZ35/
A4L9Pkjl6Nwyh6cAkzlA3I0v8gd6YjE77mxZ0VQ6WTkRzbZDmcWJmDa8DEoT7e4jCRxdIdU76dFq
MssIncUPQdnPbg9hDIeIl0nq/LXj10hD7t1ywpd1b4l14vuEDzTUjnpYkTTBZQ3Vdd6Zty7jQfme
U9/d8Xcr/vnX6xFcciq6l2QQyJmMKVl5uItQxft3nEWlTGJTHzTvox4EyZy9v8vQYEiAj4jASC4D
nUB7E6ncVLcpLjIz7F/O/wrTrsi+EN7N6M1OKqH8lULAY6pYjpNSSMhddp7TToTPQJ4PLmt7U+9J
4HFrpkVtyGmAWwAzS7U1oK2N5W3KQxdgUVz3Q9xuPfmm6thFMQR1HBqm9nm7/K6QGvrS79Co0nZ2
DSUfuDKuMP9qUi+CuaF5H966BSpuf2H99yJhEw0WFYCxd5/Q4qEVnt5DKSO85SSfXOqSZC+QnyHb
0vZUGkVHnx6D+oLxNOi97AVTaRCiU3XGywCiYqMckty9HlmIO4XWH/5g/cc6aIUltrImBilUoq3t
5o9FffNB6ltKpFQrEaejrFTS818vR2HPxz6ew+G0VJWB5N3FezLukXLKNJNrCkUZ1Ob6JxXXGCG/
giH75n4fW1TX9zolKoWDGMJUCc2im6Uo+hbOFIi78X5jC3tIxJNMEAW6o8BntwO48DjfpIciEBtl
iGvSIUYI8AgMSDLu1yfnzAxzSo6Xg6ikAHIYx4tu+OruTjZ50+LokF6e33Bidem7vn2x2lDMeITy
mQFnXDt9Aez7/Les8dtRsFkrRXNE2gLGzgQM2rvBjtFJISpYLFKK/jr66br7AxC+fWUK2o7cdty7
4nEUSywVRB2LKSv9B4goobvJFPNMFWY1yOK8M7UfjuSm0iCOZBVaaGkn7Y7ZbBmdTEejT0i4c5wQ
QhtbBClST7Rp5CckKvUxUCnRgSw0olV5Dgfn3vWTQOxlaDWWSP5rc0vrZwXvM+0oQvbdPhNw3B92
yroq312AuNLrpKdT+OEuzcjTsN7VFyypWg0CIal7HZqf8lleUd4iewea4BVKwivZC3p/cJiaC1e9
KVMoja5NUDqf242DwM+SWytmd/KMO4BH2T6sNToZwao7KXOxCYUq93Kq2WiF71ptmp0Savnu/35o
eDoaEn5ie4itXnuxutD4SHiXj49i0rl/L6jLH8qPPr+XeFNOvnjU49u8Kxfk9u4bjTxB9O4Ke+sg
9wxvS9sVAiltw6fZWfM9oBsCwPzyKweuiydv8wFBUHFs7rpxuNiKpy3r0jtduGgiq+jSJ88/gv/j
JmwZNpZ6+LtJT/Iha/snbTDKXvVEtDi5+y5I57N9sqsQjaz/E1vNh3I7FqT9RpVYYGroQA9VTAjn
utdbqBvhNjzBzrWzQxmw6RFGcTwdLwVMAtHua5D/Ew43bp2dea5klCvOCX0RF626z6VYQxOWEMdj
6gxxrQHlRiNurJ4rNkzAdQGlZOhvcYTibrHY+fUxdIL4dNqqR/GX4//P/AEQXV3moiuYmNNrcbDv
6bo+c8Y+Bgz5yN+WvLfopTBsjutEzaO5gndJO6if7XI38hazSc9riszwqEy35eiv0fS8ZNIDDDzf
ye+YnTWdPjmIeMN0EQ8dMVJdVtqI3kF8PoqkmovsJUM1eLxQflKOAJXFa5wx7VoKn96lR+h4Mqin
PCqbpWSxJMIbTjqytrT2sEj7uDFewjTsR6s5tEfkJdrGyLfaK1qcv0OCY0XNb1qpH1frF7U3VxvR
oL1x/S/0XZu1VEQgc6q8gNfOJ2pkftEtdAyv/e/9kgXZMPi6a7alLQgk7yMjAwI1RmmgLvo25hia
+i0awSL87fIL2w4Vn/NcSOh1sQAgz44Kx7IMNDk0zJSxyoGwRCKgUF/jtbanqpdvANWXgfAjkK6H
C83F/QaJGoeAsfgyGneUdSwXkHRd6cdT5OPH/hZfGMkzMls3AVfUwDzSrXm6yi0QYdDByxP2OlGr
6z3hZq0OWGPWQ/yQcP890y/X6JL9aROJlI8bNAIrsfHbqlg1jtacXm0msW1lBekPrtRHE5lZ5+uW
6HMutlb4Mjb5DnWzrEGVngUewHQ4JjWFYSOXZxAH9U39MTEyzaX5ZziujeIHGH1ylduckuePve+u
X5gTExd8OwqfBpqqUALkmbsO8GsLcRHPTTfpETht922mhV0eJHe1HVgtGN2kjJ+ke1Ma8wbMuiMW
ksXX739xr4epx1Z6ctRqh3sUR1OMvQHahwQ7PhpjaeJDwMSb8zJ+jYfKovkPlbm3ZoWSdH45xWZf
0BXXuk6Ar9MWx7Ndtr2lvrONMmTl80h8sgBiSKf7kjfqDKIU/iQQ7rrFOXILfD+caAjcKrCaNUFN
7ObQhMVK9cJkbGa+qMfeAeg6tXNzIQMoRcL7vTaTDJF4GfzO7S557RVaceBmSyOM7vjFpywVS5kK
j+h9ffpCCsyvmOIFCXLq8q6hs0I8BtTQPQBBOllOYqrft93MCGyHdvu71NivRTzXeVigTXPXy+ZO
s1alHNsJEYN2pxnLrTCf/K5IRbLnOYu0of6YvXV5FHxkfiV9r2O4iWEeuNHuGuu5araSr5sUtiLw
ok2e17O/BPJaKk9jjGH+29K5LpmLG862Icu8sHd1y42WOMidz4oDId18JakRHzF9GiRXsnjnJnKx
6vUFuKFcb5iu1Xg7atjM3kOCDlA0HM5DxqMi3PBH5MLofBFOZJRuudXNzgMVI+j1Hc2SgqOo6ggK
VYk98qCC/K/hgaptQ9tFoIVjIj+MlWaLdsgBphB6T+KHPP84nmWoBKxPQMMFIFhbe606/qdtGgtz
TU7fA+jvFTdb9mJLDXKWV4TUa0Gj3oRtDAuNzT1ePf45yOiSWZqYKMxwvV2QHZoUHa0wTyu6JYOw
jXXJszdTy9C05/henhEkJvjhqxJfZryFBYwU65QUtfzYLA2MqQ9E1z/JYajtrW6sy/30TBLlMT+E
9ggt8TaaIRSz6DAuAaGwCwM1ZJoHGy/4oSpBbhcwFnd5vF+VZcTGnvVrf77rdGToKBKvb2lyLC9d
YZf8+VYB7ttlaoGCqwyQ+Ie92fvB9So1iDWLnzLXkrImlvybeJSiAN3rVfdSZpwCP8TvyO1IVli+
ur8Vjk/S1lAHV5AG70mSOb0DnSfX+UXuZQWI5RcgmxBoQrtugvrRIDHFFQYhhLn+ZHpyXDjT0VUL
TdyU9jlDGTNMtUmwXb9F2RX5GHDngDcFquotKjW7jJJhOm7xviIMiYPLbDj5J9cdFSDQ4FxN21W6
J753goFdyClnKxjq7NHB1N1ytdPMD4WzQ/97OaY/H+gMv8IK5sPhjb1vDK8vFKtaX8yvFSUHjBkk
gWLMAUWHpJRs501Wpx2aglYzeEBghijTizrgaMaCO+ekY6mYktvO/7Pk/lfK4DEzJrZBN+QKd8oT
NMFDGsNZMCj3xT2DFtW7j2dyLRkGD12wWfZ88LYxkyMDJbHfnFbubBViepb/F8f/0M6ACsJmImkP
qsfKjXix+8kiW9B+lSQX6wYJPZBNurjBp0BFO/toIbmzoPAQpWKq5n6yolqmNHorTdC/+2LKPYLS
lvUIm4tqxGx2CJNHiVDOYN9wjao+qeXyqfohUCFA+mx3jQl5sn6BFen1UfNe8B9qd4glIF3vqSJy
E6LGzkcmTavqpB5DsxsrYjmxOdYci411JmWQHrIahz4RKVWnk4yNbSux1brD8bvrKvPl4tOqHQDB
sxPT5wOVsUeuOinD3ypD3pX+fM62xBvbD0mgS6975NvNuGKZ5Ol2h7vx/x987+qnJgoB+B6J7p/g
hmUomIWKkDbbgolLVAodtCI/AA4uCP8vMPbmJ33I/+7gjd7FppYp4Uw5uS3b1XZYVFaK2WooAj4h
t5HbC8SmEnz4l8M2NBOjZ9de1wUKGuVX2OzHoawn2QRdrPZ/VzLEwtJ1D0chIeQqAOlzd4WC5RFh
D0MRJ458wU4TO41kcvgXdI2PU+eThSad97gpbDJxmpxuje1EcVOQ2VaFHJieBJ/cNP7GIsIeWF4y
Dv/53MmmpP7BWK3HSYUg/4sJXwiEfZBn3KzHUZyoStbEAs8DSUv3fv59U38MKX6qHq12F//2AWD4
9G437GsJc5UAVHobIhDZiaMwrk0znEijqsF/MNQmRDgoppzoLxepKDk5/dx7jsHT/04+kbaydSFu
P1bSmoAvlYX9E5TYVTM/UKmIg8TmAvqypbG4aRqIE1PBHyBtjCzIbmkYhfX11zdND8kCr6VHbdje
cSov4QCY/N32XAN1NWS0SBmXeHOafO2/vw+tSgWjR4a7VWzS0Oms8emiH9pvQFQxhldak8hHGZZY
BRDO8wO9rOZ4o15z3OPNV5oRf5ZDBnP1Y0/N7pmKD6SZZCaiXqE1KZM3IGmyXXykAHqYhZYYw/AW
vx2mJKmK2o6iKJz0d6Zz0QiPmo8V/4NKeN9Jm8oxi2Drl/mnsLB1fUFWH0quARNxl7lNwLsPbiP3
XwHb6OLopSStGZ47ceG9zfKojLWA6jFMJaJ+7BJutpwz0jyPCCvIySEdKHNGIdlWHJuryHql9O9P
infZ+URtUJLsT8OT3jLJyJZhOmd3Y5f0z78KFNSdZ3j9ND/OqhcEPFQpq0L1nJDFQ02lknQ0EFH9
Kz2eT08/PgDOiAvyiyjQT8S2rJgDAtiZPLGp7XHo+LrUBUr8kIu8ja2DZ3Rm1Yr7vb9mPPw/hn/H
nnzrU37U6PwP2Wk2oUwh3RnWbKGLykKGbROBPNR3uME0vZp/V1Uzyeb49KqYoYwmC1qb0/G8WGxj
YkpvxAJl3oMWq7TDR95K3xns8JoeNBFDOmPq86+oNJ3xEnY+E7i2p15XCQI6ewAiP+M95YUVjJn1
DEaJj5FL93XD2ox+K8qOOA1HrN+1pn7GPumKDtqS/zIXqFSGBNf8AMWpBabpEFvqZkRrRAcGWFrf
80hEONdQ32rgT7zAWxAQ/dAbRlbWlR3fnAGW8FB6M2bkRua3UjINZrOT5DobMQ/XUc2g3WSh6Jzl
3vAzsCEWpGXAPdvNQ27YjK0PAk2N2dwaGn1Q3nuo4uhmhrM8/4OB6jfkmt7l6QMD9+6fjv68PhZj
XT9K29jEXt4pgDOWRppnBGPimUBndnpobzDtoimmuWEhPDpfv3wpBoubyXlXxUALzaGsbm0mV/Q7
Ta72CBvEnWQxOEVmhDPRFMwt4pMCu1jhqeEdyU+ZiIJAxRBQKAEGLdjDEA17YpJq3xH65uvzCXwd
4N/KPIBuF6DobikdQOrlxfV+Rj4ujb3o6mg8J3FAUED2Q4iHMCWfjKCeO9h5r1LTmeEJmY9ZiXJG
YCOvjWeSu7+GahZuZxPGeVMhzxX1HtaMgUE3YSrQEj4ZeXb7OGpTLaiezPMupleNQj6rjTVuyHv8
qxZXABc/3gXG1f9HUy5KErJ+uDCQlEDTr0l5pj0Hesm0e+T2JzF7224/lvd8+thb6t0iyPssooXV
R4xlxoFfkPfIIJzhco7AhES5IKrshkjspAv6X+rIEvYfWWT0ZSzwYyyF+qpGyrjF0TYRvlhh9Xbr
YR4c+0hXe7C9qWiPbzbkEMu5JO8219EVkQy43ENOB2FYHeT1Baeb6GHAw2DEui/dyU9wWc4DYjBZ
O1B3m/zKljymr6169Sq17Xzwhnav7idQblnyyDzNFMcu+uMHhesLGZmXuPkT6vHJTRYeAdoYaWUF
90T3/64OeD0Zji8xR+TDZ+XF7aBRaIKfJTxooKbLwtInBVst+U1y/qlqLRvVankfLtKRSUjazBgJ
5K9SBRS4/Dxdz7kEdzBwmOGAKDGz0KqIQaq1Ba+f1fdWoyqj92iuPxILTnNuSQr5w0Coxo0K7WjQ
N0+n1l1hYU82yacml6Szsy1j0tPiCSD5yhk3ND0lanN8v+PQNFESnBRCkXoTF+X2nDwkNncb854z
CQ9y5EN4o1usrEbvzCyLJIf5oFjvOVEwH/OIsCgr0JM7zEmdfWpGzRMpYrljx/01DfDhvd+qikyJ
1PnkCxWHA324bjo/QAG7CZyYK+Oohzx0A/jvrRU4FtERKkFoCZY8IkZ1nnLuAPVs2JwZ3fSuEwoa
attwpnClj1MV6kTESlwOZiq8UIF87cOPadberjaKhn7ktQs0r4DerWaTRrgQPutOE2Z3SgpB0iYZ
Ups4Rj16T/eZP41HjPPD0Nb/ZmcpL50ItKxu6CzlWmiooZBLrLcFbvfRwOwUijR9KPOIliOyWSlV
Wr52QuHgCqiXwD52SLaKPBN+1tWv1VUeLE5ClRvK2JNWT8iBJwhtq1KxBXwy0liy57kFZKqQojqn
VFSvM2v1jLaPitvLRg0f+YBMGURsKo3lkkKmIO4nHA29v8bTxaB1Wfm88/UmnDPCr583hQ+FvCJD
Qwa7QVUYXJ42vOCVv3Vix/bDX0Qfhwkcl/h3vZdhrnyf4UUsyOwfo4kag6x8DZcg32l5RfAAejWr
1CeMvUpSYzvJUEA22g4qKnxynUhPEJxB2XG6WG2IoF74r4Hwjjk3c8Eu1D5NC7UoC+cLchwgtula
qN2jXjrqsS3stiGPi9k7SX10rHH2VNe0eVOFCCgYVfI4I/MdPCyuptDwOJbei1l6aVjAzlcFe4sV
njlvXG/WC4Jm07hkbEvMYGxE7Mu5EghOCKZl17cpaQIeNra1csSv1v3oc9AXLazoGDW268wIydVE
iyVp+Lk0WH9Jzjry6Jvhc+EJZ0Vq3lb014ci+qTMLeJPHTobDUc8PAOj5YtIjzzk2vJ3SNbe8cFU
T5rB/kadKAMhnwXzxZPdZc7oGJ3EpsWJBUjIY95+V63sJyDWR72WeOI18Le9NMaboDzxxAZmsoNI
2TawmdisUqGQQCcoeayEbL8zA6sJNbhrpSOxtCfbm/C13XVY0yBMte/SDJusGPbomHCR7ottD4xB
XikaVLAR+gnqsppv5MwlB/i2hdLjidFC/6rQkpnkYbdBSfjYsmADyXS3YV82olAGDR+v/iJDXTOI
q+aC4GWjRdictOLKSXkYfSgf65/D+J1rNf4lnKvjTuEMTIzWP12KAs15h8w2cr+ztgn3thVAo3lw
rra/BNH1G/zFRNFsX+YbRqf9wNonNboYylA8Ksq+P/mZl9OwnIPyCA30NYwfMVru69PAPDUtAARO
XE9ok4tIKH5nkpiW9IL2uwyO8dcmFNrw4Jx0GeokpsoQAKoj5DaFUWUSP+xVcMWIxHH0y92Umgr5
PMRUHtP2XJI9fARZ8i9YZntvt//VZZE+azLHKkGRlGCud2jtQiByl8lr+dfMG4uYINlG1JdTVqNe
Xk7uXBf9YTBVWA/elFNt7Gn6XKNXd64rLsYY9fHw6Sn06Fub+twtTNOpzGHo/ZRo3TGhdglC/aG+
Wx8VwjRi/7fvCKeccXzHqwg9TJDDraRkM+rzqYyd9xBJzoqI9rHRYZtnZP3aezBH3rcIVgKimVl/
HfXl692k7oZdr1pmRHr5mZkfu5Rx0aU0QmHe9TZgjEV97+e9ABz3p0YEEXYB2nIKyY9bLXf6xewo
dn2JlIm75nJDvZ5BZ8IXQZjmwpwf6PFZKvpu5fxI0GuH9ZxE1lVBCPiRgUscKfA62eUWGg4PW40n
vNjM6LGhMl5ZRxf/9geuFk/obVfM1ar7bF4ztAhp8pNcNKcljIjaanAlYEjS0B2cgQnBGwKVHq7i
V+DS1zmpvRBSSZBsx4qzryXMXgGhhPuJdZLwX8nYKOz7/mwXoDwHLjdBlDw8b2kQ2s++ZzPqq2Wt
uKfR3FEuIDXWM2x2OtThBkcuuyc+3kQj3R9c5Ij0axU8Hzt4TiwFX0IfMtJiatCwcdZDI9fcGyJk
Leq5DzXZqjUrU95o8Qtgb2AklXgN+MKjolKTmrfUc+nKvBICxL1K1dQ14ctixJg5pJldkrPPaGdl
UQJ5aogSKe/hqR0YjPDsutpAJyyx8RV0kKJ2Y3GVEhL0iat4agWbRZh+4tMmETplSCj7eate8QcB
14gembX/srOoq1gIjfmORxLsB4btg7sJRHWcMRwVUTrBQE4+pTU+R72PVgWbc6bGvMIMA5Fl9/+f
GU0PLeO4/VT1RoiJvRbe2SZkQTK9NQ5Qh5MPi0dWQtQANs5RmKPdTJyUVdlg5IGwqt6k6PT4d6Ph
InYl79T+zrliZ6V3gq+7iKDYgOgtp/6EIf+WvPxflVrmgZCS4NnIr4xoFCUFij6eyEz3rMAtwoxI
7qbyOpyM5ANP7Y2CyX5rNFmWA/trDrF0pxGE+he3VXyRaw9YOStFMmUOGx/mUfxYlapP4n+q8Ehr
1dW7VnSfp2baecVOvOW2AnodYi91AwhviAw0E68cZnjz2qHqTmIILLLl+cWCbzZ4xLxi6WS95uiy
SijZqJC6ivofSd54VJBLmXsjYKDVs9DnK4i7FFl+nzHsGn72C4SeirWfYIojKG4dCuc10xrb512q
GKJlhqcIzmclbxUqW0RxFsMR0hh4ZGWOQCiyZJFyjRwqB6e9qOZG780kWaLf5adcostjm1+8i60B
NqYdaPw+zUjE9xlI8f3Su//qIjNpgvo6SRwg36hhUPRKClOUVVTn4LGQ1Z9qfvnUSnHAaeDN8Gwq
l2dmLXGjX0ATD1s01XQ2MGtCQmjQnLdTNOII5YxCJYOKl8QRGurZI37cDoktBTAInBlIzBIr3Js/
Eh6SrapZRZAPAc5bHSTiyLU2iRqIMHEi2/M2XE406rNffnNHcHSjnrmAZnPh43isl++61+eOaMa0
cKgq760mu0/5ykn5Y532waDSVu39H0HRGWIFKDxf0x9GySH9fQTV2Co58xvaxuHRyFF1mRvnWVVF
QB5DVJQdcSTHAOZCUNmSuTmDmHzyY27GIBOqt2VrDOKoUQWWrAFcLGckK5LjGIK2NOsiGUQVvx8i
cLERy2nszhvlwTFTWiOzXc4twY0z4pDMvm6MxJBEPOMUbEYKw2XZo35VQ0Az6dylHt4C6lf6OZw9
o/R6NcKaH+96E9hiTKbTMCj+fkXdXH1sF1k7c/Mh7/jsxgyL6zHTrP6DEPrl8RQv1n/zNFigy2ms
pDjzH6vKVbRB4FOBSrJ9ZPovOMMYtJIST821c2MXcCYn+siJ1Ift5UdHec8e8uxUK8wERTgAQP2/
pBsTC9YpkJptgh4D31SU86LfGFu74mU7p9LV7V/P10tNlTiHK8HF+NzftDIINF6oX3wWyJicX6cN
yAQdqw9d5XF73RdET/qds/ng0ls8y+40ixz9n6Dm4jmplGxwDYxL8863Fue2Z0oZFX20KW4h+mfJ
daKmHkptrgmM43++80fTtH3aHjHp0he0SDoFf8W/cjgwkwGwnIWDJkGVVNH3vGF8vQNUyjtibWf9
fKccQBvS0aAQPYnQKTmIQFaqm06gtVPtb9Ms1kai4CQDaOdY738RiYq1Gbh4lR/RmyosD8nXRB57
rRVAH0vc3WC8gB0K/N5GGEpL/sq2kkpq7IRCFnhX+LyRA8in14auGvd/+l1senXXy9FfVxdeIgS+
3Qp2+uSVC2kVMt1+o4P9lhKY5hH+OGIJ1Fm6yq93nlqIxQkThVGC3QbfhXH/d/tbDmKE7nckiHdb
PTkXWVu/j5ciNc889gjbVAbLNMHntb0AGc7nNbXlNiqrk5kAQCVfPvKZ1m7mTPHQSK/20uarK7t0
0tsyMzzVZUenx95e9RfxjnqQl+KF4chuvi8zpr8F/cfyEnKqR8em4rIPg3L1AL++rvbdPdK9C3dt
yo5ZWOmr9upY9zgwjeF6pNx82QIvkh9Kica57fmHCTWt3aDdENbBdlU6m43lH9EECT9oqpvqd/AQ
dPZ97Ijz02BZzk0Vq5ipdGOFJuTQ3Sv/7iBoGTF+edbvOBTT+7E0xCDIy9KT/xUUCgKAynCggD1e
5i1k0cIEofPhYFa7vJRC7mEPyWIrtzv3J0rPm+1QaIBMZ5V8SGFFzLsz5mXn78C/aZkIbYzqy+5U
Zk4tGeJExYSrxvPfPk3AehJodgsVfqkvBZ0U9w/Q/Bym0IhZrwT+ebSYHsFJY+w9/Vy5hEJG1lX/
rleP4S4hyMrq/nBRTMc2kpMg6huRN3W6MVHOO+DHy2I9OUqqHwxHk5x5LLhEQmjLHhFPqrgbfK5h
dBeqNFROMCu++P1f28BHl0juE4x/NDEwBZgJVvQpcR7l8q7ucqSzW4s0E0yT/B6VnWTwKefSA8dx
qQKzlnTFYFC8ouI5ZUf7JIQrBAAiCTAJuLE1ymEIpZsTvZCc00wVFqOzzLTut/VO2b53iMV+agdd
7D9dTMowXsqUJkuM5G/Vsm8aLWW1vocXXtIs1q63sgzUnD6S1Y27Nahq5BdtfOr3coBZdk1eI50w
gU/IG2lSUa2sS9vy0RT3aFiqZizblu4RyqF3kSavcpzEa29L2xqqks0+akBjhpWeO7PYbZf+/Kvo
GXhuRf9Xmd06xr1n25Hr2G9hUiak9URf0CyJ9tA86RAXhz4F8yz4eaNAMuqcNtmytVXjRlXTb5ss
rLzQPVB1hWyrTaf/W4uzA/g5iwpquwE6yO2wjoXSdhDk9ncHnG/XUAe5Gpo8HVfFAWY/CvrUFLmb
DtIF3PYUpy137o2M/v71RKGHpdr6RtTM53beGgFrpsHEKsPGwUtxQHOT99aqUfY//Y2CvEv8Lwlu
R5BMnxdn8SiJyd/1ee00o1hJQ5dtwSkYGlVUvpwoUwgfgHcgKUC95ifpzvMm9zRqgFuSrG5GjY31
pcjqC87720XiTebo1X7+rxwJumsIlrlM1gSkom7qU/WHxQnn92zsfDdW7gY9+yVP5zBpx4Fg2Jo4
Z/OJNyaobNC4DHMYCDHgRuuU8VESetvG8YBOZZKNInto7V8ONnYSMwtovdHrEkZrd1HXN2O8m+lz
P0MNZPExDKRgcTPHKmQ3vmSkNK7LacnYikekcBmkQt+7PES0NUrFlhBzUx4IbKh7IUczmtP+5ook
2WydiQR8UxtAjN7Zxl1HdILsH3fHPo+fOgWokL+qiee5H+wZ+K0FHZCodpOqGBzEPLY49h2ISSHb
1xqUPb9FfYi9nJSqQJlUyDnIoHyE7K/rXjIZH3AHZTvRUjLR1XbcSANwAkJTntWurt7zQvZveWGz
03pdjQLlPX8T2JAW4O5lwtp4WWLt27sGUvZG3nyGzRFruA7VvRF29GOUQXnGJwW+32FOgD78a3A4
kDblx/oyC7GBBp+0HRlDq3BQ2eyKKerr9UDWRf2J/vVCpuI5kMPajO5HZOFJ7yVzZJeZTKofPkYw
x8fruSRTCRmx11JPMuEJ2H9qdxSfnzBiiS0mSYuV6G4NTehTK42/v1Fw/sLr5oJyLABmtMNL8MYc
cgxu0hHJ1I2+q96OS/0KyhaRWAs+nBdrEZH1NJZCfwFlkcur8Qqk15vWryWH7wdDExb5R1b0xKTL
rx9SBLaIDcBKzYaXy0Dg+YT5AFgHzB4a0tbMkDvwCH1M2Sik3b8aiJkgUuolh1hWyIFpteFps5qu
YcUM9PUJiATg2yGXQgHNctfstkm6rEN7vegX9zKSiMwiEnR5/6v7rwMqWx/pu+btOZlOPF7Z+n5A
FdRiHDQFeynO7S8ND6jpvSoDkmIax96VtkkWAYA4b05xuNFm+NPy2c+PxY4cc4b2tT+2o5+C8EH4
yXkCr8LeCuC2Yctf6HKQSImMWXj7otXtslt/M4MnIOeTkBLuBFVBdOXjmePuW6Skg/Zy1emxTvl7
e5pBJxPeJz5KdtqqjnK59n0+0we+L2MMH4mb+6HsjVAox5r+SveWYtul+zOY+3oMJLi5/V/yEVA8
kK8cptBNltSzbH31TiyTI9nomywMIDAdAZozH5gnKBFGlftumGDtAuziRf5DkmI9MqioPJFTHEjE
gYrMLGsPfWKEVZk5jpnAXGoyPB1HZu1EB1nio0ZSpP2VV2QPBjBdUyPM/4kUbLRttH3bJohhnD8i
M0yFDFG5CPYxizqCSkcIJWxImndLEi+ccdmZDVijDZpeVM/XlMjarc5UiM14XrVjTl8rC1CfyvQU
FgEV44uIlvEBd27waue3LJ6tkKx+GVN/EEj3Jwglf4rhiqgSvQ+zbysqWjlGrVf8Y8BaEWH5xkIr
3Jl437gaH2tSs1QlR+C13v7xA4k/wukh2mzF+sayO1CT7DjLqn3ojEnYQh8iWB4gsd1pvVhhYyXA
E9htBwUJZgmp083YBbAIhqjua5FwzXQnWU6XNmNSF0K21dncfg/JrDwEHIhPtdgeNs/Bs5X9JVuG
a9UkVssr6m88/CNksiyruL5iO67ZMZJodz0MhdVgFeCNntUwE4utNa9a3LZpfjpf7gDpie7CPh+P
dboS6w7NQZ9UK08l6YCHgKMXDg8biyjUxkSpfCtvT2ZxTAGcup+fowoKWc2aevo8mAiOTimAEXKP
mYoZ+GbmfbKUFoT0SxAcageA8G5KojK0eePNpNgeUHeFDvt9qdIa3ryxqt0on16BbBvItx8rtQ/d
ifiq0P/+zTvXgtNEjyjYzBY8qvTK483RqlVhTzeY9wmun051+CP+uk4EA8MNCXAiqWRjTrMwu2E0
C/8edl+MzUlLKHRaUoAJPxpVLljH4hGnsqMm2hyXrIONsLi2XVHDUI1gHys4oNHBhlTMIGIlkQpO
MHEClLGI7/JSOAVDdZ2qg/P14ekgXBnaoFSxvefoWFHg2TQUCG1NejcnW+uoHtp1WTWgk9YGTLfx
1m+MjctKx3UXsXgcqPaUTff9S7mriEsZrklgfU5H0py8SHcnw5OoH0aTavBbMxJkt1RLgVy5HmCG
2/xaYBR8i5DBUUqp3Gdp00i70hMQolMNZwLa8hs0EK1jlb0HgHg9wHWpA7+v4WOBbagQbPqdjm1b
CvuuOB+/cFckkUn8jiIhzTWmnSxqjxT52z+rooszvFXD2lRj5uOp+xwNb8IscQtZpn/Rt24FsB4G
8Ag8ERdIs+ma3nuKO07UBLfwAGzLhw3FL2HM0PRRP88TtK4u81QchSeKCgUX20nVx9zro7/Xi7Dn
JlNJPy/A6iVuNleMxeat5d1D/ANJ80YVlensKK0ph2ltBnY8nw3u1C7EAbGognqA+ADzWThOWjvo
Y+HywZtz56aVz/iplZElslQS/k6UnlIF3ZfEM8yHltT2AKWiWyXDznkVHrAamNEA66Mj8zmx5us6
eD0IjiMb0DdGZ9ek/d4a+9D0HwoYWEcQuZ+PQQ6qJbZhUpFp2zWizQQ3ySBRRxVUpWV88ds+wWiE
Qx0yHQlwEW0qVTptJavEqN9WuE1hg5mvd9YkskzjJoXgmxFxCTyNnPEwE7qUK4GC4b6nDo5X+2sU
6LlSQ7/x/J+2RRZpqVPUTQ0CK9s32ZZjPhnmyfW4BvEw2uLxyGWcbvtsXmZEGlCleR5aRs3WehPF
rg5PxNmh7NVHpfanmw3WdkIgzUz0kiI6yd7RhrdvnZ/GqhIfHOKK7EBTof0geBhUMrYYzw9cGaLo
2LoE5N9LialFCn3u5692fXhb4NEQAasCyBBKUImbcv2TT8lYIk/YOlVGxPqOE5d1nthn28xeiZKA
0RRnxt8H8vCzIQTAiEDyB0ixsIfXw0mtbbW7uEPLsi0s8eT2iT+XDPGglsStx6JYUZUaGeJ2RHd7
62cgDxlOv47xhxBSlchA7Bs1oVmDqPnSN0TOuIDMfjQ0gB3wwncb5yCg38rqRY0gp+lHt+Vr5MTD
f9CfyDzZA/AMkfQBLV5Z4iAKrGJnjvphjVWcrR2y023qWg1WPZtnV5o6KPCgR5BlUrVe7pKaPdGX
F3KaPR49vIYtbLuCEFt6p8btGpY3S3e8Y96R89T6839ErOsYrTrV3SZULLs8EGgqydaqhttojPlP
UYKkXDpxZlhZgEvdCuEsE/0uXCB7I8gAEA837iGJMJL8fSj2EDJmvZWOraVidQM11gKMwdVm/TwN
cJJSYuS6jSW9ZNVdGxkI6jU5LKOZHfZ4Y7Kj65e4KZF80DM9JUq9bcnzvbwXMDEhzV9L4kH5Pp3Y
5oQxENW+j+ZfZIeD5aLSvgSJ65dQRSbl0imK+iv0lBcFdUIDtQYR26rzm9CGIDfZuZxsSc0HsXiQ
kv+k8pM69LJfZos4z2KSFMv6+Xo8NqpTbx6/0xlSm7JFQrC1iJhnGjv189g48O8JpQoUOADA5oAC
7pFijVv0OJwKku/SYi0A2v7C9fjRlBIJEj84R/YX6qIh22ikg7mQ8r3Ri/PVTvUl1EZasls+hyJ3
QVUqRXhWX59ufoSDV7bMhVRgGWBlyJjv/19lsK7X6bIRSqsZGsRnInfV2ar6mMdZ6ZKI1IVeJJjP
hb7Lyoo3KdIdRnk1fvoseNsYI6kQRPcHaeEUIVFsgpAULQJUvtkGnWWnd6ELQOB20sk31jWPvWMC
RKeaYUYw5Dd0ZTwOl/a03jzLBCZ+LkOazSAhB4c8rTmC1wt2PueWU1pvl9Kdc/wOzKqTi0SAmtL+
G5LE+NBug/7/STMzreVI2MosW7yrHoXCDyrJE36ni/EFQDRUFlU0Ja2KspW1mqX5ppuF1CsQlQZD
66WnJRiCZdTKbFP8ITEa1Wq2SaDFeTlYkgpw2WE90H/B22gEoiO2gltf62jf/ogKFc17UO10rjOU
tx75Kj82yspbJT5z836teB2SQnEzFJApj318IrS/HpmLfoE1Mk13Yl34VkcGc+JOBy+DZTE/AnuJ
94rXkgp34ghMObO8NBMAZ/Xfs7t4c86UdYPJDWSkb7lzW6MOGo+eaX94iMto135wUx+dbm7zBizk
eHXNC+MJPDkC5a9POYvcaD/dGwJxwiNXAupyBS9kAsn+Rg3RbzeBiL6Y86C8kqSFIA5o6yX/aWk+
5DiiB1kMkCDb5NkeJi2xfVc+tbFm/Gm+kWU9BvswkPByG7Hb69+9wKpSBmPksHJgpIYNyBGzVf0S
q8xypECT9xD675xslhtyMuT7OWtMMSB1QZjWDzMgSF2LZLV+I+19rEgsLlzAPyEGQdlc8jSAtNYp
kIvuIB9zf/dKWm7Ovh3d5qvZGZyagL1yw/cz5LMgDwkYyTzg79T49j/3mfSOHw+QkurDgnxEM2WF
isgfgsdKMw7cQMadfGARyzk4kyrcg1ivFeTMG7vb0wYGtspwRtfzOtZM7ZpKmqT7eLDYrrvXPvJG
6Rlpe4uHlhdlVylBAtei4VcfTn2XezuNYZLBSmRpKT8M5d57+nQsYQUXTcVenx2TcE2OQ9LJQB7g
qFz67OUIGZ3B4X0y9cUUhpeqGO2GqVIlOdFrauPJucubc1TLivwHhWB53g5NgqolbgOSBCvi410n
4wYEbQDjljJ0uvAm79UaVKL3r4aKfn3qdUdxR6u8DObw0PWiz2EOd1a2baDUtRKfCxcjS2MHw7rS
toIGFxjd1DTxbVfibzw1Q3MyeegCILMQ7x67pYvlg+/lohwo8O+3HgpGW0FUqQrgQ/e94rEHyXqK
HLuW8yQkfRW/RvneLHIQMKpH6Kv7RIggnfLWAa1ZN60ZIrrP7jSq6cZtfkOmp5UiRenyCZE1qfNZ
2A60G7A2Vho97c3SKim2zFPq7wHHdWjqmG0Ig+cYehGZQJ3MY+zTt0CoOQJtOMGoi4dhhwvPvLjI
IIf3NGG9Pv7Z0cBKHQabAcpY+1Dqtf1lqzNG3jmjsebyMAqOmYiRWLYYRzITc1weje2udYdkYPHL
/vljwwPq0NllMZbIQPo7Xn2/msaid/Z3+NYnF6QcY0FZ9haA1xC20rDkWd+VmuklSEIGIt2BppzR
AjZxdSJsH0qJxH7Wx+bqsSaVuigXpNEt3w51mdW8T+Fc0O72PLZBV/5HC5B1wn41OH5W/wdtyzcd
5JYvK7Sp1dpsQ82DnkIzt3weJJ3RZqT9zXgRj/r+3WeFjoJKLszlh9azu916FjY7vztCdOUlTan+
Fv6/QOo1CZg7CUEWWoAyg5auBS14Js29xzHcJDHUY3mceJDRTrFml3vHdF1EGY+aMl6HkFNb7y3y
5OWftzTtINOAa+MxK31CrXgAilTtHemOZuD4jOM4kO4Nv5PACISZF5hwVP/Ua2xh/ozK2KCr8Crx
mNhpkAzYmJXZX8OWEWx4FgUqTtzd4JaEatBf2iNZHqf1u7ZX8ZhpmiH/5UCRHPk2DIVBS9/ajCfP
WuqcXbrFFrma5A/iYdurMewHbmAI8dNz429q3OHLRRIyEulwuRsFxkVwI1l6KklyAels2Z9yvhW3
q9DHpr2Te4M0AKplaHlLsG0bRvqeayxCh73sW/t6sEcbTPXEpwP+6Dd4gB9BSf4MOwai0Ack05Le
VxswQstx94/mHqT7Gsfot8lXEKHTYx+zaUyoplYhimyX7Wxv6VG0ZxKnt/yPcVENbyStzrX8xakb
fjXHX1yxiZOzORuhrQAzgGIBic5rEv3/j7+cJQR1rjm38c4jVl1ks0Zptv9jkos/zWctWeBy2EnU
FxBHZ8S0chGhpGNrMJQeEfqkU62fQ1KbsRbBJY6OeHyNm26q6a+AZ0V2k20I25oQ3lLEh2DTDxo2
+sECUrz0F7NYZ4uWmwUd6pyvEUgSHOe4N5WKXOXr0vWNRcs9eP0s4QQ3OG1GcKa6u5zwikh+h+4S
ZZDXLn44S47Bm9BBFHG5GlTGhufKmBM0PTffInqXWBDk7+CXtR/TjK/o+oe4Li3EAaJdhwVuUCts
LiCyEf5axODv7Hc42Ea4+/4tQbJQGZCZckyxWM7smkCdNrIn+bFfrLgGepkzLiN86Hk6NGY/z9wC
2uAFM3g288dNd7wLrIuu9JB29jovi6g1Gidi3XbRrz51iDDIBcFzO3x0cYlx8dgBWFttCgaBVR5e
NHRyREPhQXx1on628/5ZcZT5vRUcUXlq0A60I7tHofqfctOmoWGa8QgIcaNiIGnrSKbSzrwmKoYM
/VnhCUuiVvH112aSzAcP18CEumWD8XEitGNm8OMQbucoHCCE8+KYIy8bUf7WNCfjWtPo42G9RlZE
FRBLQgD3hX6o4KkL2UPEzDArnvCIm6kz9o81RVzO6D76OBgu1D8iJbWw3SekiB2E5BgMFHyABmlG
NbqlyEB7UyJLb2/aWZvb6aad9s4DWXLNpgprQWYmC0Zv++tp/iOrEsT32MVTzpemmWWK/KU72hcH
BQ8WkXxuVSW6HG3X0wG7z20K6eXJ6m76xs4Hi7V9YwoLzEvKT6gDmgogfCV2aL85lzF6uK0oz3+Q
+TmSqwHFivcMccjjTf2F1i6MetP0Q8Xcl5kQwTNHE/vk6BoaWXN0FxldOmySnfjD4xxb4gz9YSsV
lcV2/4j+VOOCIS8hhSKUyHUZJg03xDOdgSLxVQwRILzQN0FAJzrdAxYB/7YK9SAFE4gaVMqa7mXm
feqHCQGKy3lweh7+7p/iJATBS3CTWNNAc708BTP3JJtr3Upl5mYPabR+pPY/WOWjZigKk1I6rs8O
e3jGZPtCj5EP+JyuhVCnb7lkhfF3ubb5MSiXhl85oi7mENlLCSi34KdT+jtQFi9pSrjAIIJ5GFzl
Qd6WevcbksvwMoQI9hcbdASLFuDdNRE8e0i5QdghFom8Nd8tneHSrJmWWqhwvaHdSUjz9r3GgddW
bisE2qxiRABAApcMbPpL0ABuy23sGTEoAJSgryydX9goLSglsSphcaBDA33RMn1mOuAyp24bI1tr
gnAu8ol/kj0+I2Stxi27mvaekIyjX/uVin0cuVfPp67HINeERKBzlzawxGpdRs3qzZkgg5/qHJD0
BKtkRf+ClHwtXrKn5jKZg0p7kqhU+e/JjvCLlOVSGOKj/3QKA5XAIPyTwfvSji0cR+gkERa8Qy7u
+/afNsinGjCYj87CVEpnwhC8TG/18KTnKivgiR0+Jv0Cg4h79xQObVBTVJo2W/WL5R2+9z0qKOhK
PyAQ3A4XWwSdfWO6S1zWzEZgwTEhwnp1QCPZsDuX3RHLZkYxd//e+UrLp9zCXNWifzc49F+un9pi
QQ1yqo7B8Iflo6dkHE+zTMd+ZcMPN4HtrmLBaaPv23vzv/50O3iLu1vVf5Sv0OUpQjBsZjY5fbkn
XBzLm3qfpxxlJ1keaFOToq3PrI2+JClRp+E5XLLhuzUb1JYh4ANBbBtdcfxoqICbzZpvCa5PZZzS
q4mkEswHqoaeXX/prv7ldKejrZw5PldjeXLKHbl/Bhvl1eyLG2g8Fuz7MffG3XkQc4UWvrDEw+Kg
+dPC0uiguGZhVndASEVtjSI7iPHqz+DjxtyzBgLKvyoXaqAYqKQFw2cw0d0cbur9/Al3GsxXp9bu
mJ+FMp3zXNJ3BZXHSDD+UX6QRcmre6FA0RISJRkc/kMsERByOKClQoBjXOFRSjx03v6fy4wmJCqS
/llZWBO2XfY3oRJTJUQEUw3JUsB6y0KZClJnqiFrqp28dOebwvex4oapzDHrrALH2PDiPSSam0KF
Sog/i0nmF+ZkCRpz5qBT7UkjHfQX5WABK8lgTbT1SOJ1VJfJOZg4d9MtqtOHYf3Uof5vVzjAInea
CeMX091A3BBCQoK3hXkhQ+t8DKQoh85L3Q4U97Fgh68NCpIQTSkPz9F+FzovzzRtzhF4CUVA7AEW
S/e9TIw6jaqqGs4C7B4lDfaafXeSIYz+YmGiy07Z+o8MNyMtcnirzmZOSIM3zDN++/3pCHrlImPs
ViVfwZNxkURn7Me0a8q8fdaCgnXVExjyzIPV91z+mDeZBmKNNbPVXJNwFQhoXzV66/Bd1B7lKQH8
H/LaHmLl/gX1ZoxdBYgyd92wkuYLTZ1oF0sZ//lQTttZY0QRnKYm8TyQl2FyXtBkC7kbV4M+0h2Y
yHT2q5krWFCRxtEv5cWqICraiWzhD2p0PZpfjYrEQZgGYfQoYEgvgyRIDZJra19MFGjxfNeEvjqf
gtgYNKghRTocebq44w9EKUBf2iohWi74Lt1f5o+oQ5pXtd17yNvS541FgUfs85sNSAXOUJHxFyO1
qgWWAYoNCJhRqf7HfRFIjvWJSVqwwqLhLpJV3lrYxCVX95cNhi94Sxn0/Y4XI/c4IBGmex4p69RJ
ObULf4V1px/NBOEQI2+MA0DpVEHO0aRIw4uYjGFYLReHvqiLKHb3tc86ZKxKrZKkrnno8rIKdls9
dW1CF94jcX6168ZcGBI0uat50BEx/BITnccwznhlRkFVCf0vj1IdWWF/PeTPgFFd/GoSuKH005pq
dyqDzjy8sXuiInffGQwjaNGHf8ePKfnhzxiSdmjEOfQ9nLnufBGTHDVGYrHHpdgTpr1U3vPrdMQu
/9akA+qkvRyFBDZYG7DbdgIaOcjkFhfBZWehjQjBf3p1acB/mIA24rLhNBK7mF2y/CjrpOeIE68f
pDMoL4jVcbjjYDhWMJDEkm+9CnlUBI9vpqgXZZZcdGcIGJqiiGk9/w9/f6wfR+z9QiHeR2RQeuNz
rtpmPJhlUfO0Y19wceMmAJYktZS+l0uJGQDXiKVub9Lw8GZ4DM7mnrdRiz2JH+TcxVJsCTSpR8JB
iM26XZVm0Sn2jxcD51MBpmyz+IQ9LDm8VozbkZ/4JgqSva21fkOZtMYDtujcM7kKF5ZAutjOrXF3
6BrG4rjdkpbfHzfva0lAtueuc2sPOQTkjRdTMPBaPUWcY+oI97n0TUBGzUAGrw+SWiL+14AeHSmQ
HJvhILYcruBd+rURCivcDBJFgPHwpGHUiWpwNhBoyPJRc/Or2K7NOkCI8qTtRhra6Kby4HLkIXqO
PrFD5gO+0nn+Bd6MbQZ8OirVRJefo266S0oT+DEC8c6lt14aE252Xr3rLsDKCJ3Jqb/6j+w/lWpz
Aaiaae5gR9J7Ecb/AGR6wYBFkq8Ve0vocywHOYGUogYczIoq+G3YAWVJR7805bS/nKnc6OQoAPxX
awH7Vi5nqlQ6t5JbgkI4mGigRaxjI2uN+VJTg3adqeJyq5PV3Eqtjb6dYEZlf0elMyHQNyCUSUKD
QA8NcHM5gh3+Iila5kGNnMY1G+ij47WvVZ8hPku+jbyeP0T1raWSfS1XFqf/Zd94bJJMLAnnb4QW
UxTldeh6tuCExgHRxxRkqJU29r13QY6y+UP8tSbBsoz5vZeNGRc1CufZgG1yJ6IhSnEIW2H9Kpwc
i8KTYKq0cJt4xbICEMQDPYqzeq+fM83O3v22koBpsrRfPLb0apE7qVTp6IN8jD98InOFwq0WSNYR
4VMaBdz6hA6UVvu/Vxar1NIYwezx7KALRoL6c0OWRwvsK/lObVSREjKLgAM1/k7ZzDG3kmSZoSE9
0w90NjfqmF1OCZwezGhrjq619UdnNtOlRU025waOJ61T4m1RGlApb9Z/QfbDzmrx2cIG9QUNagxj
rP5MmxjjUxcNE6wjcOYeYdtHXuj5gRE//yyVmNWnhk6xK3FPs1O3jSG2sR4ovb887bbNp4m1rDrv
aCA5pMAlN06lF2rSXnDqkFfMdJOhQq1N5TWBkDXtj8WKuL0dPKI+pJzb+tr8tfIaEYZVLdkarLPD
3D+4D99KhATiuzktZIKcGDikElhyaoxq3fxtPuLyUpEiBJWKV89dLdeQ2clOjkUSF/blSO/DsX2o
nixlA/tnHfDC8N6ajafOB5P2YpJf2qLVR5CJIPMVFw/Z2TpjilzH5Z3KKFvYFjJwi6PUGj3STkWf
PZzhEKvLe56G0hgA2My0a867jXOtPeUHE4F8nijq+7T2Gqq+zcWkgvUp1urILq7htU1VuWdmxo3k
zcSDiV+l+dNoOnYcSczz07ZfK0Up+omjHFBqfzMvAhUEksTMTx22OVpTiYJBpLcRKwoqdw0bNJvd
4iBw6FF4mbnAwDN0vJtiZIYCwVWmi1+qu5XWkRGsp9QLqsqD23Z17QpJXo7wMzsKlEFtYaL2TzsU
LJubbZ7IhT59mRRGMKwFBIV+HS3fqyL8ImhJa1+zaAlWrtU13c4lpTYeJubbacDkhWIEuN7hKpKA
73oydsc1UL2rT8d1BJ8Ez7tawx8YGqg/VTamJVGWKo3upUlKK5bU8BgWd5Rq3j0FtJNLku0JatqI
zNGqLL98Dbljc29TEAjnZuqS+CrJvs+6iAeHerGMpgIXIl1eZda/2MiCSuDEEPm5+Cl6ytHrAyy0
NVmz4wx2OKbxHPOs3nU+nY+ry3UOdC9Yj3/1N/pKxxcsqLz92gNlybzbg/F34VJXC7Ylv//omikN
vJNRA49F9+QRkPeOuuBg6YYlAgMQTgMrYQz8/DCp02mG0Ee0qcgqgcTLa/8rD+CIOuCGH7pzmgzA
7hfGLg1LmM80QM995spa/rnA7uEKP7YXFOfVmmrK64PBKItqIBl2oPfIee9YXMkhOXQi4V4silfI
nWoqAR4Sv+I9UdhzQDZjZY5Th1NnFQAHVtLTbhU/ak9zE899QRD8iQ8mPm2evhIX6TNF9iEKjKgp
hF0HXcyt4Xtw9+pjcOOKg3s5dlRenoiKezuVRzJd807ebiGGJ+w3S8wDyAO3Yt+BoiVzcBB+K5N7
vOkfYmx3opVPxXn6sO3YC8NT0ZoxJo0vvLUwBUSU78X/Y1triAZmFnYeiap3/nY9u1N4NNglGstk
e3Uyz7bypNSkj21sxr+eOPZm1NfWGfPguIKqJ4HoQOF5i3Jlb1jZGu5HL+lRSsdSgu24GE07G7UV
IdSooffOTueI1Amxgfd8unXXpbXw4XKcu0SNiIoLv2vlYPjE2S4NKsnsT7cGCJPRlOeNBi9HLYV7
QT5JAVhzchNjIoexJYNRo1wtFb2C2VIHLSbziMoaSmFmSIeJhvDR8G0OuMp3cTGsHh9U8VtbFGB6
4BEH6fnH9whPPvnpJ28JUt9008VGIc0WVJlENLLHQFOy/aSP7kUGJ0YTvnYCdxX1JeGiAh6P3qlj
B1epXE6PT1ASfiOQzCIh/GEWD9Qb/05wijDeI8EolKVR8Hl/+jNkYW5SHTTOfslIVyIGaP4Norab
M7pQ9dDRLp23kQuhHjanjbRtme8eHXNNB+3a1BnQj1u2nf+R9IJ6Nk/SP67g4uCNhyLB+DWLs7V8
8f/XXglIXuTRgOjlnhhxAlQyeUD/oMdr03Jz+XPJDdDaPL6UeY6NDFssERtS+/oWhMISv5nDa3qw
fMpImnTSugaSRdVDLyoAvG8+dyj2fi//z1MnYOVhlcIo3YCJDlwad28BLQdW6XKcdfakrWa3hSXd
/4YAblejS8OgeEDUe6W4tXvnavrqY04R+jF5eBc08x/jQs+qACdfyAWR4EE+m4Q88aUvrmK/f3Oo
vdNhG7+5u/UCur0IEHoA2Pi0aFIYvwHG3ADErwtB6kMuYL+Vo3hvB1QE/DBcnARV85mNJ7309JJB
1nlPmVHQHOgkt9kB5QbU2LotQrDtKIIcZRY9bcucofGL9CKkd8S279ZeMfNLgx800/eKhf/iJ/Wc
ZzFG4/p4X7roD1UwNH0Uqq8t1r69JgZoPPcKVJe3SKNRtkRF54zC58ZwRSDKDrhhF7eHIZjGU49C
O4zsVsorURKSoEq/7Xr3WfgNV09+BVXwq5yLHSMfZYGiX1fXZEFYAOwA4QTtYGNq9876A712+uOv
kWj71fGHPiujEUnk8fM1mfyn2yJse9VaFwfdf8ybee1xDuhpb/Q0NQAXTM2w6n7vdHg9J5tJyf1h
xEpn6kyBq5oXw7Fl56GlLGgExSpX6TfER50zsbPzi/lD6hw67RtLrII7+pt409dqhNypbBBJdbYz
+Tuaoh6i+1msnEq7cnNv+vgKqTQw/7mym8LiP6mdDcpoJ10Gds0NtjVuTpx8wgeO/AM6v4gyKCpe
1+l9MZp8NGXTuDgtsghqBNvT7TV8NhET8vrXMCsXBUQvRHArRRadUWFsvewtvFaYFi03X/ZwOAAG
1M53mitq4WMGo8tNFKh1HjNyMQ314cDjxMjjUlRTg4I3lNEN52/g+BOrIc8nkPwmegzQUukj7NPP
o4pw+OviyUSucIo3hTbbjq2Yx96KcyHrBuH1rYRxPYRHPqecT1Xggw2LfIakkZh8Cq26xWQMGWzo
Tn//tWq3VeS7C4vaOEBerHQdavBSAMcEGsnRKyIqjG9Rj/q/HAlHm4dPJNdprAvgl9ACUbBux+5d
kQY+l0AD7QJaLXz7DutdUWBsaH5WmVjh4kG9fcGB10Dwb8ulU/Zv8KXZaGohN8mKFdNYKkjyTXfd
aHXSoRSPbZbp9xxhY+cJ2SSxS3kkkvZqozlHxPKREGiPTJGvUSbF43GsQPVcB49n00RuMdTZ8yJd
tQyspIyc3yoqNxefWOuZ7/umu8ipOq8HfDdEpNvd4a2wL+oEsTkBFUzJTblwl5P73snXI9zTetK0
PSSUii9AkhFqGQihkx3YE1jKxp9ZebsPd1ZGXnuNbcOt0SnbklA8BNzaaPLV3TEuPaFGC9siRYcV
DIREFHoLCxku5t11KIk7zEnhAodIGtkGNFlY9ZDuuqlBkRphrW1MpeisGcI1dUf5iXZ1+G27Mizq
PWe50yB73rz0aYp7RaCUMzrOEiVV9ArpN0G0/FjI3xZggaYwVBEs0wFVEYnVVHH7ijpKqVkADSYv
hNs9qam9RxaK/bnW7LNl8XaZM5P15/NqIyPOAaNNPtjyWZFG1JrJEjrL/JyKVtHSYor9XDgrkJsc
B2cL0gVu5Zp7vre7DaiF4J3Vy4w+MuUEu4rVtgNpDW4/z1uWzfdPvmIEs+Gke33pSO7E9SXHy9x+
tb+FKpnWcpmIrt57VhSrQ45zvynGJmxGlwXTzYcIPEN1DcNYYRBJGHdoFEFFjb5czHJ5Vm9TWFl5
LJjs6ADqTQQQP3uEg5WFs/GfK2z8492ZhB9lyQfzlyGmNUN7sb5MbbrDOyKstHByRFr3Pzk4JN+L
vPIHuj9X2IWA9Q0j3LRet+KOv8s9o59kwwFZjDKe7uUlXsprM3nnCJQNl+ZGriPkHxOhEL/jhwrm
cUg1B1xLI/BWT99nozuoKschfQZL3pNyzOONDr6c0+L305/c9Hh/IN98U3/sgNfZil26T1vO3czt
BbVWLmIH3tnuiYwVcG45LkNGhn8J0+P02swtgvLCi2nhUcFvua7OcShBBeIhPJl+8fkRU5/r4wCY
aPTr9LftZnoxb26LJw1Fs+GujJAJ5kdvXDNgQifdHECdJaO4OuaV291PSl0GYL+4Pu8AU/yFrOkF
weiUpiEO+jU8Cdap4GOtL6N5bgdOorALInqLZ1IKHraBGJPl5zaSUliWInshPlDFcE8+pR/M4IVo
ecSfI6AZzHi4vpLCnh3ZB+2PA1W5yKgB8Y2K0zJUSXqlcqLrYXD52PH5rtIlr34dYbD+fBx6ogD3
BSWxa2GIh/sVckzftG641wsni99sQVffxKx4+RMw9ccvJI2eWAzZpTOIbsfKhrlD9c7pY2NHbKyT
KU81CPXiZ7jjNggKTbMjRHxY6yo2TjVoeH1EEpIicTeOoSwDxYfjpLIAx5FmT1GePpQBqLiSgVT/
NG8bfdZjnHtOCEmpEUkj3+/wul7ZIFcKfRvhweoEGF6yEno/N10hUbsbgYS+nYeVZkBwk6rV0982
H8esL5gGjxMjVCrL6MTd/rCCD9rq64eJ6SX5PIrALA42L1VPC28mF8JFR3OpUs6Tuq5OirAzFnXK
m5mDFxoo0u9ME32rAn3ync8rW4rXd2isXH2ySuu+TNc7+5hl+OXK0kDKJ/mBQD0n0rr3oI2hNnbR
SEpNAqE+Z6WuO9MFli2MyBRGrRC7udKyiPRVPPofbWKyr53qHYQCljjHUjMR30zGbj6tQEs4hnB4
htetfWxoBhDCLtU8ok88WRokH1fWjEjvPz4eK6OW98sCr4HnPhXr4if+eLQBpDDTv3NpKDViiIQ5
tjgqX+GeFIxvA1w/sIVohmw+H8SJMLCdka7HjqAGXFUbM4aPep5FlSb8KLvMZXuuwwJbh3wzcrcS
i1jyhHSk58qGxZmhciJMr5vAx10a+pEDv7EvA/q6UTm5prSFzSU7Ok4t+G2dMgAR3EziefcTSOzP
QysX0m+ip77LBWSRCqO1pnR8gECKQ/hy6yixfWVuyV67DUXC701QlAQxIIxBkXc7DtNI2lZppaGB
2qOJOkfNrmtEbl6LtpdIASr9tajmp6qJ+CrSlMr2itjOxFyul6N/2O+KIBp+wdO6wcNaVTaRI9c/
ykWpbJOgnfPvquEKgpe+saiqQgiTtyVGoQ2RuiYc1yiA5eiDwq4ZkIZFNelpWrI+br3HUPnLuVHP
V4oNsQWmNBxqc0L1Nmo9r0XLiGqXU/m52KyjEkEYCsA4jCb7t7cKgrRhp6RaRJxH3iJkQSQ6GOFC
Qh1gQbnsJiiHdKw0QNsGktJqEnOtAijomUhgbRD835o7/PN+VgOzsMS8w6kJMgu+R5YbacqhsNVf
jdHu9HIQWtqt3sjJKX0ROtBQnCXzdsVxVhRC0FqpJ9nOn9myEoA14cGrKQkZ96XQvyLPy4sqON5t
169TBtIs2qblRlH1ZSPjcaXagNKj5Jk7X+rE8MLcSnFGo1/l4x/i6BgOYvUEerMxKkU27nRBY0V4
xuO8wiwWYOV/hOLARuqJB3OBPLWTmbrkYHP+FMdzpCRsgmAABrYmFbz2HcOEB7bAQ07TboiurS39
qtRwIB7KaKasK8hmBc8YGifK306Q8wQKKhLDuAH5fNaSVDGyyssb4iWWeqQysY16shkzLzGg+DqB
lc94+U4YsJcjg0cRN1TBxbdYMKINHx9gERjRJ84W/Ce4ZENfgfGI25XhBV9VUkld5AW8cdoEUS5V
S4+t86/qBDolczLAnybxVHd4nUUOsRT9DRNj5L0CQyh8tyHiip7vInsJu5C77YZq0P6kcEP2mk5R
4TJzXO6Hm9nJokiPnnG6kc0pJIZJkhUZgGkBV8zGYKWSb46t4U/tf+jU6vpCIcRPB5c/xERRZKjr
8j9V2wGSEIwoK0/90YVLYLtqo1gNJaBcAc3DlSVcn7IMdDLZ4uweT6NRNliGKoNGdMlvpn9dyfww
HBCLmSK+Ri2DOx0NSoEdu5CKKUnUeq18eVxKSZf+n5vbAmSwTvF4ABvedexdrAsE9dZmYBxZXwod
vGibauSZZYzr+YSWyyxTuhl8jXIlZse4MjEyYDy86a0XwwRpojEXSlHUw/hepTomjyYE5zh761lT
j+hkaJUJKwHjGL11uYoAl3sblhAG98MmITycdxz9HXgPmbXt6mfNCpfFJg4MNqhcH0FK9hYUeLcZ
gCZ2GU+TGDIEJ+urH/3jHfV+j8Bp+CRTL2+OHeAS4pfFYVZ2woSm4FKhQG8xCeHfhXRYZtyRw0VG
WFlspXpyxlrKBVRRVqMnApn+L5SQEFE/3g7RobsXOY8cjESq2fhK+maQFssqkC4j27KYlV744S3f
Lm04RNq0aThdrDc0gbhy90lNNbEFPNLjFOimjZtTMYHyZecY6pD74b3ake+on4Wk+eoFz5Nc3njo
buvVANjaLkxcMqRu4wNYnnim5Wyzakm2fEFR5wCo1v17tn9jceifRfFWDaGwuLSQ0fBjGm3hHSYw
H5ZgRrv1KGCtAEnCggFJy9cIHwTNns1DA0Vq2YUdFxWjrD3Twc7PYptFjO/+PGLLw91hC+Pc8roo
X4oIrUALWTxgcpauDz0bGOZVLqxeVn9vOGDfHqkhhZagupACnwDiQY7LggQzzjbLL+K0c0+m3pz7
hUQN+NPuOabtac2wmzfUEcKr21EdiZE7WyRjKxw5dFKL8XoFDx3oLKqZflGHtYB/Rbg+ZHp7BYRB
4q8RIHwU0lPQ2kt1bNf4ObP91Vg4t9iv9WZJHUFZta4kNcH+lqiFqUEgkIym1plCkHeAzuqy/wRu
57kJQGUNiIdl2/7vgyVq96O0jtDW5r3mnbfhToatbHT0mYzmzBMxoGDLyOBUu2HEAG/zgRhQ93xn
kznfGG0lAKJ/FA3OfW0oHa8QO4GwNi58prUjRxeUAfx+pZUF9bxmIxgEEgYtH2qHIBVTR86ncGyJ
QDSX9yR2kAsILPDIp7y9bKMnWfNq7v5vKR/8HWnJGwgKik7LA0qEn8f84EW8m7uqh9zADZLcEmNw
7umRDjA4saUCYJLG09LKoECYPQsV8f1lgY4mkjqVEu3yGAzwXkwKSLlsFytBMvG6odW2JT3gvFyv
w1bWgFK72Hyz8plbeJJJt/M2VmtukRi9M0eBC1yWu+WwSemurcY7504Ag1qqaOzzQpLaDJdYHDwc
ld8u/Nc8N2SXYdzogaM+po2QDh4v43LI88w71EQRwA39ZQ6ph7DK9DjIg66PSYlBX6SMX5baQPi7
wO1f7yDSI4wYi0qu0NUbJx7SGwgCUmN3NM8pnARaDJW7z1OD5bQZeTK2iZb0EIRYF3OCsV+tb/id
zf7UmKFb09HpCizko8Z8XuXTxR2dCzP44jBoaxyl0wa7YQ2LQsXax0ooqc0UfRMMKsms2hcyiV4b
WrrfPT1yKDcDsF+IVF2kveAOUVl4m5cperNE16V1NTWMboKiHxLad1PrEfvww9XdGR05Ffvz+b6M
EVdICzna14r0XACCgxNOmio8fPZaVkGv9yulkd/EXB51CK4zd5JeFBRFgaxFa+mXR3ot6Wr0nfq8
g6TIbPL0m+AvwpsbPdhSLMzrJuAalzUaKAGPlfCCB1AwDh342LqRMG8vlIFbZ/Lsw3mhnorv6Vnh
EB/0TPduHy6sTvRPiZG5/y1cGYpWqwkUZ2d+XLhfp/XEPc9Zm6jKT7pjYPijZJmtWMf2/YCUmjLz
bD4vPqNg1hi0wxyYIp8RCqGC35vPJfw4P8UAUG15sQGNGAIpYpuCskaY8fVLnY7aBFQV8CIuO8ZS
uCyXcHBVhViqrK8E7z66nfBJ4gkoaFBwb6f2oDTEb6VVTXeXCk44tAdCPqeP8Px9o6xurzRt1Vjl
WPc1jgGtJEIyjHZ8PoGB04qdojpQaLqbwK5T67IgrPQa3kyFERxYe7UlyoUNxQjRzRJBmcJ3nLxc
kp6mzYTd7hiLfMdJRuiJ/Zf0WL4oDHeALxMSPH8IuxAuwGDIb60vrNLo7ChbnGnRDLZeBSIPbBhQ
kcgZjXhdvf61+2USikLx4C0ehdigsQCzc4z25LazeipmS3PBYO3rpWGpezRfKU+5o/mVYGhpLDMX
0q0JCpJjQ9mhl5xTUUtcRMQaPJrcr49UIvUw7G7GzNMeyvT4FR4il93E+JBDpArxYF8M6orO2sr3
ZISpWg3KFWoknnN30RiSzJ4TJdlXF+d0nwgReMGwzIo5dMtddkamSowZtZLhxSHkE/Sz/9aenwke
18rS15QAGj3HAKCe0tb8HNXvUkxHIS6yx6FF9D6L1Z/tzLZRfVBvpAU6JSjPhVXNg4lkgLZ0V7OL
NoCDW2LydZ/l7OlnKbnD+YFJm+SS5k5/+mxuiGn2zBoyf0l6/RY6uZEaEDC8I81s+ANrzHFdtwFd
uhoiRNQQZsd4Y9PuHb+HJLAI28nkkas2T+g/buU7pvKh6SKdkQbB/4h2TpFNmJxBxZXLSYmxoLvc
bpMWN6zF9v9bToPV7RdcgkJCQUzOMn0jO+b3cJHLel48wqkm3Zrcz1+PIxjyF9FAI+//Wf+TO9E8
pTzTCYVKyOLXqRLUabwiqP8sHRshuKriSeDeT3HJF67qkplHsC/tS65WM8KmJ7RdArEIchdpYTkE
TjFMG5A3pWnVdlWaDjc5kbtftN98zYYgBbh/TDQ1ZEStaKUlnqHSssFGtc6isb4gtrcUy6vTovP5
Xdjhe5Ygyo5+UBflMYNnLJTl/a5IL+MSXHWSbaJClnoX+o3e9YrJvFqm6zqT4fkQGAZOumZVfUJM
YUtnjvGfrlCHDA93cB/6Fv7AqSFm1Ej3SlyPcH04e8y0UwDNDzyjBst4c4jbCijJfe3RuVwE9T66
/rNAFkHo/m+UjqZrj9WqxVMpuob+q5cSzmjXoDww/kCYG7ao/hmg7oYQVPZQU9ypO49U4T/om8pA
o+mWstb7w9LyszNJsNkhUmBGQmciUNMqelAUhbhBfp2mJpGrotVxBv1SHRYzLfERPip/TYQKJ82b
9eR+LFjb7iTsDYs372fKqmxfZZjdrzFKQULFqqLDPtXmf1Hq2LbOAAs+9TE63fG51yGr/ALyiFMD
Q92uRa2BQw/gXLV2pIu0shnGz+We/Bb+75qm0AeATUC5B9zTnSqUBWAKJeNPvwk1pHPeW4dynn4u
esHja/E/iMt5pfLbfU3sFHGek1b0bRX+REh1qfTE0xUjmNSx/ibW1PeYugkPsbalFLvvhL8iwadK
VFJkBLsXOwLhYcVY3MjB/2cbIARUiN+2iFLZ/s2eA/sN6IDzZ0sVb1GbkKBVThl6Xe8GZZf0nPlM
VSr9nvo00qyOEQy9tDaX5H0dkQJjydjUJ+phQplT0bEv8QuFFw+4cnRPoZS4sF45P57lYnC1JgSm
u5IdHlYeWIzn5FX6Ou2qQ7NfzCQP+w3/xDAuLbTrcGz+UgdF+pZdgIE1XKQ6YgpennueQ4lLRU5w
BgvW1sy65aA3WLqZjkUDmDJjGemer5gQwivrmeAgN1+30ZjBPuWxk7t3dv96vT5w/iC/Ro2vYnIw
Qkenyrb7zKRuBaru13vcMzvQX6CttqD8hIb7lxfPw4eMWZSTlkNYHz1C4KyH1+N4wp7yTsa19eQp
gy9yYkj8AmKwwAHh1lNsqFOHBxc9ThqOFpkWsuQoNoy1oeRhESyMjrstbt0ZyyN+Oj62P9T7gh45
cQXob1aRgNvmdtZuqqi/Qbkfgt+ZWl+Jg39vFCbjg36bTcoMtSdyKzi0kwcoJ9Eo0vlhHlF4cAp7
uhPV2vVi/qd/NnwJwHM4YxUv48cseQgWAPeP0pbe8TqJFlOsmayZuGIjODnP89WpeEmlwWgIhMgR
3BXMmh7MeROvyJflbK20yb9xMTVaGyVrD2TMBYceZHvPxSZtUA8D79noGr7A3RRXgygXL+hYuGSF
6T3gnNm2beVWagKTZARMJm2+XOGyDMui7SFbvKoFu0KIfnun0nSY99yFqY8XdRyPyQQ6hs6NetNh
vLzpOJZdE1nKADUhQEZPzVCghvIm1dqujz+KUaqPk1yv6yVio+K3iHSxySEiYgVlKr32SrGiD1X0
CBAcrDOj46sHnK4uq6jyhBSqjWFRSM4E/WgWl/Y2fPKsBu51GCCArgTQMPJQabkgT93xrF1lT1UW
IWBd4pyHYvxVwrbGZqM/oqsgJjFlLfDnhv+wEQT/Rj/tZuo5lrGZVakPb6Koo67qWsqU5yNLDr/T
nUgsCptW4TcA4GlPFhTEO/BmJaAizgySqSG0aNXww0NsgIsh1rVIfP20g9bR74wOJIyoZw5+ojm5
JvIR6rG1i+I5lVu/KDIfFqy3oW7wwSAX8FolqeifTiYdKy+U1aaejyc58Ss7tu8uzYYSBVna0jil
K2/KG0+N8Rx9Tz1AYwn2oAMB+Qrs1FDkCV1Ud/XCAdiAHY6UK7r++4caXRSaMc87yG6ZcGdJ5toX
nHG3zwls6Qsw8aKxQeFoxZhAZJb15gXJqI6jqKQbybQvw5MpK9q/hi3DpdWdBHgWJ7NZcZaNyfuU
qB7St2zs/I+Pt1fQ+Zap9B0i5ITmedGyUq8x+OEJCFLxBP8bpF7ek4yPQc0HJofJW0z9HuXrVuWM
8N03RjdIsPusxCwTng55/6t17mL33QKvOlo6FZbcNqjsPuVle9hXwUS9DnqAhNCwJqghOMbI78A4
4LlqaogRAt/ZqX7e1LUep20sd1rJjLDIGw3sSWh0d2i6VTnL+yADYfXPQVtDY/Vjk6nZtkpn/Cex
brrI7+X0tNnsl6E+TipHakxh9d/PB4lAd92OZx2MM75abfeikfa/FTYckHn/2J/L5sFbWPx7+9jN
06dfUw5k245kPdTaXeT45AJT94KD8gOhYTQEzTsaCTIVSL/NnHCyYhaqpvOoMLwW/euj53TvbzqE
NQpD1iXiGxhapjw3I550TKesGM1Syfb6WtXfSZamJ16z7ukq+QRJy06usOdKP2krGwCR1UKCiB97
sj7UVBsJ4lHVnvHoFEebTxcWuja08aRLp9bJ18BLInha7h3bK1cJl2pUe94b6+XKXdgds/SMKfjl
ugC/A39aNBKAYNBIAC7xL9gGKOtiiP4XLQP7RWt/jItnSYgBy0dw3zIPNriQBPA33EqtFeBtZGIJ
2Cn9rFf/ozDOX4oTW6CA/UD/MLqiWe24gaMOZoAk3K2pZ0BVmDuzxHxn/S6NtR4StHEbULQDa+Zf
JDnPEV+Y6julMgl+Yekt7/iPSklofGqOEgqwmwTeByZXEINN1ygDyo77C3em/9wyIL+/8qWrANmz
E0413rEP3vYE5KB/DEF60eQdWDoLRbfmG3ZZ2SYZsGs8dLnZwZXL1/ibm9RE0UuB7EeUNJQYybrd
fJwMiZxk7khJKiaAhA8DUQwPSgLktOOdKYM7JyKWPMmgVX0/vVgz5lzg6qfWW8clxTagKwjth96M
e2JmWPt58FZJKqNrefzvX1a0H6i25ijX0ToL2LOUeSFRcduT5DiMzTRasye/XSh5YgKICMecEpBS
z5oeslE9cIAil+GFljC/yuRP+7H36nctftIczl4YWCcRE4UaXoJdXzk2EY3K/oUmwwAoVLBtjtPr
mvkDNuRLav124yvjhvnnrRL8w5aPdeP74pPX+Nd2XU02lT0oasZNlc+Iar1fuiNTX49sR7CiV3U3
R2h/bpjzQIXaiiZflFV6ezYz8eRHHUVT2KEeRZzwn6rFKiakZ/Kc4bhYzzGjuXJjLF0UAE1R+ueD
EVkgO2eJGNcDgLCtqnpu5TFF//wJXskkb0kn/FDeOHWbHnKZ+qlEr3kIlDa+xp2nfT+7bqRiTbQm
XnTytzL930gr+/UK7AJy0KTCm2Fah2x3b9gcjfZnIdsrEH7Oxj3NWXF9Q1BvLyHmWvU5vIBmhyRs
12uK/rIrpgpVfYMLnbJp1E2EVMw3e5AcHEN+yUhPaIFbOtSKV6/kLcmrcJwX9c/82saVui0xwBdB
kvCaC5kXWoMYiVj+EWDswN2OC6j00SzvQ6DiSur3meCMsZwySvxxpfopM1h40P4RVCtJAv+X3hD7
eBbEhbvbENpNe2Y77JsxsnqJel/alhxK9gXQe48EHqaUUpfbpIXdn1xvqxb+07g4iZBLsU7EyvZg
ftMi59w/hRH3Awy+Tu5OPGxo16OmYboOiJ3c/781vfGcf16AA6IXaE9/eelP5SEjpB6F/dox1DBe
Y+Fh1pksMQIbu51LeMYbSrVTi/y5CLAXvNQcV20/k9lv5TEqS8nmuiVLf7yCApFn1xEUqkOb727B
h5t7OTvOabEAXx57pvwLIwGSfsSSqUF/XDwcyblOUhM0fGoV/URw6N7FWAkyM5EY7C7CpaslS/dS
lC34orzMlN7v71c+mIT/nwgeRQPztO7oDhk/nj589WrE0IbG0oR3p50oxahQdlZVxy5rOmBkGOgm
KCaIElBMgo2I8qtv8fyvGIMS0Yv1RIqI5y1egEMt1i/X8++enOordxv+EWHkaBFKggM0aAkNIx3g
ijbF5wnejZgjXgPPq0veUIUc1wJ4hUZlbIYK+GF8tYiOZc/A23+8Qp3KVHXZFoX0T/VJHDovaX7B
cNoM3WMFftohsIyErYzvVODzuSYdAMkwu1pro56r/4/4/xKwWJFRFUh736qkQjVPQn/9iFKRdFPX
ZdAppChcJ00wmMOEMLPq9jup6hub0nQaPFkxCqi1QLVOKkKCIbfrglVyiz5f61EDpLaTaEcvA/QR
DxF5D9NHl4GG7wNokcNZOAdtyu+KFK3g6CxpqeDCAAbx7M5Mmjp+H1sjeg4RC5az1B49rvuRtryz
rVeTVjFza5TrP8W8w6v0JsAa6Xtzt4PgtVQaBW1H0NI/NYjwrczQWQTQrXfT0/A/F8YA9lL+9edp
POsU48lLbmtD9H2X7GQOl57f8mE7Qtjv3cjlLsuL/lBxuciCCHr7dRNz9ox2pn8vHBQ5mypdIQmC
XuU67/NYUz25MPI1KSncztFiv0mMAxSXeceqe19QMmAHZfu98tRBct3d77Dt/ca+zCfaxfLrYYgQ
azDE2mA3T2dATp8wcRjYDZm7X86rhQ8D0D0C2+Ev9jkDkmkSUzpI6H0uVFofE3E26SHiQgn2xphz
x2zIuwZPNdTOvjp4Myykei6zsseN1AcQ1nCKL3HDgrgToWTLRsHeai8mbpDISvXAzuvOmExmvw7h
QzWjMI7yn41EzxR79epFcyzNL18BiikrkKNUuNBf+WuCrxR0ZkcUpn0ZgtBU80z42EABEho30BXp
k1IRucqqIU4Fp4peqLdvdFu09YicGmFkZYE1R3kleDicu0nYnLl+w2mJnT/E1cekUXezZXPUnptO
TRYoNXSvANrla+ZbtSdQ5MCCVoF89ZAlBs/ijD6xNKxenB9utl3wW9EoRZtEfbwHZcQDOD3aJfPw
RvI6zskBAaeTrUf3uUC9FDgyMM+luBV/GcM+w28gCENjR5oxtBNtuF6/WNyyyY34IEpk+ahaBo0m
6l4rG3meUHXkfiCVcMzDMXI42VNtA+BeSQ8eIqnA5it4H+9u2w4mml2RiinF8hQODoReUYK/7uoW
VyOe8DmfW9RGo+smCTnzqEMRBDt0/oacxHW73ElPKbDC954wr2Y4Vc2soNNnPomRQUYIdzugfDo/
P62vp43dSZ6oT0+DX4LNBXvFYKrVb2EbVcz+MaLAMZ+uSZNvm1oKYQgZ8sGkQd/tJ7DChoOfE6kz
z5GV6rPVCMs+VBQH2z2TP975+NauljK9uSQvX0YFE54eYf4NgBhyzYfM2Y/bjGXiN63opOALOSn5
FFNFmSuF6XDtL77+2Rn8LT8JqYK9MMTHBx9Txg8T00d/Fv4ipgX6ROHhCJP5Up7c1+BuH7MINzw6
7L5W9wxaC8E9Ave+BIGUI7IuqjSryPbivJjwmDafT+b4cTy+oPwtXUOsqSZy7m6jDui3jpCpn3Z6
L3kJbOzpnifkW7T6Wwv/lTcnlShBzDPgU614mQURNzBZM4WZduJ0hlIjLFTsh126LxHlcUPFfq8O
+zOaBHhybxcvV1b3cFPdIN4neoO32CIvnK4R78oWWiBNtOiMD3h3TwJImDWc7gAASlZDC1Ue18U/
Kb6euM430oyfK1vqyLZyhdWiQvRM3mXla1CVxWP5hLGeY/xh38mfNs1zPWtRwRrkZOqf9JhqCowO
3DohZoITtS+IFDYt5b8dfUvQzUlJzqi19BUoMGRSsJ4yHsPukH+LunQyvMO1xw9zcNuUtq0jSwD2
tzgndVZc2t86A8QUnFlzhj6Kx3dLxz2So0Sg2bENQJKwlEekuVCj289MtDBpKfjSROMcgvoOa1uL
2G/rGwg1QxCU9DgL3+dBUCQtTMoR7LO0bq8qtKF/Rd6fTOTAOKEQxdDWM7YIFzpRURqeQgrZHsKY
xbFc2DhII+NLnmBLILiS2Oytz1R530YfCJ/4sSKeMTU8uHxbeOcIpMF6/5zFjBA43xUE7ldPClPi
ve63zCvbfQaG4YWPNQdW2ZQTIZdZ9K6SluB4tPIQrkTCv/qax9fI/gIdB0+f0vxWSIej2vi22r7M
M41p0xbAG1QvvE48vsEKzcuyOKkbrws+7IDm3iEuNDuFbok7EgNotSHWuPXMxDgqgHl/YI1KnR6y
bc1p90c0II5KJgicFQEi7YNVYC/QTkei7+enzfgX3htLw82A2cEySv8YUtOVn7fRCKB+RIv0uI1V
f+HJHsGmlnvwiawm53jRvR8quoss5tSuYA5MCZrzwXs5bxWEZwSAomcdQlw444QoC149qoxYH0Ci
lC1lZE52tWOWFceOE5YMfum3/cTDqupjeuFO6BvKwTNaTjVd4BBZAhGyqLCTWL9CR5bdQb3Qay86
VMFPkCfgYPaD7tAmSZcrcRDDji6WHQnqtK1Z7XABFUYYKdw7AP172Yq670BLRCorHhlJ/BnFGuAo
mjMQlw49F6rZ+xLynljfcfS5e6CiNtTiXq5UOfvB0wZfUbnVQ8x0grooOkbQAyR97XLMOsOGTIbi
XBuHqSY4k2TeEwMMWxAZ/N0BcNe+BPYP4XlWebjJ3XO3D3e2g8V4cu/c1k+dIbgmHNB2Xk+TS3AX
PSaJJY91KNJopxBH+TtlUAj7RhM6XkYNomYw0P2EiSe5E1GTB+6EadmbwiEDp7qF4njAmwgg5IcP
YOij98553N9s7k8BXDFf0mmJcs3c67WiJMjI1I/6oRkqy4MjXZC48AHprxqH7kQ7AB7IEUbPaMYT
+8ZQ7UF1/AJqkc/6e6zfJMuvdIRZIEQC9RFbaq0re0ojlQZpCrJ7T6IaM4Cvh8DSg0p1J4oeBTAq
AR4syAVXHV9W27F8bCquX5fkV2uweGu0wlel589GrerUSbkIb0emEj5YB2DLqplCIsih3RIJ8QfN
fUDpGO3ghlPq71lFtMDcL9L3x0fhMsgT//tH37MpDkqKGrcBxnkUFfPUiSgXtNfyKrMvEccCHs7k
daBOWIgp/10+YOIZWtXHHBWGGRMAu9IRZE/UKrthZyaa8Glt7DrZY1Hmji2XZT1ul5//HkQpl9tR
MhW4bgNt/Rin7az4Qm/oDJ9cds1rl5YLaDSB7RrJmsqBcUddzAYDMhryLxUENCJCLICuuCVzJFbd
Vz24v9k42W0seLjAdsDer+sWpmv/tA4J0L5UbCC1JxLZZuuABKTLyBVXy6GEm6vBPIFKuVJQrZ6B
Wodrean/aIw9l8TDv29KuuvFy8BxpzG0i1+7BcQ7y1u7cT/MQAeWlmZykUVWkj261NrbcUnZCymg
snmoP0seMv6ny06z6ubRXDZhToqZrEAZD6XXiFY77qL0LKeauLc78l1+bX2afWTIKA+tP0HZgY0+
uOvVCZC4AIag3hz0A3sElFmCSHkg/mVEdCScFVAOQkpuzA1zHCWS31m90/0KDnXkUOoCEL7jxxz0
Bl6xpeZCBDTy+DGCw/p0qddXyU8phIYs03IOlTAaiZWXYgVYjY3aWMAvrsCyyO1FFw/wq6KkhpHX
F43JaQCqbzonIvi6E2mvKXccNjuqWspHgseqw5prwddsyX5pnWJ9fZVGI0WDOZneIiHDBKIVpUzP
hpKqT77ZJL+e7dgGlslJJvOl2gxGrlpZQoKmDw1kPFDMq2vHyHNP4YfFZ//qBF5gaXLqQMJvlAac
L0K2gMpqK+gEpWnX0rPp1Q/1plueHqmyOTCA+G5k+/x9uklhJ/kFetUyKdwEBroiJ9lpnaVHikvD
Nn8WvUuu0xylDUwobzYEDFgmFKSrDpMVzoQ3xa5cMqe+xqczs9kloajDXCsCRqo96DayvUtcfCrG
OGHVZ0mFx9DXxyc9Ah2qMBx29IDyVp8ynYj77/hNwQgIBsvM6ufVIvStULzYXUppUrqy8Xh+kE/V
SnAXz84mFVqcE+QBKwmtUyc7fGwpO7I1w1OcFZaZ8ahGGn6rVQ2BOP8W9eJdAcK9usLRfZP96DWw
ILKvqum3MHFWnzTZFE3KlGUrzasgmpRJaQwvw1XMcsYXRmX0TIRSXA/DkX9i1UXMHUiaHVmukm7k
CHZF+xRI9x7QnkpjUuxmicbdd6St7HYkFFyIllXbfw860PULhCaoRkoYqgpEahcJ1U/7qPDkvTBj
acD47XnLRIkUthEYi3xlO1RWhkKsH4rdxqmHYEnk32NQwHQDbFRNO+lPhxLb9hzJ9ZzrK9w2UwEP
ytt88s/VGEovcVe6dyHN3MzrJSjmazGwPPeik7y5KCrW/fhgxIX3ARcjt4SpBzW8po9QDGYVAUZD
2YaTuvSZ92ov+B3JZn+uirDnWffMOSocr+TrOcYsHCoi8CykE9LLnElp+1VxICs5TqvMtV4PuE1D
i3O/Xn28RMsrbkLFp9w1LofVb3qj6jmPX1llqY980t/JAZb5W0byVQv8ts/dV56+Qoy4QqD72IgW
qAz85zEC0Nvn5EPTXTq0fM143/emfZxwxyKwrCf58sQypNbGPgI0k9esXJJ6+n/BjUz0wzH4RzsY
XxBr/2OJrnjzcMOK5AFRN60AW2KfygPcEXCMFO+QOgMI5IJTvgq7/YDM5lQlZoHG6GIdjzgzKQmN
vckXNbavzOQHeQNkJ7cXHnM9zkeH3EqEtLrAKwl3cNWD8nD4T4/bVc6eGqlVXuSaq+8IeuPOPFW9
J+QqNBeXTCJFR0LE/WepC7T4sHEvoGKyzuZzdTe3rOvFvjIH+dOfFFBN8p39gcJkOgVoFJdNR30e
6jM0M+ew1or2WyQSjHbvz8zL2bHf6FsxyNKT5UgJLAOPCgY4MRWlg0x7oWmRQcU5mFsuy9vpU4Uf
j8xlxtx92P72AS88SioukwmaBS58YHx3Q2m3goMtKXHaiWcTErKf5STwRiBwjYYU+kRwTSqty6P+
NuVv3xUKUEoeTIyTTS5ojtO1/XifqR3j7tKaVUDhQ3vFsoenorepV+OQh2Tw/V5Y9c1IKxMjGg0q
sEQqw9oXXdpSAEk7dGR1Sa9f2nQtFf/elmgSTEfGtJlfXXKrX/yVk2miXhLtWnQCY9eQoCThFhju
mtxpCsBWapw1PN8dqaYHb1XDU4oa1NTjxSoJ495QA6C8nLRK4Tc4H50C5JDwl6Mky20X14HnEoR+
9C0pMcRsyqQ08fOIqHCYy+/GPK5lkOZgp6Z0IW1K5c/CLljs8gGF0d/cLFkgDR7qnYH4/rfSocYG
kSnYcQzdLL0S1oqy1ksXpuFnVN2/qe7eXmUy2doSg893f4l8I52uADb6SSPIAkr+NPVIgAcGcxGK
oVU8OJzDw175S7A55NLjPgHHB7tKV3v2bvLOMQbXy9My7QGMUXC6nIOU7I4XNhe1yw5iEYMQ9iNu
7j7w3+ekHQhxQUuLLv1su3Uk0ZsvtEB7gCvkJxr1XVzVk0r9fSUbFYTNAr+TBIcS26dqnxjR2+Rj
aycScEwzj4YfD8/t4Q5ykO+z/bNOIfHYOhF15o/4xLj5bi81pgEkSG3Jk6PSdc4Oe1mpW2RvkJIZ
liC+Qg3sc0lMwX30JfLldyVzYniMl9ksJlXgtNtvbnbHXkea5VJb8jJlCLwChfDO2G+x1/MUUZC0
avBiXSksHcjq4hQvmKat64n7a1XArJnnP9Ftzo7NVt+kz6OdWcKnu76uEpp4PhlG5yVRm7Ic4Ptm
6bafQyTVV3mRAFpi5S5w6jrzQH9nha/YcFmuX+FFJ0OZ3020vSxah3ifdIl7D5+veN4ByK9rc62M
4Y0uw+qTdYtqLKSvjOZHOG1ruc/yA8SCYMmdiOgIhaBtFxnpsJN+5q8Xif6oASUxXPRHUOmyIfL8
FfTnOLfgZ72XYR8w9+G9xPx0RkfU7g8W2gqR4RvznhrTHcyE+MGhkYrTHUEYoUmH4GUVtqeUoEdu
ib4ANNCWwFq95X4fxhJ0Bhd/tctxvKSOQoJTmoSLSy8fxOjdKAFGkT3L3QQQQlJKvZ2hB2lHE0QT
LcnvSEnkHPkDlbyDHEbUXczbHG3yY0Xr57RmWzteuwarGzhJBQV5WGQfwVCmg/Irt6Udb+4ln37K
1fARsjNWM3Cg/JUUQ5yXY5c4Xg9z2+Dx86o9z98KPGd5aILjmql4yXKsiXI1xDHiemx8MvcFzTSA
mccACGCjBtfFt/aYGb9CBtFAq0DT8aKJntmdcex3bgDcIsHA9kXOJmBf5HvxNN5TvAnVOAsyLDzR
kVTvNg/GA2RM4b/4ZVjMsD0smjHo1roCNO0yWomkw/t8cpeKs5EfS3F/Szv0/uUt9a72fgzFP10k
2JO+9JrAxS0ttp3GqiAgBj1o3SfZxqGJmZ4z92Vf7motnbI4CPPrjdHmmCVfCaYnLExOe+2udu9/
8F2Fif3SC5rqiJlEMFeNndT9nLg5XygO3Dadf7ejl7GRm0pEFYSCJVjvOn1nFzITkWvieX75Zcma
iN7eb4elQ3XfQOrhseHEIl+FZ+EZjO+ZK54n88PhQC0hzPx97vaYR09p5ETVuZaWMbij73h22dwc
VHVcvvxg4iNgldKAh3o0HlRF1sMRCPUkgKRjUGqb/vy7tEqv4UA0KjxII7Ad3SkuElr3FqEYOlhv
PA3p4Oo5n0j1sJyTyzZ2cOtiE1EuBGJySzAi+Fwwc0F5HaNJhCn8LIHHbW7RNI/uPzyRBe8F1dUp
pNd+mwHyqaQvE60supqia02d3j7+3bXU/y3dZ+QvJNeP9JR7IBDBthNwImKwam5TW1aKBRA3xt1b
Xl3HqaEQ5ajB89BPXCuXg3z5CstPZYKzNS9/dkVj8wjPvrOnCCUNtId0lPptnX3gzoba358gMi2l
Tx1ULajKS+dakGjHsaOFh2xBUMSsuyzLggKmlDYQmqK1nzcmVLp897VN6U152vVXpqnkCxK4oibX
Ij79NH/lChcoPYEkgEJPCUsEOzC513P18khNgXeKaSNYqZq1268LJl7DK0Bt32PZy+2FGzcY+3Dr
4iIwueHNZEk+BptLY9PNbpyJjoJ8fyLeIrfHpHrXmlsrz0ROJqk0Q/krpzHwX8Ahn0v+3TRQ2Csv
0siyYk3+g8K/Xaw1Xm+3Xz0oUBVugKyo3i1CtteGWkHwKO+rdCKyxKFMmEYv5xv88VQLXdJYc8De
cou4GnN3zvSkv+Ixg7JFOanPVEMLfy/7+YBwJAAtVb3uyQluo33kUhgjslHbHJOf6qlmYCTgfEvB
ifuroJ3vdFrGWMP7b7IF3TXnq9pgOuBaYro8tnnCwRUiQ+9eDeum78/tIXDxx268y/qeetaUGpfC
u+P82/dN8oDAit9N34cxpHs+I3L+6ZrEZ3zuxYVxPj3ouJ8CyBwtQnRj6kXDyOkCi8vFGIxsJXKW
MVKun6Tf5yOOxTEXK9JEi5ehWKuKVvQR9NXBefkDiyXwAcL4ajsiP1PjFagxpPLpAqIvJeNnFAU7
e6tpr/3YHQF+s6DjQptOd8Qa07E7+zY+V5+Rz7ih+ZgSR2iv+T9PbbO2dgOWIwpYknuilWSTC1pr
WynIbJgVGi1p2BBqvXadfmKRUl+69B4eWYp9WWON03kfiTYjgz2jpx9MGuOQDoQlhYscWa/2BeY7
LaGJNMlv2T8GUwm72QnCwm0VPAUz0z3oHHtAyjL5maJdfJQca1qcQOMRfAgtpObTVVWjZP2OW0Dj
6bFcymSqOwIJd5Td/y50ea64nJhJH5pA6gQIYHlrRQSOJmbO8zSZzqWWUBVeuqa/kVgKVvO4ACDw
M2PpRl3zaQROspKLqd6XuAAbCc9+N6DBIV24n6ZiIlG9bQzsFpaLw0eYDD+5i9UhCR/3ywFtoJTi
4OXiu7nDJTCBq6VzUxBdt85DrWixMf8wB/uyJ9YmkJM3EKaUjVu64aktCmdFMg6pvRRnkaZ9jqEU
zIDxVX1G9aJ7yQcIruYeqMSoCyB8Nqqdo6hFKuFq2VjZ5kabqXancnRu2PcJv2VgD3IxvjCZrEyx
uKDrxSz1jwjscWdWSGvq5oPV+hL6NfnAt65VWqPhYSE3u3kVN85OfoYqL1Wo5rq13rqM29jX6RMy
rSmLzI0SpUvo+N8mD/qH48+gzPF8RBrVDSMhzbCcHGwg0GFrNSWIAYGFqfGhvvCkXFGyr6p0wkNU
1rluRDGTyqS9L7+2WZrr9qdHDpmcdl37DRkUjRDs95xKmvDXv/+EhS1mhYoN9+e113fggzErIdM7
/G3/4yfH1MHG091Zvm2p4fyLYX9yMjCGcvWyUlIi93B6RQKwtgBUfMPQOf5Am8KztZ5RzOk1d7y7
6DDqXllxSW8iMtTPf3jtOgOnx8FwnLY4lovurwi0d6P1pvYOPK+YpEoqSslvBqeQB2yqsw1rLeDk
IIbgHo6ePFKWeQdBA406fGvdJAviVxeUMCVYFdjUkXKKsJR0C9ewm/YiYU7hjwHM2Y/YraYHnHYF
pzqrVILH+p7YfAc+80Wc6t0WyypulHqenEyqRKkJaoMA34mPRZHVahqQ6kM5tYBnrntFyh50Y9Nz
8xQo9q5GijQn+0Abq1xSxpxdF1lOR67bx6Beb+cxX3JpGFgN6+fuD8LVdFGKDN33abm1fYMLrSs7
nocc9DMgr861JNhXhxM1yGD9Lk/LWXPR9TcIFqPlpI5g5qH/oUBVLTKQcrtMUP+LPAl8DMmbogUl
8ojg4Qk4hBqCoKDGw4Fw7crl33ERhSYDU3/mUM3Q2bGCtp0tRqLQwFMXLsn53l6rkVrKZcsgPadW
e/W+0cnPeZlwJGvlqp/xnR3vzLItdud+uby9YsQ9n/S5PCEPeKyxPNu2aOhlcjIF4PCjG4qn7g8w
p0CftOCexLRBekIw+Ixb5jVLw1UcoAmVUWyFhstXRTJAeSdYBQtU74qCEJED6BpnGLxeti9hBGnQ
5PPjBV2X/EoqsQDaUdNgWhFPeroLRVLnXTOKEmBU+6w1UwB9C/HV0g+Dld4YeoY3AaBIEgLsqVXF
1uRKRmXC/3FdFXNcQNmKV3JQXbNa9BtNPAJJ6OM0HnxO5TmJBfuKuiXTreQZkvqPMkEiw89FQ/ix
3voNPs1zmk+ggQNu/8W0BWVevfTUy2I1XKjIqQtw8oJWvKbkaeCxxvvM+Y+nZIqWVHSlQun/0iNf
zc+tGzJO5Z9FpXwvsheGu/DpR4LQ4Iohfabng8pJsyI/bqfgh/LP/HDGrCA2E0mEYUZOaIc2qMMo
uIrlqz6dS59g2J1RqkHwxYU+3LH8RBKKHi4MxXnw0g8wPTOUFG8duk7kBAplIRQ7hts/QkKAd7HT
h6kpJ2jE8p/aUp0AHCbTaye+W1qTfbfwz0ASesZqp+btXlCqE+wS4mHlzixsljy/a1/XQn+IdVtk
uqq4RqhIf8KbY0TPvu4Zt+jBOOPMmUnqVy/5FCvVQp0BQtTeePXiPTJOBFfb1EHzkus5L6703Tw+
Bbz7Jx5DNaYOAMoCxdqla69Lq8lgCQcqYpuCFFDpyPg3trb3mphNROKjqkHgAywuBxokTthf4h92
SsKAPrOi7zQvRETq4v35JIPloA358KDpYLpi/j6O2MyFACXVovG3SMsbxwk5NVEsSRyNjQ159H6Q
sVW1St5l4slHfbnpRfC+R6QY1GArX8LemAhmnXp0SWrg8B3PyNb6YPKFgqIZInBSw74MvNar3qmf
zLYDmv7z8uKjQvgX0wRelUxXi3g7W4ThMhjauGUpRFB7Q2NmNTcrDLhB7XNYyQnZrCngY/Pw8xV3
ByQwLP/uki6RPFgzPj0lE/D+wSXDdOHnbcMzqayLAQTA2IWdZWpY6ja5o7jJNyIhPXXu1rLu++7N
Es9+GyGW+5qphk+z36IFAUxdAC9yK4voBrcpY5na8WlD+fRaufHL44YLIyxsEJVyIn5nzynZ8/8z
A9Jl5ww/J8eYI+m46AGyXnkkKU3/KMADCKekMm+KfgIYoXnQkN+PZ+WNdLHzHZ9Ro+l2jayhSAnG
+XMrzpCrhQ4uUm1+rkpNcDFMLKevOmEDCcQeQPBfLy2yB9iQTxNv/2FpDRC1u5uOIDAV52Lh+4tG
17uxFwzK1guf+QoujBRNrx5EWswCG39DdXTNrUy+maGelmp99QECbICeuY5fvF53V4wj6Ez+HgS4
gsDKWw399U+eLcBC1ewVwRtSpe470T/m+ygAGqYsyy64iUhRhuzt/7B3PA2Cm+jGy7pKwUkhJPxu
daiwOo5S1Um+UpDBnoOaE9JA/A6JTl0mlSnclJGQAE5YTk/W8UFYvtaJ3jZW0UkxagtAFWn1ieVN
LuCJAljoUcywp2ugdZVVFsdrl7m8OXZ4bTE0XrnFbZMae2I6RL30Fuk4A2RFQUy5q80KCj079NjT
AtCUjMZ166tMMwmUGS/NL9MPVkffp28hXJxq459T5yzIVGR/7Gn5zhI+yPbZDozgmKTy5XnV/F/Z
v4vsX/a4Ph2OfUNIavNb1I2S8dPz8LZ3Oh9QssGumFRObDXq0PGyLRLFAxTBxsyBVa6eGTG3LEt1
4RGz3w7wmEZtgC2ET4TR3wDxhSEUHpDaHdTc1kFPELh9om9ZYhLo25gtMzptNk7BlYQNg9M8QqXh
NVwGFOc3olmk/8rrXRAq9Ez7nRPONa0drTXL8bMraQS8diVW6ggDwzpX9e+0vRlmZg/uuYGazb5a
baN2v0aPfM3ke4z7cSujwYaosBQnODU6qIUe+udzDmG2kZEo3gf9GsOqAC7m1zDxb1gBYZ0nZ3Ph
iYyPbOQxrqKp9a02WDVqqAo3R76iw27eDT5n2s804exfgPPtUz4wfZMeofHehBD4teckdlhvnEEx
ONdb9TN6xQ9AM5GrLkL6Q+FjhMh/Akz/Gl6/dayRcU+54/UbVOOoR6QUcHwET+zjnyHnNhKoT7JA
oqIYh4r97mkWDR6R3DtsDuuc1STPpEX2EQyqDxorqDZtgK+Gizcd+R9jZnHOiKkjOc/hxQc5gOPa
GNYMTyqZdPx3kYD+OA4HZALvj9xE5Kc3ktsV/SRkAp1LcPXMlBhCTnnQoSVK1JLGo3AXI9Y/XfkQ
FvUYNYEcMKDw0CrGyckx7CEtwllN+/mXr4gPy1n+nsCiXd9VlujRv/YQuXMlSE8EfFhZ5/L0g//v
AJtEQUUUKQds6jV3b5pN4ck2Mff/Usl6P3SWLDd6q2SowaUN8xELzAcpfgRc4hzLIxJQfk6N1n2K
TpO/mYaxdWj3JEb7nyC7zuwNHAfHMBamfWJUW8xQGq5vdwuRgBTZc//lPejE5kkY0/+drlVmIaPl
ATQlmt1m3uRL7/Qj5Sg4L7w/QkiTw/4smEFleQ1LnrRZOpzaVYJK2Uv6B031YbQWMNXlSy5uBS5p
uoGYfV7HxfaauW4OPxbnH/TpfhL3VoSZJmKpmcDb1GKm8aEGOT7JNqP844e4imZhhIyAcoKZdV8V
AWRfdqaSeo/CkUGrOx/f0RdSD04XTkGGQeg5JfYZwuqJwOIXyH9oEVxyWnChphOZOeTW8ZSndjCY
bWP+T6uQgR8uWrtvUIVIud/VJ4F7cesq75rcRsasNuHtD8JqPu2rXIOtHS1Wz/5nYkLv+3gRSBi4
jFzkrVFnD7GhQmTDf+lkw2hqjjnpszUlrXBykMWvVgvj3P+vLR55mJpKMbugA9ZdhxfeViKnEkSY
HDdRmJX9W2DV7mranZn5ejJ1AODcmMngikxhmriGZE1tTWqcd1cL2cLGXHk6TPKY8TGGUyyEanKR
/ZoEfr6kHc7hC7LEhTjPQt9vIFBYCfdHxuqANHyqCBovZkX6Atm1IlTCAbo6aAIwqCVsNDi1vUDp
dS/Noyow5OX26o+zu6HDPw6FwLngFR9cxI5c3F47uHf9ieN8QaF9jKCOXm64jzBE2nLK8cO2n1BR
EJhf4m465eDimLIl6GECr3aO/nghaR23hAFrPrfucYgQrxccVMJjsFme1KsNcZ0dE72ronOVnHx/
Ic2ZQ7ZiwN9jYl9U+/KoK39P808BfkwA+SGUv6Hl99yAMGcGREgOFoSsH1hbhZPSencG8bnorEhq
E8gNMZhbEB0pg3jjUSRKd1S23ua6VLL8R8EL9mYtqyuc9DVMt544U4cM06+y41WWjLVcxDYil7rF
X6/dxz24jAPldcf75ejAVrAYS0pB8/mHCPCog3WocN4RJEFttUY/maWpYWl/SSShbJolBAGhFfaz
Xy6Ms+eWfscSlLSGLG66YkjBgDt5odOsyYR8pYuF0A/XP4M/o6nviS/jsRvDWXF0BOd35vkMGRUV
+7F2ZcMbElPOMRgMMemkwBkWDLQiRt80nL7QkhUVEpZyjPvUqYo3bR86Udq55vYKN4+skfjyPlmX
yje9FYywYjlzeKlqv79h2mpCbnc1Hopf7vifqnTLhJ7ukYe81mbtRwtE0lnBdp3GpdzKEkDJmvyI
19z0Lf1zLo2IuI++flGL1xt/pPzBnanz/jBC8vFW9OnJYVzvVHMZbt2PdPKZqC/OR7blmgTVpi4j
mdHgxXJFVDrMys4VGeJSXU4tQWvnPBg5smCx5zHV0dhnLWrxekkTReathuqE2+q1OaPLmkRKMe0L
aLK9DRpd6icxC2ZUxuRhoSAPpgezlEmTF2qM0WJ4+McIL29rmXs1gf8yKICqfaNvZaAiFdFwl/xU
91p3dIa8mVZH8CI3O2c9ZBfCIyrzrimZ+X6FzINzH/E67wKTuJdj8emd/13LGJ4gZIp6q10yV+4m
VbCj0stfRDOx+fHksO47o3NB+E7WYrltiM/KsDF4RFgDZisEasU3+tlEVW/cJjnEuVDmwLi4Ve0q
3AT8qHo8oIflvTV9gvRpxehw5Y+cQAdVU1+Uds0yjgDahrjUeTUbAlSQKQi/Jue/i972y9lF/tB3
DbXmXYyI41RwYfou9qjU2RHFe10jobgvcevcdRk6JXgoUkV5tStcmVSmZ8vDXfvq4WUELK+a86V/
Av1EXqLkkUUt4hCVYiny2aFV3HY9/tSHgvlxhBOONmaMC0QERaVOfBzSxl+RU9dXyfNkTcRcLRjr
sGmKLOoXvv+kSiuLJh0cZgrbzkCyGjJzfigCJi8oTxhAo5HuD8tF18rH+aNfnE3pJIkt8nHoUhdz
WdwIKMofoA7Mc5KpUfWfW4loErru5kxJI7jUIt6STGhx06fSZeQKq4+c0RybtTx51D5C2C++G8pT
oitptwJsya2o5BiDwfLJISTrG/bBQuvxGm3cVhT++6fqfKNbZswjI4OwEKWlsgoXmgnxCuGlQkji
CkPle1iUQkxL2AW0wFY5DYfbPJ9HuR2nkClD99pJu1Wu+Diln63O2JB+jykZVphZBMfgkfLoznmC
8bejp2AHRf14LDKO+6FH4iP7wHOz0c81yN/0JgQTadTp6mTI7joj4zZago5A3xy+hWEdwwv7MhI7
MPgDLVLvq3QZ8suUd2BYrmKeJxibEa6Rwn9PGarIYsdos4y4jqojEvc3a5/y6/irkZ0XoKsS2WRI
38LrFIgz3dwyjTgTH88yCy/qBv0X4r6qGXC+7ahTT2x1vXO0Y8Y9v0uPatc/D0yq4ubCM4wzbdZO
PEfXdKZy0CJmpej80M6XOCGU8087wOjw5vCB3kdph2SNuWKX3RImvHFrv9RgnALQUwYvkNPzNfsW
RtUVNHZ21WMU+Qf825NoRinDVJSu2vRki/78zKiv7a4AAUUi604cpvpcg8cGNyJQqrvs0LhNS8cM
bObQ4khvH6jx+yFwpBeGnMyACn5LhGD/OE3GI86M0DD1rBTjRWGkgCtwbNH0Dd0/OerP1SDamoIC
6xZm/ZXT7Lc+hP0UT9t9t4SgitYCjhBGrRLOMgNv1l0Bh91EDAnooaOxs0c/gu9qUqwQFvLT0Nr3
ba/LYqoNHrwP3TBV2WDn8/i2E9Oy7dkq4lEOwYzTEUuFAILuIrMVU25DG9T8IJ3+lqMhIy6JAYvi
3fERtyuvcRqVUNzja1cyMcYkD4g+OUqirXYgejOoy6d1tX5KCe1Ntwy4gkdnm1kKwJRkapEw6Vrv
Xr+rfdd1SBNMVaOfPokzeVG73fxoTokvEnhlVAV1sqYQKwyVHo9jEMUzZAxqGZRZ32p9Ai3NKla7
G9KUh7QaxNwIe33w3sDvFICe0c78gqySs7GXmMeAR3K/b6YdLSPohmcYgdYoYVP+OijIdJFdWyqs
wizXyjKyMIL4D0aeORpF/8MYUzktKEJ+bUOnBEDsRLiTwg5kRzhmU/koDEcEKjFNgCD66jLlycWR
/rMKAaCyLfz0/YrrkbIs5NG4bXwOIJeJXtUwO3pnqrhoS9KOKSZw7KIynNWeF35EpaQRQOGsOa0n
S+D1lwl/5mmj3pE4oCKCS4hnpjwz9TIAw2baawtovTAwC0lqsD8nAfko7n5n7BmgsmzvuQBANmFY
HBethGedZ8+O/DIbSL42VB8Hzyccd/NKRul52DZvu/C69x9kF2Eu0Lq+eoNOVYYWqy/0vK+HObEU
8mZB/MztsB170mZtl8zZ7m8tMk/JNKr/hbDVUnY+Oy1MB41NtKjqC/Le+1a1lXpxYE8CYDNyb4Ow
4UyjpBUcy/zZtkXtAB1a86fptgJVDqeBGG/YIsDu8cnGEh1LCNlHTsmKiqtqDF0pYuH52AQCOiFF
ZasnBMRafWg5Kwsmwtv3DGpAxi6/GMc79cyEFdpkry3bUQPaxLonpUO8Vm3swfMtO5wO7xRZWjH0
EvUCcYzrLQLVi5H55taUFGhlkAP34COvbAb6T4rgFbTxAaYysgo8hSx6eqsnXl7bj0Q/dV9cqAwg
etE2h0sa7VeTjj4IyA063E0GenlQaRS+55gWmYqyUUYTyF/ELc807ffEWpx2/9Lff79U9R/+oXRK
JMFA0yoMKdqiVeHQPqvvOAdsTsLM/OzkkoKl6qivZWxS24dxCDJs3TEZyKucWJZEeSL/Cfr2IDOJ
g5iyp6P1uX8UDf+eNGRxqD9Bcdoop9HJqhxUThFMWXLffa7pBZRwQ1YH/IdDWg5wLlzO4XUiOhoa
aQ7jCjX/Rjhb3+/IqvWkrXbNWzlRS9102wu/htkg+GOWIZkpF8BN30Q6sBmJsVxsd5dpgD5mtW2I
GwXIArdALyJZP4QZQf9ahF4xxC2DO+rCnES+RNgWt9YehIeDJqvcAmBrxLZNkzWE4CKerruWJoSh
iy2a/DsGNdUuBRatmZLh/qtbPWqFosbsBAfzH2F6hsnsyRSl2/8XW7n8esQ2bfTdBVeFHP8LgB89
wNtG/KYl/g24gaKv9RNI2yclLpPLf6dtWul9dvZJ8NvV1WvDWEg6CbgVfwFfmu2ds09mO82Tht07
0JB0PO815FZ+YTClptXlT3hAGaVO09hfAJTd6PH/q0rtSGCU4WCkKL/Mg8HM3ybsH6CEhoZnAThf
gRjwY34owHV+PtGxu8oPHKQ6fKCMEogFIIhWfkcGBXzO8o9hxaHGIWwd+KSsPR1fkGdgpTz7sO8G
fzG4tRR7NU/mJxxbGEf/e2PwtuTNe7q+aP2kRQKlS66xW5gAva5swcEAIM2ClX8lZxExQmY3pCty
ZzrYtrOcJeZiy6ICSRUfAOWMLMDTctBaEnCpECPpy9QPkMXHgjtIuQzgRtIrweNJIFMRZvrxN+mz
1aOY0yhe/7mecuUvf8Wo+yeDN0GmxAFayrFewnUaBoNmxV/lUVoCHK9KzCkzlmyLXYwUWh695rld
aDHceivjsMpV+W41b4d31yXo05bkGI0nks2+v2kd16o9L5G+PYa0RqPJnXpUdTp9r5JZvkBZubAl
tj0pbmBUVjnRpUFDkpXDIV4SFdp2wLxDru/wJ1i1y/AHMHF1g3QLf2o6msKVP30VCgKvB0dPv+ev
udqQySeIJIQYpdR+A/5NLRYm4wbMsLbfp5Ju3j1+cOZPZOBMUFZdm5XRuW8nK6CWg1EcPqb6yzQv
oHlkobVu5tnsA6EjhkNd3UeydX5iAiLGPH8lIxvIy3I8+gzqaFgWc6jtkMnNFPlsERZY3N62zwDK
87FJO9dipSpu8RkXQnoF0t5/czFpoCTMabC7hGBzgEo0VsFwH59jxAW6aDpdQXiKOMG9inYOT6is
/zg6/NQYQUKQt9X2ZtrQeYN/NyDHbohLJX7BrVofcITTqwebLqtAu2PVM+Jlj8RAo84/2nhhrvXK
8pG/gDtVrOyZKa7ateDIH4dQ8rmmfjrfJy9/4Ml7plIBBWM2vWC0uS/t/M/I7T82l1NJ4CfbL5ET
8xDOnJrXv0wwGCY6PTKwEuC51TDglqB8pslDWuf0w3IpTChny3hS9gMUTxD+qUSM24fdAR4prcES
WrcYNVhmWFnzLXW4y8k/mRTW6dkOHzMH6OBf2oXXDXfswlwn0R3rI01QkWdUe1qcizAC5QsZHcgX
qPJADtd9xeXqPNfhWBnXOSH17z/aQYgl0+xdHml3l/tyENez4Q7tiR/+6MGIUubUKu+4MkTnROFH
VVE3gu3kUspoQCgv/zV0851TrGBYK0r1Usa91Awlt0xdTuI5OoW+SQPXBJxsynS7/OCOBC5lkBTn
yM8s8E0zLmkQ4h5ExUXCjbgqRAUrjeCC09tR9lrbgtFT2QZ7w3Bi+SDmvEx1IEKWnYDRtVd2V6qF
giyvg/tP/jIp3a4l9FdvL+A23tSee7awQvDUD2n07yVCSy+ATZiJ867JIAFAQ9z8vj28UfrwTuVT
dzrMXoNUURnMmxxSp2eT6YDZU5bYaiDykN1ic+ARg094Im4hEONFv9ra6PRMJ++Fn7JErJHHlWZe
7fSQ13Xp4Zh6wxEA4Ea+N9dAQw+hm88HGv3Sv2ba+kcjUcinZUDrH+l3ytbzj/D53n94gm6ULohD
B3cWyk7QuDJawxA6TH2WtVEJDzOs9MgrypxNKDcEoL1k8ducltckCeOnew8Z1/nGMzg0WrY9tp86
3D3Af23ev8OFyitgdyPoP1zCg8hEYj0TPR0vwfWEROs1XF0n20E+acsdhjj00CeUX/syRTzz8sOC
rZQhaMTCBgMh0d0zqiPNh6jEErsHGDyZjk7elDqBzMrtCxxokexrEeJUimUUX+efQlC7US7EkDd6
lP6a1dRf+Jz7AvfT7AUh88ZrWeayGl0kPK7hQUol1UHe4otzFuK4HBQ8xV6aPC+B+xBVgzWYcdNa
BUE1UXEJw36DvH3H4X1vjs2Fp5scNfdd7v2ceGRTNyy2Y/lCynochDMEdWdOWhtEKjwuYC5Bf+S4
eXIJEdSZB0rHn1I07IQCHVNKJYEI8QTjcIrVFZKz9lp568tuLj1vuTNAboVCL4qD4P1zlN801mo/
6v5IzDPPrIpvBbM8Od+0R/5bwvaIKRKtBM3wAXGguHafg8N6OJe7dcQsBogUzAKXZE4Qnw5NMUkl
wkKlqmws+Us+AtZIr+br8cWJqRBSEWAllmqdcQv/SzbLz7k9PDFXdIUvsQvph8nsy5fOD6ruyXg0
wx2G+aVu/RIdzlbtk/aO8r/XbYppfLRk7TlAqcgb5fJH/tLSV5B+8hpXwmVnSvFSRFloWMywGOTj
UVehUFLz98VFWKHv/iOoRap6ocJIqixT6zwPk4KYXi+yEgtvmiCEbD3xfQQqfOxbzv14P1J7UNI3
GhMySkDG70HK0WGEN+K88ATq8AoFLrztACXcVXBwBvYiEbt+wtziuQCbU6EBa6FGndCoESzY+mPT
76Yg/vmzxrHPcZAaeqFWy1gwpb2LQieSNJ7vXLa9IemOow2RuycgRsiRT0DMKCaywSOOzn54tkgy
dQuQjroL8KLDo3kUV8/wq1epC1hz2bEaEjHlvXKbHrnN2kJmmVsgCI/1f2rDPxrTKEXSIc7WdvGt
BdAYvXsGnwOnAN/+odiwbuMeqs0dtC974aoo3ctNM/OIYHhhwiW6F+7caWsOXTgHm5O2IfuLo/lT
HGdED4Dyx6YgRPpCTEBM/jIZ6K31jlgWYQSfJdlgkFX3cVLB/6VN/sfuY+v3CiaOQLLD9TSx0GRx
V+H2u/GUx5qnaAwMbSkkRsreRP3VyJkjD18MueaiBj+ZwSb5ICIDZGBzm8jgI4HJ34SE7EPuRjVT
zZICAAZEjgyF0CfL59itWEGUMTtSTwwVkB7GoioYfNh6+bm288KWaX+oLqssFlOpzPO8sDDH2bg3
sEjvSvl71AWHnDAThym5k8i5MVHyYqJ2aStYvVuzmkYdABAnMcHG6kVTkn57t64SgXMXNBhgWubA
qckt0Yjlr/0Kv7RY859IJgTkPj1PYfbPfHQCM7bmjz+t+Tj9tZQ4NoJUQ1GQ71YxbKy51bVzRfsg
RnU5jtsjfiKzGjhZmSvSdWkS0ElPjVOXuISMUKCckUng8uXWtgrnc8ynzVLb1NzftVao5BTq+v45
rliDHoh89D0qHgQNJfy2w7/qH0kOmcgi4a8IKO5qgN7w+wOJYnaMAZSnwA7j7FCaK1kWtZiATNLh
DMj4nDDFMGVZXYry6uD6Uire1JVO+QFugitkcEiqZ5TciiK6KtAm33XEe5j53Vwb8OM0PiMNcfWH
Pc+pmmgzE6G48dqXY191mR6loM0y16AZrg2GU7MUDYHCsbEIw3bQdbuRmw4OesLzntszUXtW86DS
fw67aemTHo6lxXC5IV4fDj5XkM8zsQOqUaBkANJjtSSUwTCNUSsatx65LCsXBd4Ek33ny5fp8xKl
UNXmS9iL2gFkZjmxNCfhTjGaXhhomTs5W9a9sj0ZoK6ojvZ1uRDWUNn+hO9GeGPDhrUlYGtpM4xv
/D7SDN+Tj97UQ8r1Bhx4XZdkEGZtQlaSabMuYGNBcPl/6FhVqeAqGabVCmHcp1u8DFSv06Bcnt2K
FHb1Mly6NE+enlgDoYetm3bTIsgKHtT+U7VmA0+w3zc13aH+RQhctSYe//HgyeBI418xBZnb/SJz
2RrGYkgisMw2rDgZ0NiHdEDfkNAfUccZuKkbw8J1qrRMZC3WvvSApQBviDK5Zjefq8IsdOFCnlE5
ROTKM0jwdEzKkgsZ6A90poqaBvaP65Src6Po0hBO3wa+ds3ShCjlomdFNjlcpD5ACb9mNInQUtL6
r5illnRKojvnCuG42dIQ8vUjyAr6CKwGRQj8/mVLx+sQLTZ2wfrxNTw9a7CGo34YHp9kFVaDhwnH
GzhWGI9hzZ8eGFTRdWY0PcSN+0ZQBb+VaTE3XIGOwSvJDux0l/nhb6mTK0DF4A9aEUUqJRd0yPq9
0QTN4/3AHg2zEy5d143goteH/iiV5rVaZGJoC+QN1GRRhOAZbZVM5BnqIL8btz6mB4AQSjr02edS
F2VhIH2VUvjAA3d8axSYzeScExnm+fy+F0rrywuYpqVpzDsqR7gOclmRZZ56nNrMW5fvDCqEDSTY
6Y7hLY8brSa/WHU7ztbX6XXTbwlQTPeRAENKzkdqC2hcxVqZ39Z7Hvyu/aWil1hkKnENkXenpxsk
0NjN+UqLhAN8yYf98QNN7xkJ82sdddxt2vOSj1qEllX2sguETPAEVm1UAXcDfm0i5uCq9qqcJRzH
Bf/d2oUNU9fZwsizCPItsBZYb//ZEaewS9wYDo8HJSyIUNYM7a6wAP97+ftFBL9i3bhcDTgbH2YQ
WxqUMKqvWQVxgb6028yZ7OMnjUlgDwWTeQsraXKJZTQ+e/r6FGihlPlGTZGOQ9HBTYfSuTgQa85m
FpOTL6rUWPhOoE3An7s3R+0iAxApCk8iBy6MLg8l2NbRVsoZ9FsLFAnHiG87snxde7bWqJsBx/nR
YqUm45Agy4uQ+2+zsI+HuJMQVuYJxpMFoNSqhhUBf0lrswDqUPcLrvY2/E1JPMLJ2Q1MR278rwfr
W2pAtGEdBWnLsadEOiacCIbFvfD6DCtP5+oIZcDJ/1qh5l2MSkWuAOr5JJ/JSaTVKH6azxQ3WLJL
AQyg7MgYcBXU7Bt5bsVJ9oiUIL4B2kzXxeTDMfP9vcyBHDxoKAyELShkgV9gHYeFazg4DTcplEJ7
mYUiD5wgLK7Sd9s3K4Rr/xJCRM7KTvlJgzlPQvYIteOk88mzKC8WGerb38u5zLGEEzlhvqomE+4I
/Azs6p8TR/7bfdL8sMYwpDdMy7Ws3tj8dkwyBlDP7f/y7an8KJES9v509j228A3ZTSdYNsxgw0tu
XHC06hOAYwq6zBcrLyUEK4E9sdUPfhA1xXKKW1i3/H6vkAFLQwvSZfVSHAutDIrNS3y99v6yVwvr
1HfAxamKm2PMT4EhWI6efk7yAA990R68BwO7Hq+/CkXLATn+hIFRkLG9JO/8cJTHxySMOwmmf9t4
/EVvei9cFDN1aZhXLZMh809Z+ETQiZZpdwmHxrSrCN+0Rlb1WRbHKI1soaDCuXLbY4XbVlOVv+rO
H8qsFLaxY7p/V87Fqj5cfG5UKkL+8c10QxLcIeWMNh9UwuTGdObhk/zO+MPBPVP2zDf/xtlmU6jg
MmF378xv1WA4QtTWSX20qWa18yRIJb0TqlHfeaLRzYFWIxY5X2O/qJFlgC4Q99756m0EL4vdVtci
T5Nx/ftqcA7Sgu+OwAu1QQBwcvYgi0tWbA8OzZ5TTpdyVqqeVhktu2RofKonFtagRRiZOq+ojK5R
3aQxH72kkeDga37DNR/OpKzYiRwpJzWPhOl5OiIW8N4+L+0/oRalLPQFfYzjmuhFFCHMSyYjRpKJ
sJDVM0P7foRLHGlzOGO6hsQouCAxKzidS5wJTEzF1wiF8Xav7XjvBo37rgjM0z8IvgenbhoFrZvP
GvbMsGbcwoD5/+2G97TKDBLoC8FEWXufICDr2dCZ8PFYkrOITDaZ73S+5APxdg40lRfGiQYUEp/N
Mmxh0yzUn9gIGlpy4wryxe8tB/teBAJOLZ09yizNgDMF/T+x+Pw9TniW0UHsA3NEppVBtBu1/GWE
y7ZB05Qc/c3l5NqL6/1xYxyb6efl+zXkaCB/xnuH838yV3u5lRuh6Dg98gyC6ACFRZNEevDQSzLO
RGFX5BFc3MiYLYV13J67nLTJkWDx7uaU8QLvNzB6EcdwT3Is78SnSTi8eOcdof4KelntaX2HQTYO
uAqsliXVOKlCj2jC1YNHcatYUQ4wBNiu5mHLNgjEVlRMwNUwEqsPLrS4f2IRzpqft68KIKLssoRb
kIgzr7Tgy2LPEOSFniilZtNninzsEUpJ3iIEZS/AyDrtff0YIEwUEIde81BxasmwgDXoeuXbNDnN
bzgx5V+xcF+kPPUa0nTc2WJISrH3QKnbjlK90y8Ybda0H9LFLo3XpGw/nXS5f7qzHpnVzrA4igWW
NZPJwrI8TdD5ihZnxtCMZmzW4JC0hmCxnRlHlnXrOG7v+ankOcaLqnbCOwpju1QjeHYXZrVf9feS
h+xS3d9HMSyAa95rPimcsEdkEPXEBx93kUjr6+epEOHPrm9Fzktcv2fORRFO3zR8OC+lzdQA4fkX
KN5ddR28pmsPYOKKURinS9H78Ng/CePMhdcqImwlaRAnLwsXRmoB70r4VKBjVVYj/VCZUQjVwAPx
xWdiREoN5q3NFxluWzpoz7oLXkdjf0Mv6p4IVuCTbUTXmorQ0XNDMl9/uNNVLh5aQxW4qst4sB9m
zSUCLt1nj7bPSRiMjX6ikYAaGWm09CyGXjEElVNb5zHxG7TdOmbh8hd1xqFS1jV+6jBfxR3TT0Gf
gKkSsilY6xECCM/xWwEuKv8eWmlHWsSkZXjIlGaUsFm5HBtsDeIDsf/KEcoCsHmWISCtx0tMcz8H
f3Y9wPC6OkkZkam4cr/v8jmOVvJ/C3uc7WTVmFmO0A1NA7XFjk+tk47IEiPOhWUaH1v+XDjzbc8Y
XHM4YA38fdKz1j2GiqGOo59IQ+wEEWIHvcZ4HRWHT4KsxtOaHvj4xOatWNGCqfAN1kKqHcLQDElm
5/KbuLknFsmBTGJmbCHT5ePwaKo//9kU4UOn9h3QP2OHKZPOb8MRmFvjcGh35TReybFiF4KjRi0A
ioBm9s/YHQaoCd67LA+TUYBNco02s1ZedFV23mUZQ/BYDKa1g/Vum+Tj6gQze7bOD9MU7hc9m3cI
DWgk0DeeY4aLeq5YbjePH4Jsko2O7nCx1iC5erVFv8Gn5Coq4pOsyGh0q5rtJgk2bYW+swwnOqIj
p7zuj3fDbxo+uURZL2+J6H36fa7B+LvzQS0y6Xk02/HuYfgXoA5wJchZyvuHVcJoo8BkdOod+yd9
Ngjdy5LfgMEE1tRHNL63o1gb6OoD61ZoirNeDaks3mz2YWHRBu/HVDgtjME3lzGinyh0gDrTcWfM
MiUznzMIZHvcW2WfZodnwAvCRnHSjJqj6ek8b2Uv/qxX9A0D7zkZiu/AfXgJOvkbRHh8/EQ8Km1s
+xjO4egfjNZMAuRJXLPZg+2yhhmzAb8tOAPpALba1DLKOta/740V6DCCYbmc4aXmhNMGWiVojJ2f
md9uIyD2nNAduGMpZImhgaFlPbR5cL9UcTRkLmcOeBOpiwRXMS1nUvf3MNGdZOmC11PLi06n7U/q
vBcWGixGVTiQHEe1uyBupqaQqE38x70s66mZtJ/+KKkcKXZVDLlNJaYu9GUgF3bbmIXLNFy+sWOO
wHibuTpv8gEvze/MUAisqy5I4+wDHyPX401+1qL8lSntGXtxw2QBNkp5Zfdt+IodowMaX0ApCIBt
02K8Ie2l+8Lru0qrepbdzhqJJDf6MchQ1srK+0KBHpfe5vu4u1t/vkgGBEmpRWJ1wqDdm9sq09Zk
r+tgu6HsrANrk7n7TGo/NYzQUI20koi4njHek73sLTtbUY25Qup2fwSnp/IdiGtuQdiucElhOJea
tsnD0YqbO9LLNIndvScRbTyz1G4W9T291ndqpCleV2nwuxKwCOrvBXJ+y5107u/gr1O8DTk3fqns
4N2xPN4R6sHsiV2s/vsmNsk7pViEhqSRjmhQd8qjZKYOYdvljTfNuKpbzOuuoA5nWTDOrwzMPreE
qkw4ZzwBQTJr8QTCtZ1rwx2eFUkjSDIe9ba0blJIoqXa5EUV07IwrZThyX+y59FHIREkHWZSYzcD
tmVLYTX9sz5MAkTVTupPOnig6RJN3v3duFbZBGANfmMHtjntSJUQkH/q0T84jqp9mQpV6DQPw8lE
MjM1HOi+shQXJ4a6kQbq4dG0GSumryjTi6zFaw8PaIiYI0PyfyeLliHSajWiVqw15iLjCJtdYlH6
pD13VMeST2H0Q5o3n1OTjTdtOfZUc/lG+1rwWhGzfWrcUrHXhGinieJS94v9UQyyY2p2TOHQO7tl
YTa7r9wDiKdCweG6t3vdyf8tvbaSPx19oNP3hriYXMfwFyjGiJ6Cy/0Afkm54QAAwCBuxT6vQ4Yt
aWqi25Ek0EvTTX/oBW7Lr88gY3j6IRdSbSNHVxW0Ensan3xXSSPtUymvuyXiIuQ52kHsOTeK7NUT
uf30I5gHBPGPMq5/QIXqYS2Tf8HydHsT1P4v3C8FmdZn45q/TVU61KG5SZxfUPcg+bo4iaA9hzmg
a6vxGLwl5bxP/nPp48wIcwXeY3/AEpGjtqmaEBnhJGBXOToulND8K0JiRbm1amgG8J4qXCHL/Tta
OiNY8lwZOqb/8Wx5ZBKEUVvAonI2SGCmw2IWqF2yE41BA0KRCh0jsRc+lFCJLj9i3crO+fRYHyE9
Q6niVMgHsSfBPCGRcjSKVo4wU6GG9Dz+0wxzk7q9akUZFlFNewb4BlslnFRSVy4MI+heThkehjZu
lxg4J83yrGy2t/PemYgNfLcc+DBAPtmRISQEMv2MpH3zG1B1+ok2/nJBFaYlI0ZQO+F+aw7X/l42
0bYDOtfmu2WS3NeD/Fd4QQzz5yD9wRMnKJ8O9hWRdqBLfqU5UxRsDorchxm67CrUv1uzfNSYKHeP
2qavphEpD2rnAlUgBrZNEx3MYEQ/gEihLKCyQRqz5FvhfekbfmLTyTKfmLfxMIzTaRNxse1r1rv+
FmwRxSoELEsa+ILZxFi3uZTMhBxOJRJDwBziyzxOm7hPJ4dOTkOZgqzRyqbgw9Lrj/iy5WaIc+pb
e9YCaHxZOWoUp2N/rlskfHd0BJ9jPcpoiCziXrZqPBo//hqTICBDPCW6ME3yVSUg8C5cgNkbT058
usDfyscOaswkchBlOWfxIZcmTtfwc1e/QLYpp9V+/cqx8m1M1L/DhSKmHeKgsDXSaVGruPrvas30
GHgaahUp9cA6gsTu8LKoj/hFxC+VyB2BFG1ZRvQmqFx2irM1ec0rSiBEafCvpqgXH50GMLvyeL0B
xDLYvNm6B56abKy8ZaYSnxjAwZUNyCX7Aq4+CQ/hU+QeMfgBrVD4nG5mCxdH6B1ByHFsKND7EoS8
2FfRAn3l/PBFZbzkWpoNEPDNhnnnNwDTZ+zJHDS/1h5BnsmLpDb+Wziaam/8xuidhCObs2XrjtpE
PNKNMOqBj35t+Fv+fBSGNCPB1sbO63rz3Aj1XTFx6Kq9v555SZhAZyZ3qiKL6JBmPNtzcksTsMDR
a/yGHDZYIhYxB6J1tEt8xrBGDbVUyjyukU2TNfzFguSZ2Bal9rXCBCo0G2Nf74HeT7jl0q9LF3Go
5LrBygVhFAk15Gjqp0IHm18b3xOCx/jtONBil5pFMVkxXa4vD+N0GSOYVAV6s5gPmU85iu/UmdHH
mquRKsZLzNTIKiDWDB38WKi4c8bs7+mZDXFpuAthTmNw2D+lp1fvohyCOYIjt7UEsrczvKIBVsVn
I0jeBfE2sOBO/q1j3VXl654Y2exATDsZkVTkaGAgf11ywRCYF7y0juSqDzk+mDQFBTG7kn5Bjuva
Y8G/pteZtd0Y+4ZROAdE6frZsh58KNteQjwnxa8g9bAtL6PmVDFEtmVkppbRePCReDJqYjzm/fdg
vsR5Tf0YngTHAhIZZ3lx0Gay+YnCOpSANzHIitumUqJ9mMMg++HhKXIO/nspHWLuWiJnoSWR1i5e
dbY+TfXNUpvf3N7dD5F3GlcZw8j81G1lEsrpil4z6jrtEY++P4sq+yGKHKEbX84Y2JBtwMKDM9/O
LiyxagEyEjMtnFc/5D2eXBxWERyIlrBXe5+wsP2k7J0y+VcOcIufFwyXZ3iODoiAqJ5uM08FkIDI
k/70+JTLmAQTdlHG11K8gfvkLUvu60dKBZqu6dNgfbGX5rjCytrjHyVTtjwxKVN9CALUafe6tGce
MoQABLM4DxfBn1+tsSRfnpRHWjXsqTc0T0Y9uUHIHJSdkflDAEdwPRCpviTfZa9436d3dVqOSmyF
FCWfpejlngSlIa2tiRjqNbCs4DD/CLtzoFjKUrWrPJUCxeMdUCgdeEu12ImT7W2OrwIrpHZnZGaz
mpf5QMuV6HgGn06raoL96MUdUmB8EuGW9JP/bbxwPvejqYGFbc4BQLp/GWvmPFaHtSKuORPmhRU/
pDRTtlYQSipxTii96HdGs36nY8qVIaeB8pTOtrWKJIgem74MIFy+ccY2mpxGa+6/8/MI67t9VfPz
13xc9dvaWA4VxEXBpZuz905stzozHHTFP2YDmnL3nmW+fV8pg39QgIC4bepuHlbVoR01leTc6Pmg
8bUP+sO5MOXejt2+K1EkwZcK5wYAnxhwUiRK/TZsG2r+OOZfi6S4XTdNEanxMNXF6GmRGOylVrMO
1CrnpXw6B68esSJM7ZSrBSJdi/lOabnEThUpnJwmOaQoFyhrPB8iyYu09g4q1EE4xY8k+12D9gqB
SUOHDV3OV2ogC5eVRCB60UwCUC1MzAKcTo67QFu99Lhr+f/8pziGNUpvJc5L7PlPkgKsNt3+PtJL
DLWqNTpc0kmMR9aBpLEcR7DPPr2rqo6YJTs9Y+cYJrLkapjCuDdGFaOuMNf9s5q8W+TYlYr5jF8J
1TYlQQ5MUPqpxVGYBLdWPWtsITrYoyRJprFQDltB8i1LnIFscq1xaGcAztRLtwLjrd4hWB5oDMEk
/T1f+iLi3Tad2tX4KVzb9aJ8xzKnQdHQNeFM5w/JkKP6ZmDYqh56myczlHMqRgK5puJq7C20odmC
P/EcGuySrwpCLU7ExN+LU5fd/dlouwvZvKMNcd3H2oXJeyEY6i4Ws9hAoE79ylkIWtAKPUyQIwcY
vPs3JT4djC/IguLSanH79ZQU6olPbpZItT5/Q80yBAEauxBB60pwCOW2hq0YXMrtEIiOAOaRJ97v
LZnBE/oqbiChSOw5vTVw53BPDirGicCjOpL9JZIy/cjdJ1CcqLRXxIg6utx01ezUtvABoUP/v5ML
8sol8kTf0i8VrDKZpVWTxQ9HzB8wnECM88C0l63C9iyadaETZMEsxXsgSJxlZ2fQE9DK4s6J3xD2
k3HeMNXta9GZmd+ZvyDmqXK9IqzwHShmfnzE9fwDrbO0WW4HXxmxzyoFJZ4Atyrt5gh6T4CR0Wjv
gYAfm76FOizHLhJIvDHF8wOmTIhMruIQIVCgtic1QMLfZEpnY5eyBIJefORxhpcc46w2Rf717Kc5
WiRkdL2xdxePQSymWDQdLbrGx3kXpS2Hb9/3j2RjdBQ0Kqn2bdjkHXPU+2CArmipyc4uLI4on6yL
haT5VFvXK+qs6I3b6vdiJWoyezFv8vOSHsyWcamN+c3GFKrl979YRFR9sC4snsdqrSyE9G4bDT+k
XQrk+Tr6qui1wPApnw8YDvlp3TtT9VBEoTPWoLcXcSGhQt78qllnzquctioBiR4kn3kI4qY2fQ6A
N+OyIozafkESBVCoDbjuLBXw2S1wdz4QxoRleiBpDWzgFmWVFql+8jNXsDxd4FrzFor55AaHae1y
AHB8sEY3eHyvFHbhtDHFDWGBuNAx35Vn9Un7WT3HXCOhTg6j9nyDU4lf6UjbkV+p11FXCCvRDz49
BC8s9uTVA7dAOcTgUXJsewu/G3Ya76CyqXY6gTr1dkGzBSgqzK+1+7kzMsTfIz3/gQt49KcM1+eO
BdUtXAmiRIx8YAabof72+oabTWm8uLjay6mGKU3rZ4I3ChmxoN5gFVFPgRFN2kQcLI/KKUBB7ljD
KdndrT8tfBSSw3DUHQabvEWwBAZMX63IR/W1cQ3+9OZ9cBdZx1ydWlMssKy8T4Tip6PEqn64G4Tc
Ll/kLR/e+MWCJEDxE0Atj4o92JF/Ff/breUF7+g1KmTLYGmW6/Wew/CoyLH8j0E3naAdr7BeE9Ie
l/jJwU0uq/UUaMDtySpYA4c79FrW4lur7b26hEHVwYMccHPBMONHEAHCgDmK8ab7KPzC+H9pUqUB
STAaoBrYi81M9PCJNdOCLZEe5dXhn2gBZIhrPnNo1VwAEjJ8x8SP+bKawsramOZCOv2+34t3Aq1p
tRMp6OEGnQoSZ2mjFb2PdO3uqpgrq3pAMDT5Zuo3S6h4+YEgMrd0rXTQkJONzl0Od7qXhU41BirQ
FuMomj+N/ds906FoZ4YyQ7JArCDph3JTXZQivbKI44p+t5EXTHq4TvZFqadj34/XgcERIiCOsD/3
Wqy+0ZEHiqsnJJMt40X46DAss6DXJJrNTfYNtck15jpP+r5Q2RAh9LVlRHlvyzPX0Cd/O24k/14u
mBTzOv77jC/paK0MdWMEaTjN0rktsPuvBnmKxxiYtZVJtp0r9lTJVfMFJdzPMnCOHsgDgpLAa+vk
7iqYRPMqr/iql69xLvLgwchWJyyKearAOXKw9zsyi68QhgVpQ/tTttCpIhjGOteQ1ZZizo4Te35I
W8c3WTXM/dppL0KZ9bElteSgEscofYsrrbYy0pZpYdkpvOzBQhYGhkVooI/7BeHQEX5uFXlZWf+2
QsU+Z5U9heHhBXn2L+r/A6hg7wekFcB9p9adA+KPNXv0/A8CeAu1fkrMcV2qsVdJ0/aR+7+3DK8+
8I7iNIF94FvAm8SLyiICigQXjqAS2ZMgNxzFhXRQBRuWUdtg1ADRJqWYhfbeaiB2SpkEMpXe4m+V
z0PofhwBFrDNFM0wWsvSploz4V8WVFBe8b3MO4kjFtR+Q6rxK1D48Hgw+fH9st+X/HEqhkaJJvZ/
UFfPJdGD/6APymzcHwJ23xssZI1B0JM9+mGtZSjQQWEQCtXwiJYDStQDS3P89W6IcG8B/8kcgLNM
mSq72NoqOLZR7ly25PL1f28I+a4ufLisHe7EPY+d45ETOtEiTfHFWbESWFAVFDdShOSDtmb+fnQc
m+2qyiTYmDA8CXEpeS86tFee/BHUICxntX8mk6QA3TnBMEYN7dE1dun62fAZmKL3ARu7HYGoM4VU
14j+8dnIrxGbQkCvSJNpUmYjNvr5vEw9amozvERPfYEo0z1O4fpeYOsJ8TH1v39PuTSOKjbH+xJn
9t3Dytq7jA/oeOIM53hktofZDvpvEa9/83ie1kA/jEHP9fdm1YNxksFizkjlAnOuyn2tRNav86Av
bxo0sVR6f+HQFZI98heeYT/CdezHrsZbgzDZz4u6czL33Fe4Nn4Eeby6y6kBpLv+h3EXy8LxHrN4
daz2K2GD9UCnkwsbxJkZUs/rrmJmW4tzojAZJVpL8cAa7CW/7xtzt0+BfBwXt1dxrp/VnyCoF4+c
jH6cCA0D2PAMjlqdeLgujAM2xR+6YsDeao/hYgJ2lO/oVIStlt2zrRmxxs++/kNracvf7TaVPbvU
wIkqCO7p92N/xOk0hU7KAaUVB+Tn3h7GIYmcEmsUnb+j29CAyM8UMw6E/KcPUDVO8DphyD8MLibh
esA2t8cwAvW/Zy98TeZFOPXM+KnF9ToNX4YquSoZgtTJyT3Kgs2d/2rNU7/Gq24mBUKsf8k0uEx8
pdHjgOCpaf0UrYHxNHeOB7URxTfPQJafLAfXh7Cu9dsF0h6yCpUB/iTVE/4q0VLqkGTP//hXikd6
lQG95InckoLr9JfkEyaVuKEcufmTNokyn33BBhrYju2tVYd+MvVmOMBql47J1IhoC0HJ/2y+tguF
4sViMLtVN72kO/LhCojeHIimv2MNlQFMB1fAVK6myj4BRskYgvzdlIhm7W7xXQKGy2aTnA9GwmOC
ScPROCHnABqgSzeiTAGHlI9mJjW65eF074PvOa+dKLEX682tY/S1za1akX/tMsdttYPaybcgZsHD
143aCAaFvX1z86tqcHI/kLM8VWq5vC9Afpgk+LVcIRjuO2rYroD1khOAixFxPn0xnIVyeVA1Ts4q
1wFubHVD5FPVVm4kSZUeHSC2XwVynk+40L24km2gXR2+SE8jjl9wSV0XOehlKsKk2umkNB0ZZwNC
7tIPid9YHmj0B29hLFd6ci2K2W+AJQdtiHPhzD/dcWZHiPDzaMNPtPV3er5Pr2BqHY0M+WnLrYWa
ScWi7Qbg2RW6aPke8JY8fBjvrXP2d4g5WyNgUBEx2YsfmxsbR4PbXfthEtUpi733oZXpstqFYElH
uzBcgh7KycJJY/Ac48DTTFxJss0K3dJ1Akfd8Kpkq5twxkIwnMp4GD97tk3AYTgUYw+S5spKkh5c
uuFuxk/Dv9bV7bTWdeLpvifasedtvQrjFQIQfKFzEFa5rWHOQizqlwgbs5sQ03tHId8ZKT8b3fnm
uVqaD5m68I4d7gbG5zTytC9P3Md4aX8Tm9JEDXM8hWq6/i/BL7aJ37otoD/aF6mcZxiempij2FFH
rDodRfwnbk7pFOhWGBU0PgDFaeR3cyruhr6oIxoHSz4upE1G52oHMS9E11BOenCYWNDRMyO6K2WU
m34CY3Ykh2+dT+lV7Ef1jjFSOMgULJ2dcK9csyhFH+QUakwULsCV+3J1MxyQplId2rNouC3Dndxc
Mj8ciU8wUEp2Nw6n9b2APpN2TPN7HVbFJvycVFWf4doM66Jxkl7mz5LkRGPh/bTLcHOClZAHvGuj
WSy1P1RVzl6mhleE6q1Q7A4hcZu/56mTwPawWLAeecb1DwEzRwR31t96B8OEgrpJWdObAgcQS6Gi
cFTv6JRGP59BRlquwbHuPNWBNxMd0us0o6eRFrGQjfUi9bcop36F8jmHHOthaJd9fH7M/99FQWo3
7+YlQHMyEY/M9E02UeltI1mamu+ZEqwk7MVCxuF0W1WJ8Kh0bHH/NsuhGFMFzGwQ4jWXs/3t9jWT
MGx1muMne/RArtN3DDqFthxFHsyQbyQ3z22skwgeit+gI4Ya8H4W4KH5eRVRy4IErdgKGE8PFcbP
+TMtNAsXpWwoGHnM09dgrP1xEdNX81WlYY7ky8nSWrcdQCBpG9nQkdzGxoqhQLKwx7pYoppKzUfV
vFOrE7+AwXmlJM+r7MejOeyexrrLzrZqnzunNJEWZme4yBinBu3m8CX44GeXwMNb8cdH5RPRZZcK
29qD3N8A4KmLcnA6aOlrRCh6zp15iQDNk28LN/A7XMgSaXZSzpGpO5ZBC4+YXCFhFy2eMGlGtPMg
39E88xx3yqy9gnN8ExDTWwL4ASEsKrNCOzmNugkNR9MbzuWee1bTswh1pj1w0P/yEFPjazkrGxL8
T7RJy6htk221qHA7KFzx1Bc9SpM3yEe8k1X9un+EHBlDY2+15WHc9h1vwGXX2baArqCN5TW+OdPg
ezeAfflFWrU6l456OM8rjCJ04FlElljmZHeiufNhJulFvbE7XJZUezGFNPzTB1dtStohBDGAKn5Y
K4jAN1qwaWCB2C909vBZ6/V5RIJhnmx93Mm2xJsDt4Xg5+iLkmU1Kn2WuEktpo17hiUZ2dyWHj3S
L1owMPaNublGxLv8thjMs/6TJA5Inx3YcIaRRw52sG3ts+AlGWKe92sQw2QCHFjJrNBGStObEIv9
ZeXfgU5OthUaN7Q2Tn8k7Y/WaPpTYh9qWGNTfTv65S4IxqvbMvz/BhdoRhlIyhNVQCr6jy6HglCO
Eop6xSACvo0dMiO5Z4HkueW7H/Fi8Nk4+AS8WejdzVPh77uHAVG+Nxzj8/zf8njboWmAd4j/SsFu
CdE4jhooBU7sGwS5RckgwAzTwGAv2x6N/yFYOHZBT+zwk5e5VPiWr83XLsU/n533gy4dzpRDfdCW
11eL0QmPXmXegveBK8HHXjYVThh22XmqtBqoJgvQZBM9BJRPPcTxBm3me2RM8B56VAdnwUshg5L3
Oc6hQHwNOU6+0Jjl8SfTynC015i0WXKA1OavaRXlQSWx+IHMe97Txx7HAoQ1X/Oz4s3LVJOIsW0o
gghx5NlNuZ7Dqg2WdcgNMRXEXZGuUnKZ9WCY4iwP93Yja0Q8yn4DhW6rrAg7vyBI7W+d3n4Hprz0
TNycxxIOh8WEYK/fuYJK2qcKMwI11d90vV6wLeq/R3D6IKETlTsa7P1QeRe2dFP1A10KQWmeiDje
JKySR4hMw+7wJhC0JLlPT9dhWq5zi7sth7h7AvL9VR6DG13xcmbtZPlIZVER6ZdFLi9WUieM+Lfg
cCJunpbE13K8jzX72qPLocPhVHNN6ucC0hOP3jcUXkgQ8x4C7gnSyfR5WyuNyYqz90ATO3kLv1J5
KNb+hkirh2viFjyJnxVCa58t24mOcahq1chUluGKlUJIQm+BwIaskH0KtdNUBvgNqiyZ8Lwv0Nvb
zzK7oRtHzeX2JnMSFRBxl9MD1mWxHGEEkPYEBNqlw+3K8BEcNPaXx2QabyctY+opAN6oTl3JjCkV
yIA3XmSSqY895xntiqx+Qp407lNwsY7rKfD867XPMXn8h8MdQIWLdUT9nJ5scEfV7vcdYlOpmE0P
YdxTUMmF+eTJZbafNu31SBn+v2jZEr1AmTsKNXtnL461FJzejE9xtWbeMRBRUuauzq5cibHABbzW
aCtN6xsfuXdpdgqus9UIswXme/ZWW3TqX/Wf8fs4GVh/YQnW02MgGnWs59THmTDMOAYTjn4DhPmI
holAFtYY9IBEnd/h+3RuaiVQKw2DBeI8QNIrEgIxIsS7Qg6TMAwqgeu8ONYokjwXysbGzlqUNl9O
vg5TDBNhOrLEtBCbNw0sJWmYASvM05aLEntW1URFm9gEjehmEWEHK5DVIALou8uAMu1yJBXI8Dao
9FoErqyd+GeFslJ9M64ucEv/2gO7UyC20yB5hep3g8287C76UBmkion/3YFAzIgDBWxfNW63uJwi
g7rN35m1DCwguiiR2hG6tgrTWZOH+Nhwz6F4o29TJB7PboxLBaxZ3pk75ahq6s5qK/eUH98Jq8zv
XYeuulpzIZUXDqGC2XVL6tB2dFgx0CfKoYmxLt6GVmfPJ1Uw8dIQDWuOMtB2lrk9+346a9zjVt5g
EFicxR4xsR9CPMK0i2qo/BowgpeoHlOQO/o7ksEkrsAftYq8/b/lT6TDPyAjJdyhObQ2yeBCvexo
umw9eoI2/4qlUE993jbquwUwZJyczPnS5XEMRcnm7Qtyo84e+9yogna9yeGA8UQ8fR4SMEUSCHVH
dEM0CI8Pw5QXIIdy2y9jkty0Jtz5gUZGzlXd7DaAb0ayqV1aKi1G8X5s6uDp4NmGzV4HxRhL79e5
Gm01sEjMqzpDL1tOFVk6c6jzFGG7jNsosglPy7sDwf2q5AKoO/0nVCcpvlLPXI17LriAzTXfIrCV
B4tVnphs6xyfKNWiFgVLjnF52IbH3U+NGI448KloF2A4s3g3vcT7S/ncsXqkV4Cdmp6oncmiXo5v
DbJhpE9+IkL71Q1+oCEZExObV7hMKUAsu/d5r56432ZNtNKohXqZ10QK0WsbmAmUka8FcWn79YOE
icWq58h4pgTB7lFYaaXDEIqlnnaHfwkxJiv+ASDI191LNk1oKf6SjwaUPUBYHuAvcyrsfKqupbLI
zVQrankQXLOdrj7fOOZLVBHgZfXfRK2/D/qh8wbPQgUe4IVB8iY5HwKn9vpXDMMh32oA37PnC1xH
fzvyHj9dUQ1q3rrZtujaCkiZXUw9QHvKfc5Pgyqz0Ot8m4XKC9spYKj+4iromO/Uzsfd0H+DCbeB
4uUOGx0Y+VI7u2WiABUsFd3by9OaypIppaHufROQa7BsinR9o9f+4OVZMq6JPj8TNCRqXhMDkzoq
hVLV8Zy+ylfsQgLNG2n9Uy55uKOSOaQtXoBOnGEr7XtNu+719OSBhQvmCEQnEWKq+azH/Ga0aSr0
031ChkVAsdwBgAYKfLr4h/qlodIJ8bJAs9SCbyO8kW354OCZl6NBP47mDjhn4LY08BIl79v0OS9s
+v49jTnRV8q40m6Zyl0tII8zXOr9CA+1SufByzgAi/KGtM/6ub4ZbQXBj/0GWs0hzQFq31cr5jjo
vX1J/E9RRj0cQJT5ktse9KkzCqZ05GYD7ov6gDA8doN+/+tapqLFRlirdsG3GpGXnUKwQNRnAl1X
GCd16Jr5k1AP44FcA5kz0FwQ2ubEY9uA8It/lVep7/kDMknhAlrFHtS3DBrHHxAH07tmprAQgXCC
UGctd8AcbGui0OeKR2FGdLqs8eo5KXn15xoPgjSyuDdwSj+p4exdjM4TsR3kdgAP5T8VvhHTNRzL
m1M4DY/gR2k1LC01VmTqXpaIK/TBI79/ThGhwd56glOy16hfMGRG80qvI13hBvyhSTz+B/G/pECO
CR6fu50AGmQFtBIaHyKe6rnY5dpYLLdecgQuErvlyMro4nUyBpF4G52TsL8fmxF1XYJua1K8Wqxh
AVf0vZ5iCvTN6Hp7uirMmmK+Z9EpeST5MmHXjoo//wsAZWg13jf6mKYCkgy1FeH5UxUtgHaEm/0e
KA3I8dpu7HCleLwotmnrLADhXTyh+2a509m89eIN5WFNtJbfJS0sisicb65xgg3E1l6AXFykSKBH
XTIqkhTbv7KMQlhzX1i2nFRsiDlYoQGFsRJiiQ3aYP1cBDOIN9ICATdLvZwERya2NmU25t9kmY6s
dBBHLLHtGkdZ3s4fBkOJgL6ZCFeIbs7LL0hkvAAqdPD8hI306gVNy5t/DrVGcv+GRcWn9K4AfOl/
Y9Eb2qGJKWwNfxMR+hAngT6rydHAgwJai9ve9J8UBxbNG5W7ad2HnSJtIVMhRtRnSw6+uDEq2PS5
5LFyEFIhK3QwSAc08otZ6qiFcTm2rh7f7ZJ61SK1nRIlAhHicWwv+z1jj0zC6jST4WwMGkLywy9J
KuCv8pTTbjBSUMHdpQH0+erLd4vd3/Vk7ehOJMf/4kp5p3ABqYQuUFfCQeYWFd3RmwNHUu6FIsLZ
oVH8uNB2sYH+Plv52rE1R3WosyvPO614hnEh3tcY1MGuZ3kxMFVZ3L+mWcS27ULLz37QwSXc+uu7
P5h5kJMoWewcA4z7uWwkzAqGwS3WfsAaW+wapE0uUlVyE1yLAUdgMGUC/kVs+kGAYsVpit0Tgam8
UPX/9+v/tvlLQDa3m2zeOoOe6KgNkc32dROuOafLZDyaq3g2JZOvWa295D+r5EiOFvK1NuXg9haZ
F/zXMwl9bnL1c/VH5D7Rpu1Q1ekxMg47vcDJJOXQNIx2j2dGCdZboQbecR4qiZiSFT/p66Lm83ev
2xXF6toxRgPcH4mLADgNZqeCIrqLXHilPTTpOai7p0tPVcX4gRk6F4zrOjWq8i0GMTO5MPTTfSnl
Xa6lOlj5USq4YPkX2++r8EydpdqHJeJwv7tskttSWbFNSlKjl9RNYEteXTYJX0cvQaf0NL8WgEvu
CxS6Yg4uiSFqYCHIrgXJJDEsp95JNmvDCHT0JEHEdEfn7o/jq77sotv3AtWoZ53ePSD9cWDsl8il
i3f2vn+L9zCnXiDeXDmhyW838w18ugh+sVcpktBLIm5f7E9sonJkS73S0403QHqgdVaINWVpy5qA
s+E96ZhCoaxiAK5D3XHpMIFnVsIkPXHe9FT05O9AC1VukgfznVRvEzgZ4nxs+/rPIep+Bms15eCj
3NW5tlY9NDqRo2Jzp0/S9CimcF/W0qr4oM/BlSEl3spUTRcLC/pyNF3PRPLRKwTUSmvfCSf5qhp5
aYhshjMjfHl+vtHqOEz8IFi7TdfWCYceslzTXysge0+uxhmiT/z0yVMl3X6PjO3kNYOayw46+Pup
zcUHjL3ilTAU2UvFkaDBz7P1unAe9zjCoXu6d3/w5b/VDgiH+7/EqqFP3oV4z+JHylLLtY8sEntH
FaTFHTKhs8AFa9yFcqXfVgTIoFZtApkQBmyrhM3fII09QNE26z+ZqG8QvaXnH6wK9b1OvaVtCa8U
5k2BONhYtyFcgsQ2e1qd9K1y112JKgbDu7BvITsbFNDsmUppU3uGl4YJVgoGBa10j64vfurxN1h+
aSOkSQlC2/5J2xJYTWnZCoQdsNpoCYwMkIUqvgVkDcj70CH1MLhysfLmVnlxerYJ1HN4BIRldv7b
ilZTqx1DcVDaB8e8bNNwms4ZvSTTH+NMdN8ke3NN2zrjHheqHXxU7SXG7rQlw+JiPszdxaMwu+jf
HXz5xnlVdVIRHTSC7VPsg7V+cxh5fWjJxqrGdUcuqyeYDltskqCWneoBoIxJfrO2WzCE+EkKmzs5
N7HKnCN27kwxITzwLmKM95xwz9+o5F6PlOPfPsp6mzekuonnkfZfKwD38dnTOajbHCMWJU0g65bl
R9m9dJcgJime4ZfTyHzpSlsNVU33sGzZAr7fAxhoNgH2LK+uTnmVwo3xunLapd3tS12nHduYZ1ix
8OsxUbQNxYiBy3NrVt4TZMia/GhZey6MyA7fbbjmPOAH0ODYOTvc+62SDagX6h55JM7k8YqSeTbR
tP1HvczZIg0kmoPLddRJWNOeajIRXSI/xJW1b9iFTv3fuwbThgUGxLu5zUXCGeLCnvKKvOtzAagh
pvnNy5wGPd19iaDv0+//rlvug1Yp+uctj09YlJ7hmyTgEKLNoXXkBDHILqpEsCUp5f+e2kao4h/4
ygy5T05KRgMjSGcnD8U5l7cJhu6JqtpAMljvxPcheSE1ogYiYpbTcMq6CHTr1H2+q4HIpmQ1eUTr
w25JwcC+GrqJy0JIkdZm4XXAxQzcAk5DIBXNYntzVbbcwUwDkd2WFW90robYvKN7tKxF7umD66RM
qdYH8rtR/auOR7mVRut2+oLFiZle8Di/fHtAuGhNDqWAsxf4Z3yPNLv5U+h4i4Vkn2dszFzGwset
Krdr4QyXFZA8efE3zjtwG9MmkCG7V4IzeZMtFZBjdWd/+jCibcjyNrTrijZrK9lauw7jPecQdMGS
gtC76nqParFENB+MZ+aMnZiouOviI2LJUCclzmgJmRjddHLRVnFK4Z7JR3ez4MuS5W/urlu73LuH
gXnVvDXTnp5jNGnLUOX2M4yO5hefjbDy3J1Tiurv9LIEvQF3g9zxVLxte/5ZvuMH96A7XElRTIsN
Vy9oGyaWBFfHgKx3EGNLQEI7f5AvQR1T8jMrlZEBWxyO2swRKUZomaJ7i1jdoXXjRvDMPy6V/1BU
Zyj3zDEkbJE5We9OHR8JVo3S73rqLpCAkvFx/I0X0XxYi2kmlkS96A8kMJDLVjtlp1THG3+7mXC2
z8HoSHiCw6U5AXzoRt362WfMoz7ESIdMWv/0XQwo6r1U0FyV+7FzaOpoRdFc6HJvkXl6V9Azjk9k
bPrgV3Qy9lmXieqUGxmyRASx2mdzvsUIhZ416efND9w6jevBai57QP471CG71tFanrMWmIPx3vm0
glwalBSd2qflSWuDu7CoKOtSTdW4HPpV3L3x77IAP3jKzoJcRh7BlrPAIDvtG+zIUzjvN6cuFRmz
6sGTObSkAF2tzZmwrH/ZsXiopyVCAu3YMFKFyy07R2ObyQvtIwyTM66QDjE08CqvOYlAnkLy2cNM
ZvST8e+lSSedsKrk4c0r1WyGbV88wuc/pxvt5HwsysIBWUJNABwQrqiRN3iTXotPix7ZzvrNUofu
8mbUwJNkwlTQXepuS2esuNkudbwOkNgQL+ZCUooCBf6pPjKD7WfY9ZStiiMePIWk3rh8uZzYY/ka
NrXFWpvZRj3HkMuYfZ7PWEmYE44H6ZoBAJKTS10QC9zWZKzxufizD1+EW4Eeir1xIqIDOzDCCZEY
9d1OYPmnV6h9obU0W+SVhe1d0+MJvxTDYluGRo1DUW6v6TDg1cIPtIDGxec/foj0l2I4SO4Cp5q0
FG5lxOiXMy/W4u7h4Aw2gz1sSafRxC1zs2cEsizBqSnjXhzXhbEntwXJ8gPZoWuaMWgv+Kw/VGQq
LRi78ZSIi7a0nmrp3elqJ1fGY8IzhWRNQ+Ser1i0nXZMRMgVpQBPIQaOEeaC6OT8gEePCPWqDwlx
crmtICA4Ejp3H5w8XYPwomn38IBSzRx9p6Xm6yiuYOhx8pVMmbTwvicFiR/GaWzDHec/wCj5wc4m
c5ygMf3DN8pWB68TK4yF3paCfVuFYkNSfA8dr8uytzuH75izIM49Afw5aJYNltLKLxpre+BWaPJ+
6cRvHAgwkx5JHqdg78dioTbutQ2+ntMiUTok+Q1BUSihhzOqXJse5OVEugE/8oq3kQqBRkuUrs6Z
4B6Uokmt1geKkVIQKhsmBxpmaEact1lgwQD3c3BERVyGe/aaT0bTM9T24VQFVxApMAgpa+I9si29
MuQiGPTww7Lgcf4TMH7BOmkkDdqv07Q5Vi7CgWdoNCFUwuuAdwvPSJCwitAuOpLKXPqvUI6Dt2yY
xPD92F1jka9XmUHkC9WX61h9fmagfCFx8/3AHicT+6n3NfyOMm6WbFwoApd91ifRDSctqlvpzvnI
qE0ZJRLNjQ0fmrqLrnf+WAT8+QwmeVdMIt2r4LLaa3w7LpBVFtvxsCbGlE+nzx6/hB7chWLwP+V5
1dyYB8fA3hmnfypCMkPnemMQ89vV/hmMZaCs4HVoeiFkZB1kkEz5L4kIuyRkrQmOzhWDs3kxpEaN
KmX2jr/qDYs1V7E9RfPrAmpvj1Q/TLLt6KIChLfNgzQqlzqBtLXinNnLG4oKhjEjf3LlRrMmCEGE
od4qhmJsn63IQjNOlbI2TcNQ0HtVIOjIK3pfaaKAJGNR1M/wGQBhqPRnor3dTKklk+P1KZ4xRTR4
zXgEfr2QMk1tLVB8TI1k1LgUqUkHLxrxjKXhWioaP336uxQ0ZcfMizCSspVGOAAKrNDgHMnNdPsE
SS5zyZitNnPO+DTvx9ZCfaV20Q7rQf4yaDPYYschqJrVRRjLAbXKmpRKYsrCRn/Aa5hy+pz6ejow
RRYX/vFTJhKLyAosyg536cxPlEDrHKBtb89ysyg4iLM/UgujYAIIKnbVMAGx9sLHWrTrnZJM5plH
3HCKGWZMi8hjupRkGUiZKfacmBYXsthw2WcGCSnTDmYKDrkD4oLK11QYoiji9+gajeZ7z8iz1lxc
ntre7yJUZH8atrBoEEzKpFjBk9EnU0feUQzUpMBZECXqi2JiSfUqeKBYDLv8jY4t4pqzPLYKg479
cYA9ppXvqP6KnjHYIkCU5WKv560zrKc8DlgllKJWF0ZW/HFrX8nmK7wWVi5wFoPaSDfGtFgCJXnW
Kp9P9Rs0gmElmEdVnyHpQA500mm360TFGMRHPKj7aGW7zqZ/QZj6pPwccaCeZvX805LpKQoYdWjm
mStbKno9xpIQ9MrspNiQ1aIYLJqaPEDll9LRTn81HTQNHEgKp1mDKS6qWKBogQixpvjDggPy2A3m
SxpNINVvIwUsBinHoUPzlkb0sFjBBA9OadAqkTfd+9GBONNyPz4AWfuw9R9ztymarZViHbEzam7o
Q2F0ounxX4m3oTmgpPB8zwgAhk7U319zxKJ949rUJ9ShsiaYwH/U4wUjzAHCCOc6DTzTw4GjrnOl
MrZsCiNVJjsCVhBLUX4xTugsZBypYYX0jfru8eydCdmAMZTzQj+wtmajEH6uGX17i4FMjjS0zM25
C/vP3n1S0nd31L9KbsM4/H2WivVLvmi2i6uCgJLZpPwi98tBanGhdCjIE4xxXL9bNG7LmzrNKx90
Pd/tyyWZm7G6UIrUlIrlQZV/K8YmEo5PhNk9qUVLDmTiVmJgs2taarrjsrnaZ9Dr5/pPY6P0bSr7
QhzUmhV73jpoZLZh3xW/73h16jxwj15GbY9PdN51yu955M1+FFrqNZyk2lRDZb8Je+EKnYW87RGl
n+E4BaVex5KjLiJ+Oqg0SzDbhop2WZaDt0rKRpFf+rgiEEQ1DjPujYsbF5K6984XHQ7Ow1ZCcd9d
rvc2zUPTkj93oGs4AJtUTh09G0GKYCGQKbACAmLVON8SGXgg1WAy5FegkxP6KVGovTfbsSIonId4
lnvx6VeKRPU/ZzynhfY7R8Pon6vfUgnnDLT9ZXLXglFrX1grCiBjp5LaHzCfIYLj3ECMMY++q79E
50SVIfoVenV0vfuM8X3s3pbhQm1kHCtwwmRs+VBkMvo3dtNukhcyxzzZ/W/F76Sd+wvFthjy1dBi
o2JstTvwBabYwtx0MdJrCPUBgpp/s9dzTfchrJebjWIVv1ZL175pI4ZKS7yqO5tcMo0nqaOIgz7w
YxV4PDDY26cFMYd1QRgzsVJYeQl5zOnEmyLywgnZ7MygFt41X4/tqmHGGYX5gMVLx3asRDNz6TS5
hkMfDGCyb7xV65WzTGy4p0W/UFTAopPuhyi6si0SlIsqH9lDY3P28+lF1lUQe9JEqMsqoWeU9anT
HDlz/ugyRnBrnEcDeFj9IXZugK4QtBTjZQ3kRBqnqu5vJPmBgVf9xyILv80mhVuXWzW4aSJQGsG3
wDARRRUG0AXWypPoipxmlN/0hDIgQXvacBUzzuny/Bjs4Y4A27Bw3hQyp3R9MGMQcaCyxqAWZLXe
j/MAwoywUs+UfCjkO+4Rryxv7cMpOUDXUfKGFJWmy79fHlf7Rofu/YtBsbv346xrlf015w2Z7XIF
4u0zsxXqohWWd3lkiQuhpFvuUkNbasTEVE9ImztYuUJQQSynorsPMHQBWh4aiDo37VLcQZJPJXUo
EEdiR1qnwJCLUqaAvyM9KGgvZJtlyMHNoz7OmhNLKPpYuF5OrZbrc4hb8TWa+kwJmyAwwzgvJpiY
C4n9v+1aK2gn62X9aUUDeCUmUrPoyhV2WvJwmUpYO/SjWSKHlbAq1MLkQBTPEDsc+N3R41FHVhhi
pmmkPrHGZMvbYO3fzVXoAR0oiNE04GR2DXAZiEbl7R92HRnIUZoEafDOTNEBmnT9KFBmIk2ZiEKw
zQxzlZ20GTvt88tk/EwdbIdFMEB5EJjYfXvL+TZ5Es9LBFuD2PPWCQSn3Q/r5CThNzq1OLHGBWo3
y+uND+pz0KBGIOVSjXu4qMD++a4dpQYy/+uI1f/Z2yAAs0MXgrh0P5LPOzdkD9loyikZu/KqDt2p
co9l7qjagwEhNz/Gt9X1rBBYlyGIfic80Hz4vIMgkMl3TaEuaGz0eqfypVClH7W9UGElu5PZceX/
7my/MlPuZvG0xAS7Pn0Z8n1EBud3uTZPeqZO1pMr+3YhaeNpNyAQbLvOuFiyl9vrFBtD6DHN1DbP
1ueg72bpfOBEBb+bNQqapspwl01B8jvENfV/oong8s8sRsWXpaOXdWh/cQjjXy6SUOt43vGIjR7h
7G7uvOqMiLOF020Hfame+3QztdC37AUxZdEgFAW3RhCcIYUEY2lk9pgFiZJlaj6cLs6T9cVQrZNu
kwLEOY2KQVkFnOuyuMl9E4lPMcRS5uUDoGi3xlHtEdBTOka9iYlDExVbM9Or//mIMGlXbm9YoKlk
jPBBS+QZWV++cDFgrL9i0eSle12fi5aWl8ResC9Y/AiiM6z2GWUJPhQjWbrKnSSrZ0VlEvp/xVo0
KlRn5bddUC869qwl+XUbW0IysxyTlEZHnIYns0faNhLE+qmFxcH6l7RaPAX8+jRZVcauyEvcirc5
e0+qpZ86MFIW+6SoBzr1nSmcpAs8DigchzpSX8+VygOM80XOwnfkZNMVMQ+rWyqlD73POpM7YHt0
yJAAqb8xJSot4tN7TaFm9gyOVocPxP5buXr7kbNSWHBhqEztFe+5M6lpWqqVFNh/+R2mB9FtYnd3
GVK4yt9Sjj5H3qG5wmAezxiOa5HCyJCX7vg7uymYAUXQ3pdtakLqVE172VtWBs97h7dO4ZX9lySx
avz78WHSO2YelvicUzCFmJxaubYHB5xRo74XwumheHfKEWZd3JKGMit8CK2ykFcdjXhzK/h59knO
11xYNBNTuf9GsH0iypfLE+l+YNS0dioZ+LvgFwoq/2tp8SgEssVfrN238zYvSbSqcJlEbvygS98O
9X00x2Rn/k5q4/RernTpMmUy8xwjXV+zWVYMPASf7JgIQkZ54MD0R/HUl3OOHcxX+h/K10w8ZZ+s
747BJULtELzPDUX2qMGttg16XQXWacxbiv74p6V2hLyrz6ZAWcpuQaeMMaYdJam3hj2AqaR/zbU/
YQVdKL/2pyGf1Sc4krKdx8eQyK3p4Hpp30+mpEmZGEdswGQ9qBJneutF2N1CG8RPmyBqmyZrK+Xq
TlOUTvt3vsizYMwpOnjFMH93uvhYFyvi7yfLPh6hl37Yn2Ld7yhz5ee65+kR9LhXMfMfa3LMMSt+
1wckZ+eDlC7/QAV7agZZklXQBbvbvhunN6HBo3rjNnEAt4rOySyn318T2837Ous9zrDp+sujYVaL
BTUuO/kighYF+FlzYMBEwVysmUaQQIgyiLtuqXo7t4qZU7i3bb+utxUozLSqGZ1ADSnmpR+7zfzI
bQVr91T0+37m4ReYY12YZYFXeAizdM+2Y+1YZvjcrLPU53VRzKHcw6JVfQ3A24nA1/JdcQfR+B9k
NR2cfp069tRh6ptIGcKigHSuKUrlaItdLGCPTp2deucLfouhNDSeeIizLV2v6yBa4RuUJoW5GFjn
kPeldWu6RzTPvpK9LtEJ2/M8Fpk0EiOPGAoqzgod97NUx9vD9jD6bMC04p6i+OhLFMWy3IWEMdFC
Ju+njgseJjXTZiklrYhqqVFghh/X4vW6OEnXVFW13+AafeKs1gDN1U82dT9CdT+h/i/+ldGQ0XdK
J188kws86tJVM6IVfepnPiIlwsv7sWl7z74Dl2sCTToSH5V6Irngo6gytzB0La4KUWfIGYfLl7VQ
J/08DMGspyooiWYWdSC8004DUOJYIMRS+r7SyBHBBr5udpogwpjz6BqCq5UDjww+tr57jPdCE8Ca
KOg72qGpeiMEVIbwc3qTjEGRHQHwnqNd6YE7zaKJdUo3v8wIua1ae+MeDmMNNiTc2HrxwEgdNZnz
HHJ5/kzMCYImKTv4KvvZrYgQhf0TVMWFVdmbjx6lUP/MXYiPa13lACfTfXQF0lsEhPrMU8hzrqG7
iw/zSEsddOfSUUO+EcisiNAt2D0Q3xvzSNqg8BMcREsAIaZyPBi56J0Zc5600MGy6ehNuURX1EhX
pJ9jv+0iCg8yOI9SkfuC23vMWLMHX9ZMzQy5PAJb6WJRXXx4n196BTOnkpvvOulR5h24eSGZPR3r
Lc1Yw/AA6xo7NTds1XJI1ESXKUEvxn+ANmco8Rr9YWP1+Pnj1kP7TDHF5pY4paj7B2HdnBx3jf7Z
9KMXODDyq411bBgyh2lKvnIzk6dn8pDUdmYV7WWJE2P6PgTyQHPVSGIm7kuxT1V8Tn6196X/PaCW
/PmboeveR30Tc1qTngQGBiAJq5N42iJgrTMqA1/NYFuIzBLBwR9hrAfws6bWdDKwgV98BePGvPel
Vk6lWF6s0EfDEjTu1nmttV0QZLxYFC0utqKK0qnBfTKcjSkoti6hnyK6/XRsk2Zconsjx7lgUCY4
BlgdnZN8PpGo1m9gOurUyPHhb0Mi2fgtQV7SXatqu4p+Au6YCzAp01SOWnYF6mOIe1YjCOwbwgu6
qrcXXQ9YiphBV28AKXXUiQOcDwBk5B4T3GTprUBtAvL6lzCyyzRd9aUuGdU2Jda6CAqJgpUdYIYa
m1VasHTWWy6c9Ij39yqD9cSyZg2iGXk3IXIdWvCEUqzU3A+LutVL+S7CF6LEFi7Hfq/RCuJy1Qk0
MedOA2NfsR1lRT45746kUGJn4vxOsHXKnwCTGYN/x7IAbsaF9gwXoK+2F8wrmJbB+UtmL7QkrgJq
Ak2tMrLd38ruLCrXIfNwwthlRtkSdbu2aYuyUlJOoHsuhNCuJeRGhBD2cVzD5m9jbXuMV/yL60mY
3bcReLVOBmzd2F0ioL+T2RX4nWKWrdCTD6pTKIMpImUPCNcf9C4EepnLp9OmVDFgHiPCmSyLV27A
oto0OmuwoBKj87pEDaJ0kofAVVswIfquTMBKR5nfzY4SqzTR+XeI8wkZJMPKif8pBQ8fqi9W9mKH
nWxH14HB+L2QJUVC0i4ew1zD1TD0Lpfc19wcwIkB4xqY6rZbrxNhqHdjhnc2iRD1eKzo8nOZoa3n
mlvGd973On0BEDqtm1wIMyQx553ZSLFqZABYMtuW1Xf+rOKvyEoI7ElIdsevi4pWNiG90keSwhs5
ZDBHbxDLueuP9j0DMhuNjKYlf0DiDkCMWenoykUe924OmWebtQlKYiGXlfdU1sLjL6hDIuNUqyBL
H1n7XISxBS0PoJQVxTwSjeiGCgVgtqBIekV8eeOf9cbVfoQWCMw6ksTPmh0RXdoVGLmGQauna9xA
ti4aR26f/R1pJ7ywW+DQyGeoMpxrMceBjzw3ycnXOLFApyDTFh1PR/2zvjPr9y4joR3beGsujhT7
G9F9MgaoFn7ceB1qhlYAYGmNhp4pBwdJKqk2l1LD1dmocT+LdWuOWTIE5FMyCsV/NVdA433oat+1
ZEihPbOr3ViU4S5Zq00NMaTtvEXEGRWnUAcAvALn4f/jZkBP6RRWQ63g8V6fX4WFR+W4sADGOxz2
A2BJrYmW5arR4Q4zNTWWaQuUVvWhgy80sOZVduN3d+WSVUiq3iYzJ7Z7Qb+/Fr0n1kNz2CpW7/eI
XkVWEMU1oG2RksJodt8cFZbOaUBggESftXqODHxHLcdM/zhYBcz5vrVAMvmEyn3/aVdiR1Swxd6n
0wwMqw3m/ZQalV5jerx/tpSFP0wR8oePgLtw/AzV6jFDNpgyldC6dYeuPyzAv7tT+LhfDAbEtc3U
hOus5hOYbFTsQ5eOpvLTb9nktKnNZPo+RqBtGHbXqcSHkxtV/hd3wURYiabce2fyUj07UL62zPce
UtUxUW9G4QUX/HanmEqcQl6bDra//w+J3a0Rq0tOqBPe0lTIFag3V74mk84bz8hlV0Np/JbxiyqD
j/t3FrpV65+amxqgoEiEfowzTbv8wqYlCxmSiTOlg5BrqFzeYvECxxtrpRgWSetF80MOSVToFiWR
UkZnJyyoHgXKvUshmNaXhRqkQWtKK2QZ/CdF/1P3md/sZQIHVSJ9WRBM9cBRzgyXQVqE6NM0rCiB
lBYKtk38uPdN71a+KQHUZ7FiNLKiRl40BQQTfOiYcM7oOoxVYpI85aX3BPBmFE8xmDKx5PjCts5j
dWJTOaethEwQ031tKRIdk7zJd4Ds2DhFykjAI4bvAzJd5XChSq5PmEzr2Q5KyQKF7kdrWiYhJweH
W3lykMxQrL8jgxFZ9CH0Oedso2O4qeaBdX2XBYkyK+weWBqXeMtj2F8CVcJWQu3Rt80+sOGEKDEc
sDR71I0jB3iVdFjgjHeqqZVITD/7Ce4+EYeuq8nO/oE48c73g7IuCfFrxNx1i+a13DL9R2SlhZu2
goSMfch+E3zr7tBUnbr5fNGB3KX+Bi7yZbm0ZJYKMCo4vRAeVsjXCbEShpmfLeLO1XKGGHQui6Nm
WAqHDjsENuTJUnz3UH1Ci1XNjR1ecxun1Xa4+te+TVDz9lFEp8GJiCmxUkshArGinRw2MyuU4Vgr
ReW8QB3R+Ekm/1+rk5OHz3AJD3PDgzdtjXwkEXW4Pskk39X6yNKgjk1Brqzzr2W9bJ6FbFkR2Xp/
WsjdVbedzh8BmKd8ByasGRv2f6T8SsnwpihgrLWf2XZvZVf5EXVvTi63pxCzqqVoJi+qjqowDruj
AgQd1X24pMi+ZZQmN0uwgvkYf8GGN5qOYEzADotFZ88sSpMOsE4VznF3pWnURCOnUXjX3XiUMEWw
jeebpS+QTZnFcWgU/knxbNYzT+OpwMAjw3xtO06Ipfo0ldFVUSte3XvEmT4lAx/FfLkNcTUaMH/E
fZDDkHKZ2EC3yLdB3IKGVpYY1G/JjMRxWTnvStRqtg6QunNFYjNreupmfVF4yoKlF3wxMJ+KwBL0
rcVZQwsDLYNCqLiELkls7RZ95T/ZTcApj6CvcpYfVXsJLJN8Muv7kWkxnDE7aLo6sG3P+nXHDdVA
pqgosaUDp3qmf5HdrZ1wyl4F+G5fW3s/UFy4l/pVj4BaP2Ga8Ul9v4dQgTHRMOpIPunbA6zPzexp
RskOO0gzeJc+IA+witS1Y5D5aqke+QNOW4KzFFdJIo7qFKTcZvFvPLg4pv1bJJ1y9FtTrA52v3A4
seUQnkjp0lfRc+c4fUtP2rq0Kb439wnIUhRsbk/WYaEjzLsjz/5hmjShUZFPUFXxt2DTq3eU3Pcw
HZ4YQwS/Y6YEH/+TO/0WZ3GZUI7kudVnaX5vAZTSijUUF7BLNItnLn0MuJgQ/qs6qHETTGzfS2UO
HQ0MIZrrg7S6eJvE0rEbFNKZyapyORTdRSsDvTOpcEG7z5/a9j3DaOle0Knq+9fTLwcDacbrzcu7
0ywRDR5gbZNFJZQve3l9nY7k84F4VVhF6t/T6IM8IZaNJT71c+VkmpKu41/M2FzU/HmlyySwO97L
wb6sRmGUlx57UhPrKzc8of6O0B8JSRCKSL8Zrt3nuzfojKAvxqzE1554TA50sIxWn0LKTwXqPZj0
CFJe+OGmpYdEOGfs1p0zGphvflPod3DfPppLvqHOVaiW0M1jjIIsF6LNnkuFnaTILSZ32p/EpR7F
W/ECsvLp9+NaxaVeVAKjCJ8ZFfCgbbNSgdIDxebqv5xj10BmpS77OS0rMXqPeR9PoMmwQTr1jZUB
zLA9TNRCF/hQYoXycVV8SI2Vl9Obf873M1e1l3Ry7zdscaIUIsEuYarGFUZTTk91WpVjI/SV9qE0
XFXmATKPJi/Kwoy/+wRLTQLytVUWx/5HoYo91c19uQ1zNcgDU9LL76NkXRHTaUtvbxNSRGaBj7Lh
7C10WMI2lGnEQlYlMuuzCXMfRhlHgcxtYlqPyf5iABJAz8Sjr+UJ2lb8Ij7ZibFrnwWn9+5c/MO/
/T5NkWvq7V5WYSc5fQAKVKHL5e66KUApmRLza4FKUK+KCNVpjNAjvsqLvs2pq8HGuwqEuImiK28q
FbsxBTvTeHsVFYHSvGndHys5wJaS8pW4OhiX1fvWHQ1mm2nklaO0ou1dbxTkALoa60OSsHA1dbob
xNIRUB9UsrrRBlq76z1Ecw+QftXHVWQjgIIGZcPI94NF6BglW7flOPXDbA6o1yM1F6eNfllSZJrt
ME5zLw31SjLvRaPJblT43ZXC9VgkJsk7Rgv2v/VuZM93AsIl4gHfRvbOl5gEW8zG/ZmtXZVCk9zu
RibgTYVZBPnYzAaSm2aFuzaxXQKGmSx/BvsVOHinxuoDPJt7IyLve0U2unt6lfcfDhm8aYpNcylb
klXgK11VtesM/6HEPCsWMWrXWDOKLE8idH7L1B+HxCHE3nON1VxDp81+gpima0EtKKBwxBk5zyQ1
ari3j0SOCAiblbd54Y0H9iWgXi4Zp1fVfAdJq2DGdHqDewbALPe6FeYO9k45al7HjF0ooQF71WdT
xeNmJPGQrCNnaoWPgqHyHDBMd4K/DpFVuTpMpbowes6i9NaOsvgTouxh6Fq6ZxU/F2UP3MyVFMLA
k8m/3Zr8BFUoYXix/unike+49Xix1xaiR+TU5kqdwi5nC3Bv3A+0X57KRCazhUa1/Y7FbIhgcEda
CzyqVbhr5bQkuilGWxgV5V2WCpPfs8M36PsNuGeLfezHNXL+v6ykGHJmEs2AY/Nx3SWljSwqzNGL
tbV7VccRtkvn114FBEHwbUqcyNhjvQORR3RzHIChKrQWdtJV2JUbNyxyBHANnVFMsT3XHvvTmYXl
Rl27p/E9gk8XFumevzqw9F8Mv6BbyZ34vBOZa1qTZ7R+YdGYvdqhF0GPGL9YnKI+gePI0PSlDn5/
/OdRAtN7GVrjCNMuSq0RSJfz2vVzMUgzithXl9EFbGQ2sUcbo84MdamZfi0HoSA1Po+9XqZ2Q9EA
60nU+jcEDyL84C7wzag2nLmeRqMypWKG895egGYAZ2Nnxi3Cd1yqgAL4HNkz210a3pracmE7RSf7
3ngyjSiyFwQ404eKVodcdlcs7plkh1fsN0zugWVqbZwXZjTI5OMZ3EO3nYZw6jrixucesex0lgwZ
axXZtgODaBvT6wk7Mx4ahqaZN1e1fwD2QJ+ZcJ3/ib5ByUbF96g280Eb5ro+3+brfqfNNpZjxG2r
C18yBtU+Os3EHWNWI7lf8X/zgqszmxkFRX6ck8Sg8LKpSMqx9jOWz6N37KPZ9RHSBWgAcG6GocYy
x2oaf1GO1rK/4l03Chhj1XbPN5BzZEi/ef4M1sG6FaNA/OPb4f0JBilJ8kN3LMrv/wsxIII63FsG
z7rOb8rXSldiJFDwhTWHLKWHEEQ5oNcFFkn6XEhBtIKI7sVItCdS98QGHncMO0klnz2CTWo3Fkz3
5FNmZWjygn7O03O2tFQGXDlARSL5b87QOrdeshbcyDFv20YukUTek90/2EvHOkUlm8bkMZoQBnKV
+y5IjuTdBhraxz7g89AlesIJzllk/mpqdoXd8F+36Tlu+oye7LGg2uQh+aEvJD/eZoVLA42N+7XD
LssZtuQ2YMbL1nu48gQ2nJ1GKKR9jjPyRxoQDfDRdbM3Q3KZU+ESzxU4gsTSuOJmxTno9+xlucve
jllXg9bi50S2az3li32tucWfdt+YgHLSdGgoZTLnvaQakbXqNSd386MGQrueLJJ/5eYveV515uzA
vrP6oLtKoe6V1uwUqbo0m5m3S49J6xHTafzbr3rRfC1hAFhnsWuqqp+aP/4Z1RN6/+dSobWz+3px
bV19V5k0pGPgzNoX5YPenxLrfOJiMLI9nel9zOg+FvS3wI3bDFtzpuvgjQ+k1xqmwuOMok42pf2d
ygffY1DSUEKhjHXBYvPyB3jJ02v5pOTBxkztWgY2F0GI/cl4usdp4qvihbqHc71/ukKLJbTPhDNN
FYdMZlGHPQi/4lPxfsP1x6oS+mkgdNVMt3jQLGdG6aEIBqJG6QQbAaTvjhdNmrQF2tfPNTDvTY3j
5lEMCgrNOzRAG/izeVUHdOFAO/C8YtMqD/bBbyW6Rnr80qZjjx5T03z9a6jbbTTuU62P6Ks+kjbo
MvybRWBfGy8v2krPrjkab+xdMlcQcXDjltUAMKNSwUvojOVtYpHSb/LJeRsJSJ2AAMGCqQqZB4kZ
O5kCCz9pVOP2kf3H/eOU837EQ4DMZOvvJ/pcC15ouAlFm3FGzKqa244gsyZLhbkiJZpo8ihUrG/m
gZHhWeEshrQyfRwQKAP+0/vcbeQJZfAV1ZkY9GHt1MKG2jr52OgRqngRsxnR/kPnk/a74yXVC3B3
kLqtdE4/mWnPq8EowEmZUsfSw6nHUxoZsmTq10np6OA5GmyyPdWQk97G5PHe7b/UULawpE9gSsO3
rzWBmVAV/rYM89VVJe9t1DPgghc3L4A9Eu+7EoNvKe7eUkk46sqbvCq9s64BE9YENauoqHEVipNC
Gmta9ndDoboB0ebYAy4Oug4CpXjCYV+xAvqrvXxpmjDJkirSmftdvUT4lMt35Ia7zpycecErmQzF
eEopbtKm1we9VGlnzy9kCzIdtWoTiwlsDUaqhnqywkfWcIx+hGA81Txvg2V18h0M8l4GqTOfW77l
5c06O/J2HSk0RJavN386ef0/+W8wBJYKzY9t3pkWwOjV9L2ayAFtPviRD48lV5KmOFQ2gKAvM6t4
BWhG9wgpMkdZHhyWOQTHmfvyD5AoEzMEUQuE+TlPQ7bp9DIXj5rk9NSAnoWQUG+DdvMvKHRH+wLK
/oznDm+Jky24O7y3jKnlvpk100riXFkwOlQQW3VqWa+HgFrB33KaxjBaV9TOgsAah6ocKUY8spe3
BdzwapjKvfHp1TvkcOnQPcjJfeBdL35dIrT5HR2O4lbdf7kgPdzthkPH3gC+zTjc9I9jpS3V0usN
i9cGp/fIPLdHC62C9d1mLB7ce1h9LU/X4wA/53KLQxRHyplBPl0yhBzJzCZG0m+GNKpewL/TpvKr
a21bDqjSqlxNe7kbI2n3YRPwkBqJCDrf9okokRzaPXi5YTHCo/HRzI6jENf4SZO37AKubAM9CkTn
iQ0q9zu6JDROzDRGvC08tH8YH7gd3vu7QLvEZiqIrRndyvr328kjzZtNRA+dL1/7m8QjC3fDdShp
0azpBw4hzQelGtcexm4CgmT4kmaeQamQIvPgVMhyPfF9FzQGQXSLZqz4MDsq0D/8ZAyESuclOnZm
Jrf1e18Lx5s2IHvtDHlBj/vvKRNELCrhZqnbcrJZikhLppsw4pVruWCxdrs8672Y8YtHaJiDAF5+
LaUIyQyRj3bcJTGJQyVDVTk0uY3ckYAqPTQfS9lI74ElzAUGRDI7mPEodalfleAdZURmJQUf+Z3B
QKa6dhDrnxCcHZIptSiiTDzAcpr3M8+imHTNhQbRbDzjwmtcuj5NKIxYbX3YOyUW4m1Sl76Kce55
9pde7m0Algc2HOdu2vYdAknpdG7Ev/0PEKSk274vj4I/A0/mz7cfYYk+MTepjCSkgMxuuiTYGfOF
L1FTviwC3Rcs+dvVDwS4DjcGc4k0m1CGU3mnN+k9vBQxPpGwiLn+rzKpHvwBKlUN3/oX2Oj99q4q
PWKG1rhHdFH5B3/aNTBhgrlVvuKzFP1aiPmFG4SGdBlUa7nrflONiwn07nT9hLRNsXZOR4+TkXdt
sx0V0wy027w0ddDiYyW2E4qi/Ytw77p5DG80EW2XTdXMvputWtoCGsyFCvW8k3IlwUqizSKC7QXA
5YpiuGKaM2zorvys6XyGQ/xvQ1vyvblB4fDIB1u8owUcwaxM/zJmcxBP3MeC0lS+aw2i0lo63wFo
LJMvrfA1Vq9uB4BlTNuO+brHHRpUZuhhQ8s+h1tX2EQix7isrCyaMU/DUR+GtKAPNmVm2KDe2ZDD
HNDpHogJIXOZPjtXy84SCwphjvtOd825VMTbEzvSK4cC01tlwoO3Rq9VyqpPtAiL++EXVw7w7DuE
vv6QWMxyTzc9EUGj5z5tVFogq1qK10e9gJNbZkovLGuhlVvR7NpPm3eZjyo2QoqLvH4A00wz+r4j
JdJgLwOCTz4tUNa+AV9Ez1geVlOKQlFqmY19mjZhfOBcBcyPmxQjAiBGblQCQ2O3Ff1GuKx1fuU7
jbWged1DBSKD9l0aFZbufVUF9AVN+Qz0t95zDiD2ce6HSz6Ir9PoGOfh97WMUBIQH/vUS5v9VRJM
xSAGaQUOR4YXxc3k+O1zSG8TAGva4Js0hVupWoEJfklMbkyijkvPDdPGsY3jeAZaTlnaLz5XRQen
aIrhjVVtL0lOipCrAPE5di4eVL/ZvBifIRCRDTSC8Yadu9d2LzWwotRgSHljaBgUUzYbEA61pAGo
BFDQRKRH4vWVCzqOUsEDXtgVsFeWP/WNnAWgbZ80OpKWkX8sVIeia8yWIlp0ai3XsnCauDPA0FKY
0H+rZzTXUpKAhOv1tcWy8DChsxwOe2Mkxm618NW4fwm03gNtdxmUuw7kMgAXl4tQujQbr96sEGn3
1O+v+FyAq2dhJHNAwDyXoDmabDcG69n00GETriRh1uLaLD80mjEgzmGU9C1p3nikeYjx1NwR/KNI
Iv+4Ut3hrFbSa4CNdHmALNd4ML3D9mI7AIPc0glXMO1Ep62+RlsTT0HErPV5us5maKOgoyghxylB
RyDsrYLYFrRvZGttO84AXVEErTc8KsnzdhoNcFMJvWj0wVo6/TE5rERW9CLIg3edJArl3Czaz1p4
Q9IbRmyM9OfoBhl8i2Dug4BUfupeJKddwkOszJs2WLKWhQJIbiOakIdf27Lo1iDRUjE+eLOBJjb2
25x3gtlo3nrqVsQ3SL7wC7yIZEdlE9CWFPrbkVQoPNLQCy6Tf+d9QiDkDUi66cML7OqZubXNtu14
v9+v2mjJZGrsCBpXLz13yD1GEHoh8AjTU3/TwuoF2huZuYEKfdiiCFJZ53kbmwjUB4jaGj3V9m5W
WzXJMOY+TmbsphM2SVNCow3t/YnZalIeZvxTRM3c4dbC33qcs3N1SbIib28EXd4s9TdypbgivFT0
yIS3z6e4SSsIGMMnYqAiPuoi8tCvfbsfoB+7CeeiafZRpesHlOdLckgMKOt6qew8FpnM+jDOhJQE
6EiMRPv7d4ba82abHF/FMKTJCGSqqxJMF4faPOdPKnLxdo+qOWNiK98lbk6U47PWONlQqjm5HsJp
n5ja8lLTre00VfItOSyBG4HxUKpRBt0vtV3k4IpTQkR3RFd+Y4Hhiqt0Jcq8xNUb+MnmjrV5vaaG
otnrxaKvK1AqpwGL/K7JoAoY+/QdaK+yYKb2s2ANr/fn2spE532Wrk5QnNRNmAQFBHia5pNmm+iX
qAVVfBFcIo8NdfPdteTB8u2Op0eRvFOfFiHKj0rNRauk9gjjpn61ZcoM5XH4xkbwDjbdh7UOJoTd
kmB6h9okhD7vPpZhh3BPJpQYsrfyTW7Mw8c2BcXpWZF/8weYEfaq81L03s/BjRNFX3Rj4GFpKaT6
RlF8Ya5jK4cWBWsb7SMm8D0ggA5EXELI7+ARKWoPjugorow7GCHqYbffYsZwU1pSS+/iLsi+29BB
mk08j4hG4sk4EEJwOKfN4lg37W9Ak9ynDFZkBI6uPE2/K90LYV2H2MstelDQxr0Gw2+uTDTMqEnP
jEYIk+gFKPcSwxCwZTjss89TeAeud4B0O4SAZeAoZR5rmPF9ZuEFJujIulUUHYm5HfFZCeBJhsmW
Lj6xRi3imGgKhTpu5DFAaGUoy082BPKyqpDHYNhxc8TbRz6jevpK8f9VtT1FvDF2qFperq89ObWn
iRa79nrwcV1Avrsgd0RyFucbKBNy7ubopCoWDEpTReF8c4/+JT5qVFLbxyK7Mp6x2xb9atYxKFjQ
bHo+Uq3ystvzIeuhAB0kfmBk/d0apzTW8cYKQhnmsrGzC0FcMnksw3ZgycTNCMpACs9ysOIlrc06
9TrNBC+i4WFvAm/A8XamH4ZZGiVSrDkFZ6sA9gpkNzawGR9cKw6DqwKKVgCBSkKCGEUbrxz14taN
hLbkuzt3gM5tnd17uMcoFnTVMEjpWKhvrfPx9f8v4SafmlQ7PgjwXF4vkiyu8YraBbvxJ5eO/1u8
YClUqZQUOYyNV78KyYoLuwUjanratfQUfaWNPhJN1zy8JVQDt0/iJ4b7iFImkpuvHgYIQeR15QHx
HR9NbT9Suirg1ItTTjL0cqe/NE6poHcPtYk7YZnAhCq/iTeeMkumS/lr3Fnr9nxYhby4R+aDcb2m
b/ADBWU3OdAUS1FLoBvxvwsWGpoWHpeek43fr1ndHx+kJ0Rw5Kwv0hLerQzFcteM1d90Gcad8/MP
adoyfiGEcldOYGCnIFWEoyFTbwR/rNATjNfrz75L9pBgbjaKH5iGmn1Dn9pKyxMxN2SjBOqWIdT2
qbfVlShXk91iAjVRr046mkypMh4wiKGJXA/rHPOJoEJQ9W/IbknPLOshXv1YbMvLR1FC5A0qQP1h
F3NK0jWEmbzZYjNlz57PNY/Jj/8BNoTBpzFVGk17YvucSXiVMDD4SrpcGKr04NVVpVEGwgjy0WBL
5H/uNKsRKNJsHE68IZTgY0yygeP81eCjtXd81oLYe1iIZSnGqwUrYvsSiBACKvA5TafJg8Yx/2zi
UNOvSBEM1yLgvLqtM1YDDatGi+6zy5NJEHjlr8kprwCLu63dokA0GVlO0kR0kzXACNMoeNwHOFMy
6uqPkkuXhgeceic34masdzlPv/thOg88hlEAB4lbb7Og7qrDDiejqEK9Aw69oVYNAYtYejMcfOUN
ltBUv+zu0WU9/DEaxXwYqAGTW+QqETSq1hdnelBglY0Wefb8FVAMuNTj4r24AmUgtQHaT9QYA5PR
rXetXhk9+sqbFzXxAK+0R5MqGDJTtmEpCML9OMXPJjJX0E3/+zTPxQHU+PBKoZ9D4kuKjFvg8OYh
nmmkOwBmVrd+mE6k6zPq5uCj6rjaWYBJrNUYV6QND21YSlPi3o1KToFcajfxxi/yMYO7FKkKGrLy
aknNRUs9CkdASnKkchUVmVAOlQQNpwuKk5FaYg5k7EE8Ro8DXjE7b95kF8d2DtvUdeBx8TtxcQYk
8bfw2n3gE5j0I391MUsBDsB/D2WF3NP/KbnyckT4PS4D89sQ/nTxDvnbieCPCeG1lnjj/V7sN4bu
cblQrTsC+kE4aRJyrqDSCKp0MA0OgAz4uLOSdwH2yQkNwhWaCzfM6rQyD8t0LaDc6585Gc9Ao06Q
IhiDE1HqLf1EA3Ul62CCfYoQ9PX8gZYuXseFd7LgC3Hpb6bKQf83JErYDLV1WFSjKT0llB1D55Kv
cFolSIK2FX+oqo8lIjIdPWNmjyNY0WV5D0SNK9/d8ERn2TrZ5T6RmfCfeYjQi43h9x5sCTFGyZRv
cymRNGK97baPLtLi7ehCPnhjb0DlKPbDVOKXCHZ+kPe4MHmCwqqChHt2W3QLs//KH58nwIaXqM/w
DunlwNa3ZHkwSVxLB5U5VofQPR4FR50iCMDe9CO4ib6791Nt27B+Woe9vUNYsMVjYrOPi0JYkifM
YGDOAf60/4eBQD/rokMQ32JR8EAhZY/8VqpCaeT8hirmTLnOS8KVP1nJ0RrHxloxZNMg3GH0hy03
hA9ZY+gQS0RGQH3uiLysR0j8k+nvORs+eIzgqv7906EEpgAVsbnXI6gXk6nhQ/xP0sf8E8YkrMjM
cEx7uKBIQ4DIXlx3MGnApsakJXvTM6qUlioyxpNUblaBlDpvkEPpSWlQHQtneyTIS1ozycgg6KCh
dLFzpcoUQSkmKkZOdmqOfd9fNz7CnPbmbHhKAAfnylV+AhCPH5V7nkOMxUOey6gdvSVIYg9q/xtx
n28VLPzGlJRGKIkMxtr/5IbIQIUPbsCEO+elzlnsg1XKx6wvZ9LzMWnL99TACG4Z8CuVe6OcdvZo
xN2Tmq/i
`protect end_protected

