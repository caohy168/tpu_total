

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kPMKaDOi2kQXuMCKSdPBKatSDEqsZbq8dJQr4x1jAazoyE/zREc1R5J/FG8XDiEZQa8nw9j1ix5C
oQvQGXZKrg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qLeApUbY8ZXxl+1uDLQ1NsEgbqOrFXLgNDRZCtdy+tuQcsXM0AJiWUKY75eR+midgoNqD6w7EInO
ie3/tp8VrUrbZ004xy4XoAS9xgxtpDK7zidDI9umrl7fJtjyo9eyTv2JnFiF3g+9pTZrylMG9cyL
Jqdjnq4+UcuchR7QuMU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xnQyIQHzqLl8QgvKsIJHNSu65sa3bd65FP8/+jBDrvhjpx3AFd+fwTGyhqEGg0LLO02WqW6Apap4
SZrmb9BVlAXKAX2FpWv8ZQS2DyptBZUqKJelwSN1W0GK4SL3Aypfzg2EBF5/q/OFQ6+flxptDiNG
EnKZiLXMdX/1J4Tj+1tjCxDXDYaw07o/YKctzqbqesbUOb1O9e5Pzhq+fA4LTgW/YQfuObYcctm3
liRmYnsg0glfs40T1YlZuMnsG3VLcf6TA8Qd5w9qhSCFabAAalfNy1QkOkm6l1gqJnS7k4Du1tkw
MlgEyUV09+sefXYVTQAkq54DH5v2E4QzMjJFjw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
USCdJYK3gibHILCG3SZ3rb4rlPe1EhirdeqNsVg9b6Mgq3qJKWqbBaAuKwIjo+Tn4o1pD2pgrckC
cOQ5ofiFQuZJojzr4wwMCwaBuvhfgI/ph4zv8ccFi5qVRkYlJ3TIQmkJumbPP2t+QDoJJvghELjB
psgLGLrk1uXjPvrZ+AwGtIKiK3PQ+76zch26VX2KNbVfzFf+zQYvdp5Ucf0updVTApLbEt61HHIS
IEPPXDO5Oi73S0kZCDAXxHz4AGX/EQlNMwb+ddqAkYTcqY9FaWy3GrnMD3fuB8LtD3O9he0eZtEy
n+YGhLUj+NxpBXpKOMPjHH2MeRRn+cJVH4/Qzw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fw2Ueu/tNez3Yov9HXY5IljhQKemjDQX3jbPt9ijSgyTaMBDw5Kw9OGOvX/39JbYv7R2dcGbAP1P
/kWEmSQMBA89GmYeaTGGt+Y83GnY/mt6zlTgS8D/ZCCbHHXw+qlNNrVhfSARjlSKhj6VppGZWZl0
Z/9z38jibEwD7vn6lrW+ir//DI6BfUjYTBLXmYfppC3D2/3udy24bIFP0hfmY9zgR3bc2D1Rl5r/
6waaZQkK4WwH5lKNGqHdDOUvySiNCfY2eI6+parBeBu09U84j3/aBmgL4A31Hh+KVxmFG2CmPiSo
lrYFDLXO73zRYbDZ8IBU+S8cPzXrNNuT1Th2xg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b2uOQkA0sbcvZoGixYW/raDVvukcDKw22dxp5j7Mw3my0is9Uc9JMBTxHWTVCo54sL9pMpsNrr+1
9P2QNefar7dewJDfc6VsUYsuwZvpLkPtPyKJdFmhbq0tfQ2vaHAr51xPIRE8hjeIhAqGu+hpa34T
PFAblWc4afnyp+kRycw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nRBwi3FFmJ/6tXhRn1YPnZ+j7GNxvO548dGI8tBZq7sGV2oYbdspjCmXgEAGFMB6Gn7qV66rW8HW
i+8pOmwhY0+xr14RuwYVh1ued31kJp71+NEFBpoQTta7c+m1PwuinGxE1dVA30y6W5BpysFvceHu
kjixM0ey4iqe65QrViOc3aFMoQkyNG1jDnNPVU++7Gz4W2wPb/sQxTeN2+p9uYz/OZtk3mEbAXeT
wLx8I93uc83hkZCsbBWkiLx5skHPnhGWD3izNSDLaScE+bSw8hwv91RMtLF/x/xcSN5xZmWuZvHg
m5Lvl+vMZFztzpt6D06wDkAlLioGDe9TeEzkiA==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SvCVHEI+mCgtjsQ6p8gRD5V9avjftzeQS4O0q+g/VoNHuvya7RUs9btiXNIkrRJFV5Aj1b2G4lYB
F8F4jkkU3JCdC9kJt5bAYq61b/I1sy47P+BrX4VfWtcwv0ZU1u+hliYNLweMc4nBjnMLai9JMFHi
tq1VxNnMGx3tC82dfRlYCXwZt9H9Gzr4QFVY0NH6dgHUeIr09XKALiJq2xoTckJ4cEosT4gQrjwh
JzehJm3/WLtM+ga7ihKtNttmvr4EuWqJV5Ts3CwI8No1ulolCG0+PaZjXyXaAPYs6b6+HJS8xB/B
JnUQ/C6VU4hJXwTNp30KrUn5Zx3ag5/n/nKodw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121872)
`protect data_block
ldhXRqn8TZQkFRALxV4lXnJGyO55nd4d45WoG9BMyZy1mTwxHTFp9zT5dnOCpLpqofkibAvEeTH8
r8WnmYfAJ27LQvwZwkTiWpTeoHx4X/Z+XGd6jjqCjfsYfs693KvVaGCflP04/Dz3U3VDCyBM3laX
K7gEFQWs95TpCDzVZzA5caPJKo8pL48gMDit441tyYZoBUt98PBTbZSrZQ2Sgaw0biiPm6ctpnzD
Ax8j4A1uJw9iESXFSpO4HASR6OZgY01OrVge3EqafgDA2vOzjpTbVZ/k1NPWlZ00HfFUIm6xR4rr
sYYdF875MZH3xcXxIk5GupyjO3OL6bciSnnRQJlQtDksDNh9feD5ur8mYGAKZOYSHchInBK7hAG5
QxESPBriK0suNbhgpSwpob6XqI5EtYQzcfs9QiykrFYSoCJQmb5Zod+vFLV7YfnHKSDKSZX7k86W
+EhWkLz8FbpiUMjJYIG3b81933OY7E4+LT5DBuCN9jVoAyxsOFKLpK6KujacXn/Bu16IPmYIUhXx
rLctAj9cnxr/eipmku+ig2TuUCTKHbkoeAkSJ28SC6YFTYyN4GZaDSHmoQoUyWKWT372lI0cG3I/
PoJ+UAnU0ycQyo6XUBnvjBGq3AcbOrxyjmza0GsvdkFNP9ZBqzyibWxJFRX4wWcL6QqjOIK6PbCN
9SvK6u4ZQ3NTCxl/G9Vo5J6eZfL+MdbAl9XNXnE24Da6Urmgk8zIpLqKybrjblw5zgQFtABnhdvM
AwBKL7ZBv/AG5HnWOVJ2+gRQlvGGeRE1A8pikvn7rotOu+SryVtWcgYW5qG/qXJESyxTmhMKwzSj
zg6GS+TH6v+2LGkewmF1EOj+sGpiLKtNoi66UQwS3LT511g8JCj8cxvHdtFYGGdm4yEOlKoggvIX
ZL9P7urtq6SCL5j0HhczFX/vT2oFENKhC1A33wOGAlyrRNq5ZQeCkd5uo2YH7my4PjWzREsZd8Az
YJCDhH9QR8HgmPbq9ZwNApKivToi/HTlxDelLr7uJIzkwa9ghUwxdeq1EQeNkOvrMqda3r0WPv8s
J4HgCEjvEFRJLGsLRnmo92L+VcEBn+oDi0s7O4GYrs8KUZy4uwRvhdt6Fd4YdVpZCKbyT01XBMew
MqTtP58549NV0mDqVcehTOysHVs1htirYZWBmbTm3zkfvCpRa0rd3+Zu8wW/vBuNh8XUtxc17Ikx
r50uhNhU+qhuN2ZYbFZ8q4mc45K+B1PvnSgUKYhj3X8AxhoAwjOscIViP82ApF3OWQlPnsXTByde
mXkqdT90Z7lneGgoyWpB2erJJI4lk0Q6RYd9NP0U2zFosL1KTivy4x1+MZi+g4uqRjWCVo6lqN8U
AtFu/8r8llZmvbmo2toHwDKjJbfjKqhVVWyjn3J/kLgcoxMCpE1zB1eyJvkyC4wVFh+SBCIVzbMA
70x8e34pp7qq1wkHsY8/UbABRtyp9oTUCrJ9NHg90UCCV9bUSttVh9rPl45ABSgBdyfXfghWWvim
l8WwuvsHnZcEmWpHhXBLRWXTFI1atrzSRX8sEJQa7cv+F2Lsbc7N2m4IC1mGM+Rj7fIOR7ZQJ450
+XrPJd+7mOTFXf6+kU1Fg62A/ODmvpBgcnODxCZH6GLtsgBMuopdVObTcWiST5/z98ltz9+wsXlt
whcEKStMNh+8Z+JrZ1Hekoepri90m7c3SKsQ3iRUH2cWSpTB4YojvOWUdAdc9dAF0X2ef4YrbtXk
9GcLv3LJtbS80z5AO4lzHlt9B3UJ7wml7t5tXrb+qC/Ks2HVdVzbXps+nB/jpQ9nLNHYUN47Im7u
HLNH5IZPSPZI9N0GB/WfvNfjs+jQjR/OLQlQQFigs1+5Q5AolexgceJuLjhsU/2HQcxmysQj1mtI
hu46RCBu/26Jd6SDmEH8PAi3/gpbD9nR9gA9URk47mU3QS6UIIdBV21HH697c1vU8ZM+rbIG8hrw
HQJk3LaRayZsgPpSoEEa4aeKHXP4OzvBTAambKelUzoRMEM8Se/47toDu9IT54IHLPtmRdAUJQDZ
PdetgysZshEzCnM8rt2IcStMAzXpY2YiMruXA4DavlB4DVm27Jj3PEQ2HJFgiscZpXfxK0p+2ta7
2lCC1vX+xIqV49N31lOsWFbqTM3eFXAPdlELx7gX4yoCYNhxwTbdFskaThf2L7fR20byiOODJGjf
snkLPFf+uCJPT2Ro1ZWfdR0J7CnT9bf79jAjcfpD3OtxTzqE8qcZveIn98VWNC4NAWtBSIttER+w
pFvc2XLv9xBkvbWjTntuxkSGMPk5RKT+bkjS0mIDIPEaNQxti8v21MkL07vIlq70XrI2Hek9+GmD
t43/rI2CduquUW+XAGtVfbuc7oMQFmpuhlIjVL1VOJfBCR3l2/ZR+ebtpOwZm05DTZp31wJ37D8u
SEEcysjkkDSBiQI6/uCcxzDfVrkIkFW5283EtsWfLa+bke84pbqFFfmSKtctYwqonH4P/2wDD2PC
QKFfOK4ChwBk8a7m+QgJYFjKcBGF2IWgP0e9xz8M31MXd2U4OphpNSH5sAPHDLXK5mn4TT4chCVs
4l06N+Fj2fnUqcb9L6w3ZRVr9DvXi5KwHKfMipuBMRfscvw94jJlieYl81pc7qVMBIP398TxQgS5
DLK029C3TB9u76rUS1H8CYDfDp+R2BUMcq+yPfdNHca+hFZCjmwN24VEGZwp+thkRKHZBQu+6U9i
7OdwdoAjDVCkgZDBQCWyGDlb8RDG6Rh5drXcNo/Gqr0ac4mZhk6HO/HPSg7QHLyhDD5joSpUE4R9
daRRfZlUtFY1j7RgbUd0e6PIeQcSCZLCwh2eUAttBOdobLVcOeLkVSbuNt7htHABjfp0Ks9JA3hN
1k84N/hiKaA+tELb32uiSppFqqXY/aOnsfhdrj1lQioGENDbC5vZiSIp6DzCC0tAm+4F3yd3t1o7
4aauVrMqP/wZjOxioHVKjIAIxDnssw8qea59hj22/pGXR8xn2o6AgYSALwfwIFmbmZst9hK9U09Y
qaTKwRN6nAQka3EteqgabQDBkSg/IXZi8F7JZA3D87vzbTJuEc+oTbC6V3RpjPh3ViotDcHvQKQ3
Zh76qs1tHSjQNOuNgu47Ih5oJmWx3iDmefKhgdq/E9LBe0yKczWlGB1evomI1EkS6xF6j/uY/vbG
UHa4yEi+MpbBKUihkaRF89YZNBi+PcNWHkuM2gzKNSq86FfRvGddYdI7XIK6TeZf+IRCU5K+ulrp
BqJQDllVdfWN/zL38lhfbrOlIA8wjdVZf6HAnJojOWjY+6gkHrZsl6lLqrOTiDCx5c56HY3318xA
ZsMjKIVLL/z6X3047lKpdRSHD9wJYg/jZ4UYha1PuSFGSxOaUfK8Vs5uZwu2+D9TbaZ2K4woYo4s
Ku8X/ZYUZCyy1vcsiQiqNAIplKjmLOCwrlP4F6UhsSVv/LYu6IvHql4W6tO0AQYIkI+1EY2kwkkC
mx+P6RSQKz9KndiQ2KcSoEklyoYQpkwaRqznaAz1CYQPwngL+Vyj2VZfp3B78RKdJgw7vCPZd3Hl
xC1mtiqiLV76LJ9DOADM5qsD4s/VkJoiBgskSTmCb9rh8rKjrs7JGdJaHmf0YHCoFsVt/m0Rl0YM
hxltbKc0sVwE8xRBtQrLwcQhI052RXbdIzvQ8vKdrUJt9L6sg//Kh8XBu6xYvlflJlIkifgLlCta
Djul99wTjK/nryixvb9drTT9XqQkW3IF05apzSD+IzA3zY+oqUix9kZ7JsqnWhGVR84XbeF5CRVX
aY62akdRTAa8hnbHDE/6uOvEtKzTEevgIXcQpA4dQgtPzvaV4YwlacpMj1FYaM0fE5sFW4sOgb37
orbiXbfn1D2c8iACQvBdlB5EGyGPGXmLKMz2JMcVRrk5mXeZzS19N3QRBKAZeg4a2UTJYy0sFzTh
akhRd+mtEF5OI8B1ggmsovrOGyqdrLQVY0GehREtmG0i6IeGlenRqV7Ah0x85n0jhfPP+DVPXVb4
qS6Q2VI3neJu2XsBqDj62NVCjcrkx076BnYpgOH5Gc7J0QrddHV8h7tVdnFWd1Pt6+F3xTmKuYK6
fPeZF2clOi22KKxaQDe90ccxbVcq8Jwxt9G/PPD+37AvAya5SF0lJe3pb20oyyNbdZw3pTVoVE06
AoJXr9sHMe1UnPkpprSLFVJL47GH8p7BlUz11nrgJ1Yu6rXsPCvaZMoqGe3ce/x8Gu+NsI47Q1TX
QXWWRRgYCkQ2u0wkV+egxvYfq7id1uR6325g7/4Nn3+aLvFTOD1QN2xFCBHwz57CO8QHqSh5jaUq
RcRhAFrjBbG7NeXIlZkJ/1Ayz8qgJGmwZ1UuF9avSr6b87pu1FucdyikCfTfK2XRP40tqfR/bEHX
gHo4GqHInkuld9Oo78KJa/2s6odSHSj9au/vdYrUsbrwwEFP2nEUza5gYYVy23KSuCOljuQ0VupZ
n9tK/5oYwvzH9oCg6QlKQxLWDzHqeNQ8/M00v4J2oH7u2GY8SE0isvEev+oaQzFsRI+j2Ea2nK/S
RaTqkJsbHqD4uaQ/r9vOGthAnuRi1rzAVexSVfJBU+DCknJAshC+ErUGmyYkegragoZxd3nXzlNm
FPW4tpFzloNa8FCLrwoXVx9ds9NBblxLix00UM4kyEyXBMHdsHspCemEPJ9A4B0C3jbtwU4xAcyH
j7IPMQKgsjWTMfofn6okLwOYIpbdJ0JqBXRkN3PKMzZUE8jAjUoGjSQjd5N2rHDcDaVfkL+5yBXd
UqMfTQCMqXj19fFx3cJ4fH6wGhj/69s5vBM7NgIbRqQXPj7TH+CAZm9tXQfP1CMC7c8ikVOGxNWb
bIMIVy+8lwIpYElGwwQZqgt7oZtbgtoW8NiG5N8ot4ncfJE0edtnZEyaN5nS4tQc8n9Lf078dPVB
K5MA+/3WrsPHwGN/h64W7P6z7+IBdfFLAh2DuHttjkFk4NplQZwSUwUBYJ0q3nQv7OGzsfUO7cbr
a74kFuQL2GVpIL1TzUCcBu3wx0/ulgzJOcxTooU1TtYmJkYvh+zRjUF53cwnNv6UHvsbkjdCEZBB
Z132c7HkjpL1E9w3pbDIY1j+VYqDA4kDVi8Tj2ROVb0/7mGNCcMRnMuDh3JGEpiXp88zRnEN+Hwf
R3VeSyL/+rWcOV5amdmgeFPiEbIIZUhYDQsra5/qSNm7rScpc9BZjvaJFsaCXvrK6yX34qF4A+iB
6VSXJT4W6KJ3vmSA/5gTNe6vbjT/M0A+y5vlizXwk5xFM+FWH5jGB+DLTTC3BorqwsmIlnpWiMAf
o+88GaAfkcAsKUUR2zDX+cEUML9i/HyAYZTZahTcT2NcP3WMyhNXOGthNwqWHutiLcuC7pVFgRvG
lMNXj4h2bYcBjdFjn/MMXJCTaU7u0bPHwLeBwE7MyQVwQ9LNHQZtrZyKM7d9n5loY7MZA1b4HXMm
Y0Rd5gnDs0p8Z09SlA+4fC9ffmxK9UyVvlqcG6IRmpWk794dZlfYrHFKwbmSpE7mjxgFDT0XMQsz
H4cLrNXWItbRn5o4yjp2ZNpAMDwfWzqhYq4zg9I6+qtuP8HQdBfItffwYaFTIYN73sTCrIN1Z0Mq
g3egKV43/zdp6dYgM0LItyUyDdULKWNerUiDXrOruULc2kYAa6OV9syEFZiZSBcIJT4YdlOVsnKo
BOVz8pzh0X5FSYp3OMZJdc1K+sbgR0p5M+kh40vZasOy/9DLBOoU6mZ859czoOBinfvc43ZFS785
bvVqem6y2UOB/5i09ggQCSyYcWKvbCYyT9lT03CwGplX5bPNfFMjmmRSRpVFYb9aJhUQQazW0orZ
bkEEr9Zl7y6poqRONfdWmroWCay6iMQk7mdzWInZzQyHSktZbJFDOAUxw0SlTvL06ZKCuViAK+fd
pTqTqRN7YVvqJeznaLT1GGWiiR/2Z29SmEh4y+CrIYW0z3EQR+cTUdTmDEy6JHoBZDvStMsWalfX
woeJLAT6+h1STNRzLx/06A7g/NPZv3Lhgrnpa+uikjTric/fhOM43NUwISkyYot46VAdVuisUrGu
gsE/ady422YY8tf0t8oBmmq4q+UVfiuG004eF+nM7VwoXDoE1FitpmvFNfMdGugjaW2Bi6XRKB2D
rtMtSTpYxBPlP1kFOBD8MDwdpB0GTG/vFcNfQLgPzqMbsdwkrYMP6CQwsYP8taEzeSmcK4BfD0SX
CZiuHUqXshVGZYOruXFeHAD7oBWlY8wzceNGFB1FpUMVkBSrDARMiF3RDM7/WuevW3JI8Tcl5irk
+RQPVVDOEOHi2JeBRbHpVfjT/L5izMhv4qnyy95/jaqhtM4c948D5X9vXzzX7GD7XOAYutclVtOv
1BtUxiLwj3Ba+C2iY2u6uwM33UPihIg9fJ9ThC1mRi1et97+YDaPkJl2zEZnP7xMu7ZtZ98zoUB2
yYxGC4U3ACOTNFhjpHG1GenhNhoioGkxPeuWh8Plat/A4+hr452FvEqAAHFinLAgzDWb+rZvR5cY
NF62VLP/1erju2YpWVlADxOfuMr/Fe4SqLGk4pmXONT7hz56qGZh9JcOiDhwLUcrVt3okRJyQmeU
cdSgPtQQGB5gTub34jTnGrUIUm/RMQEVYRYWcKubWruou9d56DGCMetXU/XwXvWRID7En0KQJyHW
Ft6FRQ0T90atnVhDaK7ymdG2ZGANmx5K9VerKT8oBEm3unLDAxba1C9GLOM8EmrhGNzvLwJTDfCo
sHmZAuA/+6jYCCfAZdcg9W59VHoxobURgEjvS6jJjSzK5ejWzQ05yNmF6jKMh0jACo1zI4Frki97
yVRHnMnWjE4mTl5qQC3Y+60nSlOQ1iVEmeJXNgi/j89s5TqmOmIkEWDshSXVh2So9+eScUBzREJ0
jLwfmOdd2U3QXlWdADNafqA5FP+kcPmsKsH1BJ8Mulvt4Ny3nCLnowVxlm3w0NMQJg9ghGn+PPER
lej4V/ijTRSGz/RzG+twtpthFU+Xz3GM7Jzbo4SRWqCvfmf1TGDThR+Eqakw8QfCeQjJK94wpdQq
1FLr4BdAmje7+LXez8hgJFBMej2L5BEchHTnFs6AZUZ1/UGGbigcR3QNq1JeekkmPniR8nI9U1jK
M59xQ9I8Nn216RX68s9PF00JVEMp5sYkF6/cLGk0CS5dIkbGwoKXS8gSKlhaqNCXfKtm/SxPOUXA
Sx0C8vrTQ4yZ2KQNDV5N/fFj+jRr1gZHf2oBakvB/lGGILY4bIKj6w7J+1zp/nxcw29wH813eK4c
NJgPfS+gupQduElHvvhjvneWunHw4NvZpKXf8/VuNcroiDZi5gX11iUfEfM6+Iq438/yPmQC+N2u
oUxK1akFctOMEuydv2ebMwdTnWK66hj9NvXvgy9ldyFlKpLlO+c7+zYKGHqUl3yhTQHQ/Regdeuo
ODE2V5Oi6BZ+5FQbrthZqqJ6ty/Mhvt7T5XAT2Yw3wwM1J2azBKHKnXrpY+qx7IOo611R12/DTzX
L9Y37DmZLZGS+4LyLgFSBHIH9CdUL2c0AL74QvKrW2x5s7I9Z2ak0iVUWYDz7uUd/5XD3OzEJezd
WK7uvWQUajOYLpGi5Kv0e2e14zSP6BuiGm6ztGweWgR64NIKNJBwKV4v6Dq5hmak785UASU4kEhj
NjDCfS/laXOUBYubCkQo1sIfO/hWhTH2B5YsuGgXK5JnsCbj8FQ5bKbkKC0Ne6ibzdDYT8DGqZQF
diQxiYDXAvZi+d8xrNyo8WHYHZQHXaPaeVkx8FRaIqv0Vi+Fo+hCbSOhyNvTOTjI3yAVYR0DAVNO
o1PMOrJhuvRaj+NtsDGlZQjg7slOrtg0uOLW1lWrghdRyFJbmwMqtqHtySXpm8pSsjpunBhI8rg9
XyntMx2Dk7HSWxcFsVqxTPVaksfuefot102VnPJzhBOdHS3pnrEhwtdzIT+gY0TYyB6e6zMXgO1k
ZoQpln1OJ19vYr8J4To2cOOWuySN8wQqz1KFgElEIbbW3WTXmeMewwihqgtNj3qvC/IXFpi2KWMU
LfziaShY6a/aNAJYbJvyx1k8siecdhtfP/J43OBCSDbFUQWcBD5fp67BcdjMYTpGTPqxhb8GUlXA
bTkEU0zhESqu1hzq8ae61ZSdGVNl/z+MexfYxYAbG3q8A4zgLMVU2tt56Fn5+UUhIN+0x4C2uuAs
CezUdNWndahHxzBc0Slt/Fpc1Qm97tjNW4rfOK7PtyOVciLCk9LUCEbbzvRfLHRRv5fpd/y8pxG2
X5LXCIpC4kS9eDYKPdqNFqXMrgbJL4IuIt5jvIOqvBDKNLkpTszPxN0dkwJnOo+rAaqKwz5lJnFf
aHYjzCgg31H85HHxzCUN15lvR6NDcGUvKuoLQGSsjRBSnvsoPr+/f2kmp380aKlCdUS6xU0C+Pv2
BcGOl7D0yB4LkF5JfooALYo+BYgGs84x/TqNJ+uq6DX45aF7TkPo+C5O4r+t7v9RPClV5bxzO8Bd
Fa8xMQZgceV2hn90pU6wjd/RKUWObQuXArVznbS9b69SWhESsTb61yhaY/KzIugWtUMudQGY/e7T
+Ul2bh3zzpGhhnnX9AK7Yn4xURlLiIaE+fBIvkMoFIOvhhM1oEe2qJ/zHCgxGcXusd2Dr7Z4TOjH
/N+RbOV27WdrOZmh7OrxyeiNi2bXKcC/POrz1rIbYbbR4EIn9rgBQWgbv/+rkD+UMMUPTAxRsXLG
B/xwqL4bwEz634nCCySC2hTtW0Gp7p3tF7fHgrzQckP3CXvVmZds7AOGMY7je8h4HolgGEGzlDTd
RjqGMRM2OW/xYbm4UstfObPNLC0FVFnQFCwPNL/YboCdJKnRB4qwDs9ZnvaRRcAyU5G/bVlwKKuU
NbILlQ8hkGcwvC8i2aWwjRmK8UKqzo+Q4GZRPTFmJE+20nPq5Q1qC3LOxel6+JSxn6zjXmaDonU+
ZAe8/h3CLOxgGm4V4xM2McM7CiVqHdlOrYryj8nFQ2AW5e8JD05RUivTXwg3QYfb15rHJ/tNZAZ+
xACCgtrAX/cWznCdqzMv0PWhUl2sZkw4u79V8fDWi4u5/nW7tA5BM9Ew6Q8UxVLQlMy67LzftvDG
gTCbhcZ4CFDKuHek7/AqRD7d2CV4fQOGXyYF647G/vxVZb+f7If4RF7/kn6tVx+WVLyDyLTq4Tjl
WOWvS8vHry2y8z+mJD4XKl1vzxeBnI9sbE/ZOBEKRCSFbRi5dv20vkoJgCwY28Nc3BdyMIhd4J/3
AxeMWd6gzH96ZxrVai2QU4yHLn7MRVwF+YPF3uQFe7S20bKAvrnRlTwj8qtxDZy61xrZau+UAA4w
CUm4g9a67qfsW3Hkl3aAUpiKt3YGWP13Yt1j7BuMNHNoQaYFsYKa1gvJA275fd6MK0xcMNYjLK6z
rdvXFQse7z99iFJgbxLpStVDoLMxcBh1D3lD+vACdxAt3zuUZniWyZsFgkK+ifwGopEjsSzXZXr5
ivIPtA7kccPc139NWPHlqUOh6RcTsVL4QQm31VrP9c7UBEBElnNfMpkNTy0dEw2FRc3UdUzwZEzV
/uPmCoRdU4g1SK991IUU0WgkOjQc57tYofPEuzEN8yDqXElwvrSfaf9VnPu5XNwcwRhFS1TN40t9
X9eKZ1SgGwH0ReWvBp7OxoMhfFZuj1NT7BEcxSdJfzfiSKn7DPC3ilGGfIOdaCMs3ZEh8Hg4hSUm
2WYt11AbKvDtumYvm1/Q94giwXXC5XBTcxWlDFjmufd0/gaMoRWLfSsSUCK0Nr3b+GwmRBHLX8LU
g6HpOIpVK+17YUrqQIARuPtlMF5PXwgNAwKtledeZPERMG8B9N/uUw3ToL63OiRPmz+o3pASaW3Z
c+SFWHTvPDJJftGOsL5iUYxonkZM/gAM2nMUSfxhlYi3I+TZEN+NY+OmLExFkz32rm1sVyykOEYb
eWhM5zSWQIXQIfuUNvJQYLnSLrmAwlUDgtKuf5zatU2DIyfHW6xu9883Xe5ziVvac1wcTiAKiDIk
Lqb/RFz72N7LmNqHHBelQHE833LWXZOtGmcnHsyvjsyjV1g2rmBUJ+BMooJPT5/Cm6krAyOJDTzp
uQj2fViW3nn7igChB0n53MsN76dsIH4mvTr7hOQmz44Mv+uJwmr6l1i/BsCpY/kvul2zaRSExwMf
Ne0XKHd+UKUrIo208AueC3Z+iung91vTRWYPJGidzzafIGTCo3dAEy+mtxsUKPau+iZ39J6dbkQ5
/BzmV4eajq2ZhvbHX7Ghjk0w4/rzGDA74ul4WmDnl9KL52/yP055JvfdgmlBD3kQJHwZVCVw0o42
RyWK6Kz97SxrtJBpFZK1yLlQ8CHi53JsUzQ7DH2+Aqf4barbGgo3Yz6N738VPT36FN6fKCuKnno5
fI4xTemF4U0X3dpRLLdxCt/TQIa34MRyUS/ZIXb6zsRDb+PBtBfWZjKFkM1N8Jq9Uq19xLlSDZJC
lvSjPo3ATi0xjye30B0NVhAF2/0HvtMu7zWBj+qG3K0Zl5o7sKp41SnuXwgq/9lw0BaxdaCDbzBQ
0HC1+fZpAplQ6snAWB35RmN3pntjA4FnceBLrXEQ3JVvB3XY3Rw0q5A2w3S6XXl8h+NzOOsE63K9
dW0En25dV+/9ZMgsAgXibWCOmp2WWYsiuIgQ3oxP7MZTg6GkSBiCtwyuu2RsMAIJzUQPkPlh4eO5
ggWw8E4nqj6pP9/Wd7X0zcKb52IZ38D8ABuqtuHsmoe3CuOTUyL5UX7rZP80ttfjkMKeOj5KNvXs
8rFzLm5mi9t+u6kU6ydgOJxLf7Kmd91pXEUSn5WcEX4aQUJU8MEWw80PjWaKX7gu/U4J8GNAj1PR
mF0ZkR9D1Seu6XH1Z9auKIWBhxiXRBR+a++mAPhs9u5wTIZ+gNQZWfXPygx+nLWDYbCUldszD9C6
02MCcwVIMdfy37bJcmlz2LOiaOP+UO60q8kCeTv9V2IYRukAtSkFIwEUeCcfT6nvcPNSA8uMM5uS
e/dEVFotvUPLmKSZpAinkz7k9kfhWphVvJJUQUyB2riC7zjslO/X9uJIU548ixWAL4C3l25fTPwA
sfjoYDCpNaCArhRubsGdDB/5VSbrYHShRzVNX2W8FQSgOr8GvXoRHgOiPNckwhgw0HDPGf0C2e+e
ZEV0e1Cs5dXj3LS8LIVKv2Zgq21HwM9y0S9I2Xfchp9MyViw3jpPiN6CpA8y60xX34SxW1ntOshH
vjSs8/mtwfF4JP/HEE8FlvpHM817Z5yAltElIbtimIyJMxvlUUsakezfOjt4g/aQ46U4tT2uDWTl
G3an1WFC+RIht9+90wTFLdBlzNT1ATAuH/5cC1Ql1xEWBSnl7nkBjxwOdRi5Is2IbIHBjwv9ErwB
4hFnJ14giH2nluduwACww39xZDjw6fUfQk8IhVT9x7xaKNMXYz9GjkQ0l9PK6JG+NSR8/r6f3pzy
TGmCkX67/guZveA2MURbsP8YBUpQSo230+SZF8ngokYBVEVMfsWwLIsVqtr1r9+9pR3BajR5TZcm
F9RBrTRMT+v0hphcrFFUd5H48FThfCyxRtj3pf1gJLMVUZnXZdRB/0IlwjeU1IMtdek0CYOpCMpE
etMn3YvYZ0kuvkGXVbWzBdd7w8Kxpm2JsTUrHmvNcvOP2Eq/KkgzxHqRx2m6rhS/RAI3CMsJIFZG
vUz4/GO0il0z42p0VvssvH09l6T1UkPexNkz7fIpC7FEftnXwu0qM9JrHGy308tjN6SbEGUntX0K
n9hdQEmA8F9DHYd1xHIOARPfrkGIUU3bIhEBjkw0S30fe7cRVgm9aRcXR6b2a25NoyZQGBZMEN0e
gT/rxd8jKle7Dt2CUzLPqGdapkGT3n9iqXK5dZrDAOJ4uJ1xncfyEsvijqTYhGQOoiuRr1kDPZ5a
lr62VJUEdl30rVs6iodznY3JS+gPOGvNoJlZwdWJFFMpwH9PGC1SbzLDCjl+W6+1Zp5WGYVEpTOp
K8DeAnyqPMxQOwTNJvanRvgGjLOsuFilMiPPEy0byhiTJFTtLs1aq7JdKQuziTNAtqAZ0B1LJ6WH
2GxMujp4d4LaliqnFbDW0CzGDU7qCq7Xb5sNrYGMG8lESf8cPog3foHK2S1jigRAjKzZ7xgOccAz
7dlLMQH9fgqDoPVHH6s9maic9wn7LaZnum7fXMq+dKWHLY/bmAr1VBmV+RDjxkuImoxbgLoKp4YL
fY+F2qjLf1/dk1rg9jI2wgLImthxjwKYBBCwjnzDw0dhE9yRP15C2VP6R4S0ttEpAVJ1hcHDSe+Y
txtpaapy0vUe48dHTZugsNo6EIpYxPivE9P7Q8q5zjTtU8XSdL3BSciD0TvISDcSumqWIF9dreUo
cqgPSnMifESoVRdT0g6jjhE2/IAiea8gcHSCVFGyiHH+KTVryIECVYfUMDi0sTmrmB+jSZVNr+jL
3qi4+vNwISgYWKVzMdtomG3qDGoanvrJVsKhV9jX/jem/Hz6g344ZTaRFYwMBDmFcO/PDsnCbr1l
Eoq1qCGU9Y+Aii28BNaFlq77wV5vWtWP6MDRRMFw/Auo6TPHvXJw5jaNgXgcvBCgAfMt36kG1tsN
sHmHhCMOsQkNBMpxK60ESY2IxNvhnOMMg0qgAL8ftRi00K52mQXkHNBBQz/c9G0Hwu0uTOsYZTh7
b5Fz6OMhFTQSpwSOvx6S2vslH5rwx8X8iTAIH1XgvJahKM5lQnwsrjf8ScmpAznRO4v0HW4HONnm
SdeyYUnKuRoM2sd8FVo8tbMS7nkOQJDKNzEFnILoE+v+j6rYfYezpD5vvoZ4vfPrzbEFsAvJ3LaL
10n9/a5Ap8bZmoaHdFtdabZM/KT0XAF6lloee2z0anT3Tn10frG7NOXALCDu94rM5RQQe47LfZqk
3hqoxBM4g/6SnHy3VeMftKSjGDQFaYwiqQa3VJKOLL7qqdMIU6Kp/exx5G9VzJ2edsyCzgst2onH
e6g2lk22RwP/hiMM/6pQAL77sd7WsLj267XNTGszhgYT1JTh8alVuMXBTednU7m2l4BaVvbXckMh
g77r+Jufx4Nkkny/zU3IjM1JQALNGhtRJCVnwm3K8z2VBcsqOZaF4tcMSih0BhPXfho9erVlkviS
ahl3/sKQAKSozHbf/N97PPy2V6HO4bEb1TdCzRo6INPaviCII+p15N20gqePhYLtHXaoCT+4u6TG
3+wSCt8asQTZgHnieCigJva6jnkqScRC1Byg5jLqEcwDfQZ8wpJ3oOuoisY2NT10rTFGfQNC9ToU
GCoM7QU80B7aK/ErC1jOGGuQhseMMtq12aZ5xfhtZ1TxUR7Km97xeIbXNSQhirxGtPkahcLdThRH
dmxGXxdMzeQhUK3k01VXsE0OA0d7zwUMhf97yAQy0Ar+X8c0wvC+BOcVGKwfzkj+E/cpxULBwPCs
zhW5G7OKwgprCjutjtyAy3SQgPMzBdDfat2cp3JaDdy49zUBqgtePAC5vrKmWNIGffa5ate0/Znp
cs8rwkrqw37wBoFAd9F/DtJL5R6N6fECiDIrzSXK49tZB6vBmF2rOxv1NR6A5E+WuYFm5rUv+aI6
z+jDtL77yubQ4y0yHdEw2Uxk9q8kTkBd5qcilaC9kbwyI49wXDy9Qa6Gh8a+BJ0+sQpWAAMV618q
a+nP2QRDUy9quo626T/6a1suSzY2Q/TL9Bact8Y9BqW0m515C6Ek6Vl5gce1Hzyd4eH+0rKL+2g8
7ABAin8wfXoUePDMkqAl7pJL0gVwp8NRBxAYuDufuugu9WdacXuodkKSpH7wMR0XVJ9J3lRsAy9h
TVdWBvMnyDyADEg9BYWwQlQXyBgXVvlsx11r+QQxGjup3+vKiqtHDa36+aUoihROmSv4hIt4R0dR
7aAjJNcvVN4j9X1MgWtyW4iMT70smU74jCN50suaDYZOEVIpfhqyqb/iThJNRXxQ4BoctZqA6sCN
LqtdqdY1uc3zIxfT62W34l9NmdT+TLpjT0I2FEQz9FVmGjN6wFUSj0pRYXTa5L+/mIpvj0LeISXD
2WhfSa29ziAd1MGOPugzihaFRu4gXyhJ7mDDVjeT9sAQcgCfREg1KMfytDbdr58fkGkSLgRRF/H2
ALXQjTdnvcvdpe18VOMUs/sraRJ8ZDWmPejIKYJKWR63nCGH5eyuBN1z4cLzxItwMuIOR7Uv1k4u
lsJHxtVrGKkGGKtgA3V0zrT2ryhadsvg0uFGrkqxG52/ad6FLflC1MmpYToxKX68O0Dw+XoDWSGR
0/AlvZIq4m0QXifOZq4Sh1ods+78EbuHjypgoIsHs609awrBwab/3gfZkHu+xoDchA1pNhq+xYdg
fe4s8YFFC/mOiL9V1IUQQJ5Js9EpXaBfxmvsSFA7BydJD5cVxV8MgmYNO0SQ8FXkA+2yWFWrfktn
tH3y/sPK2tCvI56k5Ik/ZEVhF0u0owho/ciFqIgVUZEjVEdJ6Z9QWiB/e4EIOwJHonl6tJDAOwU9
k5DV7llxIyjmYuuFDJdIvU7dEddhx6xEiOCqHgVvvTsLD7JGop6o6R0pX6wVKiysTgfkHe4Jlujj
8crzCxTP8EU1Sv0mmIamTLEdofUJEtUSapDxc1VZ26kD+5QuJ8av5k6rLpQJjOtb3vB+Gvgmd0BR
Lbf76HCUPUoitt8ZaiQ5IyR6md1TF/r7TKdBxqLYe4jLWwVgNkk1uw1SLTB8gkYbgZHryEsb5+ds
N0+VVx0WWslyMnIT7M2qN7Ry7LZcAO5pR6h4wSJx2q9XaoKGEvJ4JmVLK9oVXySzDQFIWksx0V4I
G+2xEOg+sfzguyPDy5csX4lazWaANDSScEaZ3Oo6bjZ6CqgvqrySSxJdyjWUycBiT3UF6ylJtQoM
sMOZ+1ATx/M1mfVf/DFaH5C2mEIIw4uHmcY1MWrYoja5RqzbPEAzSEeMnQ9rw8b8jb0+BRTJu6vH
BaVhcwn5LaXA23HiTX4voykBKf+Zq9cM/dZUY9sYXteTWN78lW8+IbgqL0g+vF8C1d/gwqh56h0y
JPJHZPnZG2ewN8pgkRCGgcSJe2q0tbeT38UMfuA07hD8HNZarVvfQ+bBqkDyGvDDX1S17/9u1+nO
DRMnZ69tC6EBs6imb0P25lePzNiXakAp8WTQRI4SdB/g42Y3NuSPuHB0qfBrIodZGyEkl3wnrkIb
EDHEfAo9Irc1P9+mbBSNtDwpb77LyKXB+cLfvrQuv7E5qFf+bf1Gf8+D3DoP+6hd42Z12umhk+72
ynaDkis2KbQGA5dtTyJA2ctqhGEwWVQxdosAx38byBKY03t+TWnpf14bP2Pohgb4cjVbcxrIBCos
X37Zq0k13qoZrDJ0OsTUegH16O9i6U2kq39hAodNtQIM5+ZUZar5+0F791CzcRIR3/VW39v0+8k3
dr/cFNpvNUSbQBg7GTepLg8i7xNjBtuj2/Pc86yup7ZsuS74yueUVXtN9aj222mCRWVcePdelQBJ
fV1fjJXcBuSTzQ8xZ8cJ1SEGcgBGgvwgRmCeJRyVuRBowAtBF2q/BraV2A4b4UEtzOVZZ0tX6SjK
kP5VyhGAfZXkAtdkRawWRooNZpnrSUz+dfESdvCDSK/niC0iEfP+3f1T/RJ9n3XJstUSsQM1Raga
Ownx+wBFhyfOdw5kkV74AM/6N7oS1zl8n+f/9uQtKilR9ob8Aekef+E61wKuHXFecKBxOkkR/bU0
mQsmTnJ17lNcKr9s3JKXOG8huGollJVrZUt5MkxCRcT/XaizTKoEWxwCqvvCmcEG2mcCivYO1Mbe
c1b1hYk195MUP+b2RWgmf9EwM2P/JcB3/Z6I0bpAi6C8/LmJjpRErfiutao6RpP6AOzJPS56ae1/
A/zJiPm06oT3sRhjSbVwoyYzTsSTwYHX+iDTIp+p1p2DMpEYJkymRVIBbCu0q5pMEWmzzw/ohjOk
08k0nXnc9eT+GGcSFXJRLo3IERcHqNzlqI+E5dtHVrPX/F/GFFgPqQoQRBhiuIwlVlbQaNI23FjS
MjWrYCOo4NyeOStFApdaFpAPds+DOYwdzGkjVanQhdw7yDPNrEm54kH7hK/C2xP8Vq5a/yIqzPyu
SYI21/uIEWR9+yUTzq/CgLLJNwsZh7C5cLaTxIHxdFo5Xx4pQtarbsxgmGSJ3jtStvk36lwiVPAZ
IRvRMHgaXPfk7EBhmRA5fkSu+kRHkUj1vHsoIKgPeI3THjbh+KYeZQQDBJeLHPtnRRkur7YVsu1A
oBnY0lDebyS8w6UFK2KaTRcwG7ePlOn7LWXluLZFWlXIlNa8yo8x7NegyrDYCJDCw2iBxVWql0Rl
HNivy1+g6EchFsvvGwlbpaKKZ0VKQyKwc4rFyuX69Fcvqyiv9waAk/WVbvp9ntw/gZs53lhP4/Cy
0cQ7xk8vDQ7VfvTExfM3jDqr1RQfgKOXwAjAMSiFStoYgpP+A/E7cWQDNifRvbaAN4haQMNobsmV
W7CfssDcvXoCK0pOxR3sO4xpcy7gZLk1r2ISJXCW+kB0ZW5fGohKi0YSi0GCeX44rI1TW+dMi9Gz
AZeiNPP/2VPWJtCqWgug6cqayVwK39mXxJgjEULdztpOelqfdFBGhA9EHijCFbXPP52wr03yPU2v
GVQcw3k5IH7tC6l6YkPbvXv8DlfGXYIjDbj7Wpjr7oQUOhMPn5soGTfN4nes2WT7weXJNfGKrOtC
AhFj8zWqao1cf6J+n7H+NBVmIC1zX8AUmJl8YUYoZMfvSYimTGyRR4y2GpTCvydYQzuJXPIXA9OL
Bz2dqZmVwrTGQmywAZe6Qs9PV4uXNzZFzD02n2WgnNSPJUWF7+0DIyMAdB5NjdquVEoUqBtg7Jad
2kZynCVstsdkEMSpFuJzM8nWXqmqsjAEiKaVzSDsyxtKNeQ+IJUlz1NamO+UYQU4XVUkYQ0wLC2v
3bMIF1wE93rYQGQiNc5S3O699gN+MSO7pw1vW9TN5Jnmb6ERAZlbf8lVfm04hSBiawBAOBHKUpwQ
6Uz/P114flK7GHRn8Zv/7sz+oiNElC6fBUCtW1zOYImy77ibKfv1ZU8yZJNlTTCKtgzWIM69aCn2
AKGl+8Tm26RIgcTyYqaiBgtKRRKh5Y7YIGQQIKRydEg4LL1VXVw3q1NsKX6OmHskR+mITnOQ9pf0
SeC4CtSIQG0aTlKcg8I1TDrhiqLimLIOU2sGHK5RKeNKO/B7JdjHu63PzkV06dp0gFc51w7RHDXA
u8wipNlEQGYQPZFOlsFYqfo6H7hUCm9nLQ6I5ubo2xwPjKRU2BPu5aereS8ulTD+cMWI3+uerwiA
Ov8clA9yP+9JZ4CzQVIiFcUh2R2ZFg3HhO0gd7r71Xw6Ftx5ExbTNQ/BTcMRuC+0aGeDWnVd80+M
T7MKzjayJP+Qd6R1NTivbq6EOE/aCkrq+3dXsBEu0uc8plyZRPe6OhjC/YrLG9/4gIeZId+Wyg2z
DjL9mNYIa5EG3YifloWYP+IgmcbJa+obX2HqKiEM4TfawCpPj7o133AiMz7wCqpNGSLylq1FCfq5
bwqWdNp+PZ2Z9TJDmk/3VnMUqZLJQ9LKES0HAXLT543MsI+7lIf1aQwNzFuzOMR5mfXRgQesbCkr
p6ZB0CPqE7DtpOjQHu5CXHNnMCVUSMPKbiGecr3eNCz1qcEaVF2VmnMIrJ38xqrdptVWVpnbKTVJ
SwhZMyyNtMZeHncukqwHmZW71B6pVB58n9maF2VmmPLTh6cDlwlPqeAvlVUirPOs/SOi0MmIme9i
Mmv9/ybubjeV0akxbT8LEO74xWgDfvQZJVD395xykKxo4lDXAxM48ADEPe9kqOHxnkD0u03i8QN/
EoBj+wdaXhtKZ5aaNzs68ASN3iBZQ1WyRtiirJyIoKIiCQdoYY97zLSRGQ5umCoGTXfVzbUbQUPO
uubxpubrj9yXjauaM57X0Or6/oSLVXWqlwyFHHGkM7onvqCuX/joCc+0Rn2oQ8qTrlIFJ3G+FstX
CxgV3qlbh/dxcW39DiC8BWwaWZhFKwrzCB878U9QEAcIKpNhFxew7LMFKNPNM7rJ9hRltq+kEeXl
X89r65tLmpgJm4ZEfF/Lc4zlVbA3WO4v+SsKkrQAVithoZBw63OM/apPhblJvrCGNGUz1fsoV5ig
Wi0tfcQQUeVkU86Im86Xsu08akeOSkGy1YwSFbVjsVhGheuXW9aJJo0WKoCpnBDRpavTQWZRi4i3
Tgu4QQ7g6SqUGKI0cjM5HMrEC/SDPb+vC+X2l1suHlOxb1bMNCb0EX7cNrX4xFeF4hwbwlYXc/Xw
/coJUB3HBv8+KSCgtJW6mm5ufSsrxNitox/2HuSXRjhsngTQntB6muf/hQW/xdjbL6/hr/EYXGQO
Hg3BB0uzLZL0ukxPRJYrYdTOTXylAuowZlv1wY/5uNcuCBzrhs8gNf/zJLtUsM6h51zwTxOuAzBi
ELNqF2akkT/N4if5+hFQ/D+5FEazPbcizJljUiWezcevKfKfhCElIU3e5pMcMQiGBUaYykJpfpne
sAkjo+jF1UeNaBrU0k7+vuW5pEwvnjkzafpPi409YhxenVnOLeVcrzCmM2QGBctQ2V9MKuQvA8Yb
6ZCjEpVcSxY+kQDwa58LVpxZpuqYjAJGM3M4pdgWn0Mj4+PBP8SYUGY1/0sEQfm/We6FkbmC/zPN
EjKfgLyfUDgYrHAIgH9EgYrh63weCAFbugX3R0HF374pTD/n5adICHk40jxVgCc3yHtz028AfH+3
fRlQIOO9YLrj2wtIbsq5igwdabdKZ5ufDckZ2H46gZ7sLR48FgQ/t3ZYbewGXKdupdcn2soCe77m
645+YftRfzNAUFcvyxaN/NQqxF6sT8QJvqOv+34q7wJ6mtr9Vu0t9tgg0gUn/knNHNoyEwZSgUa9
zZlqPvlqBZWK6E/CxjwW5/RpW5GIlpSygyCYweufxy/5yDBq9yRFdU3kiSSpMNGEzTyUhos1xp/K
EIODY78ovIKqnuhuS+PFPuw/r1LIAUmb8yO0NKyEEhp993VO5zRtcv5dAcfTVkNOh09NNNoINEe2
RIqihr7k08UT+U8iwBnyr/y3qL6y73/5XHB7iv4Oaecl8vdjRK72eSTVOP89Zatk0LBE2ZTVBL5w
7t8/TLTT+3WQ7SVv7LjWfsvcbP2UovPDy7sxc4hHwp2Y+1QCxWXg5gayf7cOWiI3t7yLxerX3b8e
Lat5WkdQVIBA6BLcfUgSPdHJloU9amkg3WQ5erzjDSdVs5hrMw4UmibB7F3yWD4dp/06OxHWb6sL
0f5WjVOfs5LV2BzZy30uwat4IUoLTIe44VkRDAtHoQjcrNM+/Pf+A5W5f8tbwpwUtb9i4mEv0kf4
MoB15i0OPxUs5hl+zF/23lyzW2zIUHKpP6o2qn3BmVuCzCr3eZz1hmoNfyZKjkLUnmSCjf1d9bw7
sJwwkUDboo1phAT7sfnWHInp3abIJaG3spXY+XoijXvS7JnU4PSpHRb1pnoqvT6aYGhgtmCCt0kb
hkPM/yxa5C85h9o1H/j3NIuXFtyzqwcCuZRwK6T/jBkiQUY+VNyDkfJp2iXBIbTSyg7LWpHdgRKj
UM/6O5L8R6i08ITxCtwupYHC/dfgy5z20f4KktgzUwtg9uLAiMe702vh2g2Xo9WS9tVYFYx7Tt6j
jiI7R50cvyWkV49rwAtEXGNDxFYvL3JNFy0lOxV7OPjdYtgpSNW8wdhGDI3N9M87qEBMMkrM4tdE
hkji0dJyXH3Ha7G+VDllZbuXG/cK3GnGdi17uUWqPYVR/z9N7+Wxz6QOyOstv/FspyTvXytTArPJ
mXDpgZLakTNbBbeJF2Fuko0kaWnpFuMezHICz3od83fNFwbaMkrnuFEYPskyuEbom3ulfA2VUHlU
RWGSWnY+GSvmTs5/n9g/CWRunqJoUJ1+ysZqO4qQqUiUFwfiNKNtAj2lvp2Gt822+gpj2IJTl+Zu
KDoe+uHV+jmmoOdiXgA7YCZSuA1Cj7oyXJLsnRSp9m46+fZVVb1EPqiYaavgYMHczWCYdjvHBgeU
iZxLaRGjeS3rYQVYlJQcUxrax1h1X6QND4LqjmqsP8pmdno8iYD644iNn/h383tFF8IuBv/oBDxW
rH9N4bXHJroTdLdLaJz5pBdm6gs2yjXc0L/NpPaZ5skRlyFD2AVmjVxzPN3+yICY9qM8iNKOa7pj
PC6JPsftHZs3sy48AGUrQv0Jd1RtZA+doh2ZAoj7DlKeRxdNmTGlDpSglORcLqVJxE1hoLYsWtUn
lsAwEG9az+qSY8BFifD8uCCCdE3/W09DyS0qxTRrDhR1LagQnBU7K4Rhm8cEnCdDJ3ckG9V9FUWo
PDgcd3nvZP/AWZLZENPe5oR2D9hA+oBo4z5QXp0AlesKe1SHlWPNqwP9is+5G4BPGb7g6D2R+k4t
7FZrcv6nlQmYfaKFkqnMcHFhXDPMlzrr1pX3REEurf1EE3B5/9voJhjouD22ECg1TJIaeizMztpS
3NYaIzQ6EQiV2n90TvpynK+EN5uYvlsPrTN7e+tN6MiXXjo7EJ16uLJVmnXJXu7E4S6jSqOt/OA5
TG/0pqs29oMNvW83JDaIlcCa/Gon1RjCeoiTH0lSO8vhAGuxO/U2/iJeHjCDPWc4VlgjNkJUBWdG
do/4qMZAodR8bJjZ1Nb+35fKSQFEtBDYtPdmWiCdbc8Txqa7VCiq6Eolv7yigmFjyeaehOHf2K2c
HEsIr6/Vn3N3rGhEveXjJmVVuj3/MtJeAlWbmwRtXw0E3MFq6cNr3lGnO0TUFffzt1L6QLuaCG0O
cti1qStZcISuWHqvPfGOYdYN5e+9V2E7E9Qs81bZmQbojKXFZmB2ocAX3UhBycllyPAsH6ccS/Re
LI5rHD9zjBCt1ZcyrtOeckK+WuvDCdvOulmQ+rhx3W2YI0EnffqtKgkwB6Vxrx+l9SqDtRsvz5U7
OZYcfq63fyrxdHgoWnBJyh/9KScnBoZi0gLQTLhQb+S9/pt/fpq6i6gcnvxa1Gew5pKZrj1V2CuK
dPwzeq4ZQo1iVfcc/OpckjWIBht8r/IpL37ldpD3ScjHf9hATD8zAwdhna0Shh7vLF2Ndt+WHANY
d0eZUHRLn5aorbvCAi9kKIoMXrtFitQWJpOjpH0qeCX3mtbfAeiHpMA41zGjyvbf9kcwyoKuUsT8
sotQN6gwXeHNpvMONY9+XbuoK++us7LHAIkTpwOm47S3Of2ZB5zxOytlqKHaGSHI6AXiTJf2bbJW
tYfkoi68CHI85mVotYDnwuxVNpGxzvoGR1FLEkJLEjUgEcFt98yB6B02oLNxwe/XEGLLJ3QrZJ3g
+UgsraaN5uCBOj72b4ECmem2nKAtA+CITUvJZXBfZUTs78/DawsexXJnZF58hyBXEgDtEH0NDaVN
mKkHzlX6t/teZrlUjCmen4KqNaVtXvYs5YfikTZlrUBrQTNrNZ7BKpQD+nUstuj8DoAt/G9SNaPd
OOS2scksC2O4GV3TiJlul+LHFZCmByrVZGI6oDsccE+nusz9/7VAeWDbYqOpgHJNyk/XK5wSAnRl
6+XHb9hroN2WkNmSDIfroWb7wpuEey+j8aoMzIwNx3FL2M2Tr+N1TqdGleWAk2uHEv57sJi1QKF1
YjfP5Ghw9Q3RzitnbukNFgOwxHghWfxnFj1r/uwMQJ/RbJZgwenbXKDkgSKWK7OI6bJ8Nfqi0lNx
PC0+2vgZTrVaqpFakM+ArSHfFrXYfWCabCyW3pJ+DKKbENFGCC6/8hrXDeLaSQ4SsZNveLkllphG
gk5dlFGaLXU2uXK0glViebwhmCMcLuM7AvEeDsqqFvI5LjeEaSCCa8dzP8xX/8WzhR7+6PyJ/Ji4
knU4O09YOGeWIpudqget+/Idc0A7wJd+o54da9kPUp3a0PechQhlDUXSvYkiKz3LlUIXvBQcIaV2
U+9V1EKu7NQsmz0EmrFNmGJGSpRTTA/M3uFy/QZog170QiqR869bykeC9n42crCKoaBx/ccofBDj
PZbTyi5C8a+KM6IMt+LiJcygUwOJx0XmNNnOmwvfZN+hTy5K0JvaTJrp5WLWy+K8y7xgaR6K4oBn
G48PbCOOHThGrd8OrOkXftgjDf4/5K5NIra8BJ3vSKhHf2q44utd5j4Lu8s3zsCSFiL3D3mseyFc
5fmxEkfiODngCqLtUJLG7dPoDQqV7+jsLCTOVWEQm/gpypvymBDzydR9OPQaAy8xM/Lr6X1Quqzs
QGnCyd9WFvXYMmoTE0/tzLC6KmjeElfAVCyAG1CjRIYRnEbUxmbTbLBS6jiGIFhfa+fl+Ma7kbDi
+gPPzFEmHDt8Xije5LwoMGiJgfWqMQVJOI5+Hfcc8hGeAW5YXgynIaGM2qcJZ4C0XC/5t6espMcl
+ExCgH164rwtj4sx/llTvwKF9vmnJ+GQAkz5hFtkoiFg2ejKMXgHl8lW+nwFeDDspWICKKyLWFuv
hjLTNcZM4MOo145CrYrU29wOSyfubfyXBF4R7QBYrCP+1Hw5zb37iBf8bQ9Jc02Fcwff45fJUeD9
QWrZMx7oo1FQQ+rTQNDyaGUXd+nq1Daw6+FC62aFMlkdt4zaUhSKbC06rpsl2KvW6W5fyqzYvI1T
0/nOoS6mnVbpB/T+r9q0MIlhlPfcG/YtpVO6nvGCaUTA5rVxZbyEfA4thPFbmyEz75Dr5H7ZFOzr
UCFcPHM5BBsran3igppF0eLCXcUxP0n/3Is+jCAXkUyd9W6/Hc1uzn3vk4xO8qnjK+7vZ/dYdVnA
0bXqzOmQMyO/AnWmlMN8jusr43nZKM9ZSR7LzNs5p0sIo1DYO3xw6Xjzkc+m/MNCBYp4BNEQCB8f
qWuXks4rDFrHS7r8V58+xldOx7FZ0w5cROy8Kkmi6OnbUUsXp+IHxvyk9dv567VjC3on/jvdmVt2
TjNFagWYZHnDYWBdsiMl5IUpoeKbLGDlaAOthAPCVd/dYAsmI2uEP+sF6Uz1n+3kpoAZJHYgxiFL
RxQeKYEOtes/CeXkYz14432JKXHLVuagKYe/Hea7S4HMIU3OX7CD9XZu1NUWuWc5xLLOms9ZvOxx
LocBTXs1t2lfm6Qg8uj9melvGrQHMREaGOTI7vesgTmQcQa7fqSKdmG57oDIhgYwWZhEFLrZjj3T
bNjyaU6WEzLam26eEIWSFJSYBBAiJRPGmO7AhN++l68qPpks05hR0AI8YHcBB9qxfT2ja2CKSqaB
bZFQIhOTguAuj7QA8clAzvN0qu6aHA0X6WxNx3vsw1puvQ9ls6/9SmvUHk/SmDrUFkezxV3RJBpf
5A4D122lTIcb9p+5dlp0jDhTHHbA9A0v+DKo4vnXerL59IdIuTSb6KcNVrWUXEYtrauVT09mYQkh
Qux7aR4RFQ9hZtxykGX6XqydG5/5jPIHThHexltjFv2fpDygZ2DEp8LGKsSjpsfYxDrWSlO9svYr
QE7CvJAKW4XCs9oQujIonv1iueWVpCR3hQ9wboeC2AE+3WvxL6lCHBVSTR/F/r6XeNARkJAib1gi
vtMmk0GtFkLFsXMxXWFg3/olLC0hWuRij04R+9H9DOIjs5CDEi8gNyrwzlErJZmUwi6vmRz4BamS
JnhMsSYCTbs+M3LXFaLvJSjqLjzI/XSbJhGSrLJNylXwsanVZGb5H+pm5FLzB/7q5I56Pv9ecSB0
QRSVMhrRz+NoHoVWopSwrRMq0PGajWysuu3+NUjqU8jPgq1bsr5c++ay+0ti0cs6W2RsvfhDg1fs
3M7fDn9qTRT3Bm5suE+wOghVx1oOwZ8JR3+kU2jUK7jZbnjiqb4wwVu+EdOvtc8717z//vIt86oG
wZcD/qriUgzQnm1aNKRuqvpGPj7ZQx8Ww/ScbHQCnJHuMf5zg6P/rWQpZ3Bu57OP4w62Xj7b0m0Z
JJqaszyud0OMYnNIZi4g1EH17Sf4UgjtW+kk2j0HhyCuU9QjC6wM3TwVoJBAF7Jj33PmGj2x+qIS
MvTbtcf3SE4WKep1yfEyfDeyiUuqyiTPN1b2evAvK/6YlM4yNkDYHWy4XuZ4xnlkZ9Ed+Kvjs6+e
ER0YpMROkOxvyD7wV7K7i6JAfJXfTRk1AMsuw2zoJkxZkY4UjnlDIiGmK2MJQNnjUgzZwu5j3qnV
BaW3ITCgkTbrOqgtd7qwKwGsq1zFffWCG9ymlkkSVny6L1mDarHlwGJfBz91dB7K6z7IjdQB1mt1
PJmfyffN3Z11Bqaiq1CEadqSy+5hMRY6mlk7c3FsbeQu149ILTzbL5qX7VfyY5ebzuIsdEMvc3ai
Og9tUXjmKYpQmjSvr7qDbfwVQf6ekLIXCKBAQFlBkzzsJD2UNNIQYh/sEtSjZUkwMGykXhRSFYRH
qcR6aoT4ofQOyTnBtRAsp3D04t+qYMeVpok4ACZezxYTCLUvBslw8jvKO+j2bQZ+yEqzgqzhsTpr
bC9EuR8f5eZDKUyeWtuYTvGcMI8Hqrs8sXyqIsuD424fM58vys8fNtfBqMXOkjNB2xgVRr0w+aFG
O4Z8XnCuJgWr0/LVr8f04zEciFSpeUfwrX4cq5JW+sAtmhhVoDou75NMMMDtKE3YQCfpZlr/R/9d
HjHrEEfkI5v99gV40hl5NoMPTrqKlqgGgd8y19e2OoLSH82e9Evcqexm9A012rGlk4XzT70QIBaW
cM8wXzZf3VPleeSCyPlYXUC8S9l8tCiEx0iMzFk6BFVBoTr3kpcc9H73Y9TUjl1Z+FVJkMt3ElXY
C/dunf9ls7qRhutmUSJ02uqChRO/r8M3blZpH80ofVri0ZwfZYerZ9PI1a6yX6mcjn4/mqBX8Is2
wXbA+H3J3PKwf07bv3k8GUhMSzyXzlmYYZJ09G+9tvKNMhvihdzBbox81fq+IxSRwmAzmQlLMb85
yaYm7hBfwLBZCWtnB9wQpp79OJxcaJTt7cpFrpzlthxSwCpkxARxDXDdsh+zTiCSrlQljA9/p9pN
MrWfN4hU0XInQh6L9qjv2x6X8gCBWOwZ920TfrLaRZX5osxLupEs0N71PiS4TZkkxnCDevG8Rvrx
j5FqciV7SdkRQOz0z6BU4Utjvv92LG6DIXgnRgJq8DQ9bnfEoh2hCqCGjGzdDFMLQS+X/8LnOJ6f
UoeiFYZaWkfXT3LUpf6DXHzu5UfMmNvbHI0B+AQDbgQJ3TFfpmxMcYYpEGqupAl1p30oLsQMEvbZ
mB0z21NSLfG7INlY3ADBBm8w+l+hq5Y0srNkBp/A1g2iIiU58FvcTiIMT85axI1KIgkmXeE2yhqL
T/n551HxpKLF8q5QE1O37UxxuxIM7BxkNIjXa9g+KmJ5mibhRkmjm/R/li5aObmm2a8usrB4EIjV
SLfEJbvxP3eIutlfFjXQGPtv4QHueFyhlaZlPhH6jnfv7IHC+6Cqc+6Ng46Rvy3O05CUxLpr3UOO
eL6f3jFxGGqJo3GCg6qMGNvCLSkmjWlmaZw71HZrqyMArCG2aoNopyoJpguf/1FBXPer2Sien7yq
V5NiCsqA1IVmy8lMGlZufIxLC6Q86+EBa9TAk8yWNr8HVOwE9oCkPqnAikanqZ2f67OhrIjGlLOU
2EgJUOpA7fJ5Ez6M0oTHLmpWizdWaV2URjhZ9yRBaLfcueMssi66PgXPlTrGy4Z/JjirRHQzLf6c
HmjNZ3TuWUX3lfb6oFqxfF5VSR299sANFe51/+mLWctNWvfv2ZiKuZeRw+clrZX6/wPy8+8fLSrQ
2CQj8PbMOR4JHMHkxSq9XTJBoD2tiR5Q9eIp4VChQzCp11VB/CTtnwFuprjLulaB7f+rx6XGQi2Y
NnpJD5pxl/7WgCnPMFYoGQ/VyEc7uPnXDINYMu2jLCy4fvTya0JRkdcXp3tPoCEKZVPUNVPykq4x
vPgCsdNE/NlK0aWlh6AsLUzRhVj1j6oXLcBgUbyp5V3VXXhpDQ5qFJQ4Ws91+FbRLSPIU6BIpLHX
XnkHDLyND33qD4QilvKgGmk+/tz2qeB0XAhAL0wIiok76yEntJRablwRuvFU6zZH1ZppCEZi9W4m
KEduUixobs8y9glcdfIH+rhzhmHjuSetFszl9Xpc9/OLoOAmsa7Sm+r0uy9zq0JVbMUKhm+r6Egq
nu26RxsJ64oUjqRMXJixwSVgAskvWpCMWK/oMShB5vpC6ZbrgflXTm+mdtc9dS0f2oegIlXImNBK
Juqgw9c/7czQScMMkP0cIiUr6B+RCAviCbxm/ucjfO870Gcopdyr5Emrf6xcbiYUI9YKA15n1Xyr
+lORBq2ZrduDH4RMLl7MZVwokqV1jfgTYIAOf9/C7iVKSl+49pKsRfV8vm5IEAYsXU0F3lEpP1sA
6ec+xy5LNwQrg+kjpblGZJawWLH3TrzMcESeU90HM3fXvdCYF+SfN+7bbbhXaSGn/QTBjjnfywHC
+U0N02zZn+7I9+BSNixZd56jtBMUnF5btelg5b5nZaulhLs5Iw3Y2GsxgExNwc5zEyClyxfWZFCH
Bf8FH1fSosjtESl8noyMgLvaRdLdrq4Tqe6ImfPHIXs5eoAmYScXofVM+cmVGqqMpmGKF25omKNI
gFoto1AiNvs/iP3QNe6AObZE3YfCw+2zRoV4TFT/6C6BiJ/r1C2fc4lTqbdzxPTwyalWRUPgND4Y
7PivtODt713PoAC9FHoMAxfC5sNUy0U+m1CMvCM0Ic6oBnO1Zj3w5uLrTipjNVL4muZQbufjfxGW
tOsb2gt62123XcIStgS4hMTYue/weyDm/WczQZaa28SDWvZQAx1KbhDtyqpdSw8RYqgDFFFC+qmb
2j9i8UFlFMqqhGOwUszfl+SrZyMPDYNAfGZuHK5JGI5oysENsRhIM3bu6Nps/T75YEij0upY/36i
c8p7OqYYqw0aQReyhc8O8oFkEr2B64YUso/cdZZTtPWfxQdpa6d/HOtJvrI9rkKZOQYImNttv8dT
fNC3sxIWAy6J1XF8wnzCnu9WmuVPcUcA4rZmFOj7qHIxLz2OfFNgQMOJ9kUOCH0UirCVLPV5Yz67
BwUsrzgzdup+9SVv+qWMQ1v2cTjH8iKV+ZDq8z8f9jzMTeeVx0fIA4HthIcXcbuyD9tMOmcsexqG
Us2fro9mUE5Glfs4Hjjj4VsVFWg2aQFxE1wuB4IetE56A2UFVnmwSHo/GB+UqYscI2zJeN3TrmXo
+k6ipVPY+nQTN+H+zeo48Zq9QtUtDunh3Ru7yvE0gHN9wjo6GCefID9vWnxHEtNg6esKhL8P0uom
UQBb9T3deYPUHt4DvtkMb2kV36lPCLUQjBKlQNxhpo7d6cOYXkaN5WBLiHLZIwwvd4y+dJ8pXEFP
3EZiwFbFENfVjdC2s5jjZVPog9D7NurPXjwwlW6drMxOFbxYjBCOBpQA/QQlawbc6pCp2+aQvxKz
VKz1UmDWGFEuFHgNno3aWAi9BFDe1kvW7utXA993BkJiLZlM3WvcW2ORGN/SvQ/0jQqnvInU0+Cy
wm/Cyd2Dfs6tSaRfxr+EVux/4Ji6pKdcYET06ZBVly13D6t1ECQ9lRgo+NbQGYE9oge9cnc8RhF1
VHZrGOmsKNU/5ki6z4xXF++b2hl0Rp2kxtvWUHDKzVaZewacOshvkYqtd6RgVSX5GnkUOXyGkMEt
xGjHGG1srlIGBkx1TQeVicJbcJo8Pw5cEFL1H6hDahq1KQcOwW61FyNWhJgG3KNbhRiCPyLyhrmp
yDFhAivqwC1oB52yrNN5m/AQ+MOyO6rSKQYc9fYd1iDTN60LTgnnIE7c30uzUPaFrOAgj0Xp1wOO
9T+qVN5fnOm6M+7xaKjy618f3dGlUGmgkX7EUYJ2hp9O1ZIsfjvkDGjGT8M9HsqRXmQZE7dl8EMJ
6hJJzGGPRCnaV0lEYITmxDECkTTZShFcgwlCmJRjuty29rbqaTHx0aRkE3pfe+OJknDlmMfSlAcH
2CzyL8GQLzaiuMB5tZ5llj3rHk1MXmrYMVl960J+Fs/E3jasRczqc/5cK5+bF4UmAhRf6PTHTfKC
n2whPdtXmilUh/xEkRs72a1iyYuABlW2qtJGDMGHHmwnyaMIDbwrbWF2IhB+9FeFcgIwUZWVyBLF
RL1KBWu9ViX8lClHjcbRx0ITyKNEHrEpxV2TiE1YhVQcKh0v1Vwi6S3Jx+26OoqE/qKoJE0n+jSm
lWjZY/KyyV1zrJKfSO1sYlpt6rR53UjaIXY1mLqFokfX7pV6OSmFesxTyx+rm0oc7zOjek8gVc6o
pZX/wrwl3GFiwKjQ6STQLYrW20j13h56goxGLLPWUzjF9M+CU39LPyzclBOKp3lzOzPzeBCCDbnM
TxrRrDT4izqbjFitbZzHcUE0MkZG4E5yxtq/lgLEu1CrcUe/OuWsyZPlx6GbuFn1srGyYbpebAXc
z9zAVkPNgkDsrlVjkVRW/1GglFJeSet3uXGC+IUE7CyAvHky0atnfRbsZSqHzv4MYHLNpnDYpYS+
foU/4hHxshfK3QMVohnkgiO1tAZunQqUCgOwKBgXilV33N1Rq/LdKkoHbA/HDAdRr9cMn1Syrxzl
hn1YYFbjJya++35KT9/rOVjh47uguBWR9HwePcI5PO2yyoXkd6TkDA0KIdYahLLoUEOPoTEmwwTt
BE+6XWjNOcN6iTRO7ruaK59GKtGwSG6d160+ZV9qvlP/AsR5F73Req/tB4YlSfkwaH21JWVKZpff
sytsRDEvXEtZ8c9jiufE1DPMl52APC2WgSt18Qgx7u+00LPfetfv8Ji7dY9kSsv8LZpI9rBCtm6P
Uf0UwATcLOF25b3C/4CFONCEGYudG8uAqaDJ+vFUARJo0g6Hzx1cGLpVuVos1HCqwPMwyAM48EeR
rL4YoHoK1oKy5n+sbVCrifuHHa1T1ROl9GBgnIHpv5fcLHINt4zUeBh3VNFQUUFzjSpgqwi6LGoM
ZmgNWgCWfqO8+kdMDeM2/Pv+vwjhsMo/ROUVly1P+3llt+0qz20jBv/hJ9cQsbtNJJD2pVHZJWPq
lQv6h5VN9VMXIjnrap5um74bo08OcnDQk1jfxPknx58CYw5T1rtGwRW2ip6YLWKsS34k9XPRYcxq
/oTcEIJgf9w6hqDHaiYUNUylxJ62EbKQm+Bkku44smR+aBW4KEQ0N7WwrAV3hC1MAcgnNNZT1Pov
RKZIYSaAGDvmfJox9xj7puMZhCzEQbaBuXiq9asDEgNoGS+b5gqeQIDwwEeQvinXyVouGSL6jdLq
6Yl8F0p9vuFXponLT+ZpC1p4vQiItinznEtVGIBUAONaP+r/r3ity0+fvqie3EK7edleFLETQ6+I
c65ePDA0AkC/1+2fmHS05JE6FoGnNeeVE5jC+hoVD+3Z8DpWX++AANz0EJYvTdZQcT+9rc/hpEVh
8ejfVProakYeqwBelahRQtbxtkvc9ZPjHmVHnRY3DCRbpoxnreXb+Mt2/sVIRIre5ErodNJ5b7QA
C3FS6++1xboHGp3Zb0P/eaWOk3/YQp7h4EyLR9K2nkmKu3OQIO1SiitAyLMEflwU+hY0O0IKVrev
khhLQrSdcDwXF7pm9lMsG+GKQ71ccwmpz7LqI9r5Op2hXEYcHxkK7yDxFqtvdIBTzTk2YQQkWvj4
kcvT1BBRkZOMvd7pkiWNoBHabezLIEHDjdX9OjnBKyAIMlMkzv96ihlgf3cu4754Eyk7RjosyjOC
WEmYlekb2QO82FFBfTJigHS+E9LWYHmIaWFFQr0qCLY4sd6q0/yiZlBD8XvoKLI0GJuROqn9zUry
Etg7qNcxics83EmV44k7vW24h/BMKZTkz2a8RNga0qtGNWj7U6D4t8c/B46dltaGKII35I9QbPAW
9c0DF+vZ8hB13INg/qalo2OUQw7Py9yvhVzcSn7QRj9xw+z0JkfphLpYTrviWIqG34eoTmwBfsCF
dMVR98J7aEZgjyC5toFrLQQj58IYlr3z7j22KxLjUmYWbwWjDosO0O2Miuw+IheX9Ows4Y93hlwI
vpD03dbq6uCr3gNBv37C5llPQhrGQJpR+QF3GhrFapn8FP6m3mZ0j3vVKwK/gJJOxMUEsp13xLRZ
KGzWoVWNzpcXctzWWiIJTG2cHvvtDpC8UQaFvUP1XHB40lBJK2nUZpKYX4uRBrYi+u8i0wHq2LEq
1C7FsqH/bi1GLF0mLpyjOJKAr9XYxLXAPRUw6Ao7h7vPShMGkkUn37pEHoHLEGgHirrQhaAVczr5
nNGkKeIvgCe4w7Nx3lm5/xFKdie/7oxOqGC/4RTzAxlKD9LD5DtPuBkbh969Y11zT8c7lwBSNON9
8CnohFOrg1PyGnrwHNSmkRdzAJa+VCODgaizNDwIB+rKDKL8H6EdJJW7hjJ+XKO37N/AmEWqyRKs
5fWCmGtVsQpEkk7X0CD85jOmaNFMzQLCJDcRXqH00OvxxATWbtEKJK7pLmQ710Rc/aW1hQI9cyTh
SOJIAnZGwX9SgwSa4KqkhEmLLvFryV3qLLpmanKAs3hHkDMZ0n4buh0TvvyX7pcxCzNob3WvtVm7
EtWRw/gEP/5ZN6XKPimBAS2vad+Pd3YMJrcQUmtG7My1XXZCvwJbyl6N4+p/N4KDBJkwqlaGYrcR
gqmX/n/bppCW+L+cH5+4dHW33t7kSnj9LdGmLkyqi0DnIF0LT+DrcY0FhMYgMezB5WrslnUEbr3o
kly4L9CDF1S/UbP8zzlP1Pm1SbGFdEWFjfviDYLKuCtaOiUU0BwS1C8/WNTbDANkgZzYsgAYkQ8q
0i/CfD9Vlm6+OdzO1ukslvDQ5c2i+HWAiD8GyuPPaebYrTFYOrYEizEbsNGEfV1D40brD9AHu5tR
cnFqO0f51EWuD+zCoGqJxU8HHi0HTG00BlxMTOAakTsBCMsEYAjn+5B8OQ6fVVyFwieWYyLMA24j
3NuBc06CEslAzLnSI2/+Wg65IZkWGVzmpiIexv8mXMkYP2B1TAgXkaHHLw4i7ppShQt7SAkEE2DU
yS/1F4I9mYcLd8J2pX1O5Et7GTZaPJn6gpuRLli4e8fzhfZZJPVDwPKVYCDiU0Yh3Nxko8JIaDXa
WMmaKsLselt+cacRhxmSr+mPybmemUCBExNnyONuh1R2i5DcU4ZQu+we0oPm283cgkl5tzMVeZ4D
ENg3W3GuMMTsY5fXHYjrUmQzVyOQ6QAzMJUsaxlmJ4Wm3WSlgjHVqpV9ay6rRAiHKiDl/qGbPc1S
3l+/ICjW13pT6FJL23QN31UQpSoBgnsPJyxre2P7+lc9cDcHk+VXppWePNwONdZCfi5SlpFhCMcr
SnN/LVkCQZSmvlmbS07MPjgoHQJp+pW4wjjt4+8+cSFn1/dqcjkz8Bdcv5JlmAGjGxOy7q1AFBSD
ENv9OEUROFHakMM+BpzSELJdrWDtB2FFl2nKjCEAdX2h5v4IB3b2J1uAWx/KAzgOCuzyImYGP5Iy
+Ei1J1QWfdZ0qmHFGsfiRayj6F3Beul830JX8J0RdSDpWqgdnQjN5CcISGV6MnA/rpyww4xzYAY9
8ZWkiqRbHHVfM1EuDL7A666Na0F5r5trLeRlqWszVjn/s7l6dBUD7KXrVU/CFsf54Q3g0WtcSCZk
k0zI/TDkWoERiyJ/CSUd7gB3CUbCTYymxSfeG2paCKreVHn3TFn27HP2XYXfcPqYYnHSkZQFKeN9
KTRmJpBUN/jKqcDdGqgqHeTon9YTyVf0+eRdKEhQBB/qm+PJQIbDmzE2zqDO89fkQENEx1Yd4siu
xhubxDf1VzlYsScWWMoOC2Tn+yG8ucIRN2mJmP+2R0HDolpAbxl2sArYvK2o0TY3pYr2tNufsjTE
O2Wtsn3WCEx/fTyyMx1cQatl3ti7XLEXIQcFN88K5nihGLsA821ypqG6m48TgfJ1mt11F/rw2YDt
kkNzDQFJMAq+HbZ0UHx7vjsYOD8iujESTNKC6+vCuEfk51KrbA4EyvYJFBKBWKwBY3ttRTgHUbGy
wTracKi4KOXZI+nZ0S1lBEu2RVpHdmvJUfgJKl08HIi7EkFCgUlw0XkUQAlVwWd0C4hBGHkmVhCy
FRu2gZTJfrSsH5fdu5KBC10DCnBuAXANKA0HGk0koWrmyuvrnl/9guSoEP4aco8Tdc4eVyzlOvOS
5n5pjF/tAnmequWmomcBERrz1MdEBR0DY0qaFinme2Bn9sosYeACenEXpbDAD1hWk9vWSZfkHTP7
YaVmxTW+6KXLYeEBYNb84NE3hrsQhBkFXhdK48nlAUT9meH2MQL6dPOeX1IgzgbPacHUoDQKUsPH
ZLtjLXoAsFy7xKl/azeGJx5S7GeqT9aRoaMho7B7AIAOF6de48qe6ozvRdeLAw/gdZf0RiWYPIl3
bsWbdDUaXS8cCyILDBm0omvFrHosOq2K/wvFG95Fabu3onOkDd/26ipxjH2KflBGclCorR58BKop
wTMC1PeX6Tc1eo0+9LZ84Ws1ClwYooNAbk6isB9Io42XG5w5R5uQH4/iD4RCnTqtJiGRvTZ+5QC8
Iacu+9fMJKCKbD5tbjato5I1QT0uZI54K5+z0bOa+F9Ti7IylbqrghHBMw0/DC6dSN1qhx31zbTF
ouDvM3y55dJ10mNh+mnmicEF2kK+Ka47eSRKwDXrjgwmAOF0WIk1t8nvIj32ADv066e51d3WZ/yy
gAZv1AA4WLd9qcnybR3Ej6QquqDrv6hX7DBbsuZ0C6p8kZbS2GnjNPTUGNoqkORLEZ0X09X8e9V9
40I+c2WGDPPVM/neCZq4Dbfro0JBgUj7DiNeLb17nPg6OwfP35kvfdJ8XRMsjlzOyndGVopwxwZV
lG77luiMmeHP5kr1St8iIVLCgvzPICAYBbGtzvNFyZ//sqN+mtvo/vXqjvLTN3brd1JV4T5EWe4g
QvK0k8k933p7Uxy3gl5ph3G3+B8HaeX5kZNiI3Ky44PfO01NhbiKsCsUYLegSnDh2NmfIaK7BI93
ALj2q0tjZEPa6qPDN6/9r3x0YxytYugAmFjPXI+BolaA9tysxsR678Pm6ZXo2LBWrpuA5C3jt2Dn
jkTlOGoF8cp5yVQo3GnBV36D71YCLylQJcxgH4IsD6hGjYbMzLtO2ZtN7XqxNN81//0L90Kb1eH8
8HzDOq8R7gyg5JiSSfnT+dS6LT/sbLGGCzjbnvQ8YN8okfwHeiz4bShRG8w65/0Xp/uBKeyEf4/5
k0QR1vd+swDjkqiptIC0MO4rVPIMS5pp4KZKqLFpfYKXFcpLJkzCG5oqqqROcTzqpai1DDXdygoV
Ltacef51yHnxh1Z38aQgXxtUYqPzaqaC5Jf8Z/0jwzayqlxlheuRUXj9ekUJ093OzvwUeFzr/5Cc
VZgS2U9iKsQSYE1CUTXi5Pyalk23M1w73oU3FwhA4Ezl0cSSozASc44JZ/Bt9SA51LrfkJTSIUu7
4G/f8QsgkSejUJE9PcByr151JdoyUf6sFBTYp4mOCs06BddHpo3UHwHVx8qaFyU15gi51I0ibrQJ
pSCw2CoMhYNMtx9YVGOkufUgh6XhPw00L5+X96X6qAW9ni/IAVplFj+UG7XQNqoVS57he7Zn58AW
K8+xUBROWtkI6SUDiICWTNPKr4mwz9h50h8PSzpeJWo+/KONTNbp02ZoCzaJDJBeHVOhcv1t/TGl
ZN4D4jTypPecHY+59UqYCyfrhGLswDHV1mdmtnPCkhxOkFjf25NGTuUgLaX3PPZIIscML8WKGs4G
22H5wRuDKs3KboTj/56PGP5skPAN5MXJANByqx0qdJnXGvPJHl/1jfN2Y5PyTvg7wbiA73Ei5vNV
K6+ULefwwFqRqhLUZa3SecDY52waMjyFaURvOwxV1lMhx7v+nxU8pGjlyytiSZgOnSlNMxachh/G
NVzoBDniwwVpOrJkowWWMoADfVUXbjWJsCskW6oMqo9fDOaotQicV35Vg2hseLWpagGv8GcYJqoI
0V8XJxHDWrF1+WZjidpVmF3L98MpvSKkznnQaPum2TPJNCGrlxeEK5NoAVP3i3IeQXd8nr4bTcea
s8flyLGhdoN2766HLWe3Bk7kcwB4Z9bPGTuRcMX6ib+KLgm7PmCK3qv2Yf1wdzOH3LoAl9/GxOeT
WFTywK/r7mSruSWhUKF0N9v5dDHt5k6/O9HP8GihuYqYjYNqF5Xy/dxBmHoIteP6IkWko+8E3OvP
iEF0TBOdgemLXrOYsrEXIl60k0L76JPuJU8syCZT6ZeEV1Y1+zo/9cGR7moS9lswozIgcCvRwkAJ
RvbvYsgEnCFFK3XRPMTCkPf5+YuG5yenxWIMwPVCwsN0XrdzCMGMn96TnRq90xSjU5ddD//ynQZT
4t/4Zl5zsFN3/3IN49otb76kdBwD6klgb3QFaxAhwiwOliwXjXukOBAs/nlR4AxP/Z9zUa/4lwwN
in8pLgVnNy9CrJPGk+WF0x5R/nlK1ndr1rtLf+j/RXlixRVUGCl+RhkquyXv+ddOzorQcfOdPWum
4oKGvJJ0RX3j9ag9wdnfYLlViKllXg0dMxjBFAYK93AMhIigYoNh+pVckODeSrObC+CQvqXL86kf
w/KQNaIkAyxlW2/0CoydZBpAV/iRbMUt9tuiCb8msK8osLY0Jh12vEnZsBFtWe7L7+kGyOL1c4Ql
SIe/yFuIxZo8OjvS5iR+RG8kotNgl7kF6qJVF9eacocwB1g3C7Etp9sPN+Qc4aWjvBhRgnvoHHjf
P04dQr1iQBf7DdGVIadbpbvhcwpFxczqPVVYu6xepQlgH5LvlcXqaMhszNbPuAWiShex9C0NBE1w
rRwZsA6bmgY+u2xSPyFH3TLyVin98HFL0SCTdahOFa0M7CD4D6peDUFZw0xCKez0yfV+5DUipOzh
SVrfQA7DtNyLdXIxPUwdTC+JN0S2+CSYgj+HxFbhTy+Hc0bxPjD9xUXUAaqOoekEus+LxW+OTbUd
nYC8DxsCWUahdqQm1nQvLVS2xWTjIMKhxRrE6JaMlUUdqsxfzZUF/a1dRiOHg11jPwY3SMs/PuNR
D7s8nRZdTUOFNaZrWKxX5S0ZlZt/7hywyMk/nvJe0biX18XxRxAGUIiA0wFsJ4w8J37w4/GmzbjP
in8LFQ2hYeCcjc5cd/tW3YIP18Uxf/2cywdcJJJ0+EjwomCdhP3J+oBvXTn+WEhhEAepLA13YCnk
Oshgc2/zLsYq145WHpd7BmFmRq/sPTEKHKaWxIleNKEl/6gxSBiA8mFtuOWQWa/Ox/KaKCQE3AeR
jDfF3/ZyOUuIB06WjSZcCabizAi7VWJ0uU8vS1NkwdfsU+Y1FhojhX12aEWt/eDd5YgxZAJJyBSv
SrfIzT1vqAJzq7DbO4eE0Jm7oSncg1o+GBwcQeMkbi6dhM4JfBo1ef8IKbvOAPuoqqRkBtOXhazT
3uITCWnAEmQFxWjooKn9lktKImbRTSZ4Pi7xOeuLVfilnJsRrWZm9q8lDXY4FO0lHWHgB13GLUeg
l0uerAhLvE2bNHRo64nzp3zkCT/QSPlEYzjO0qxOtdBLbbGgryjmEA0ET5FqWqpr9WjpE8VwuB8V
hvK+y7ybgXRhoDqgKM3MCtIfddY2wBaT6rCXLiuwIfuv9KNHZ0uujRJo5MhA4fZvEAoZ+0aFgPb6
arTTe18ser1w5IPatOdrRmFhv6bzFtPXrjrUYUAwE9YjgJOM0y08uRupI1sA7MW+UyhxcZBHRWX9
jo0aaH+DEM2/Me1EIqWLfStWHyHI1VSg/Q8xOzBcnsD0h5LXdQ1catKk5gzboVp5Y5QEZg3A8EmM
XlneCOG+6uhI4s0XuLfAC6xpY7Ysg+IqZsg6/ZyfOwEM8JZQrKUpuEq9y7STjvqOqzQUKbCkVefB
0JWZh55azVU5JGCWzdCkVDztoE6R5mRiilKurtojjcNHLlkX+kdItbmtWy6vHSDa8SlL5HtBr/Sb
TYs0UBKQCm417dOM9hlyhISAdEqmvAPNaXq6GT2UtnOQHmDdt8ldJQ/mOG3QEbZCxzF480mgKc1u
kXiWWH8m1TAurDV0B9W0/UlIgyHoI/8DZXEY6uQgcr/v7q+5SQdrV2REDRAs1L1MSBb1ZFRBVojj
W5kd1kZb6ameI8rj6VNjz88oA492ef/jmO1XPeeLVIZxO9s+mSjgkLvEzwsx/v3QK4ohykn6RaAJ
3ZTu+UHWCEnOk72ANIXb85SPf+RRgN4+yrOqi7EJHcmiw8HMtvx6ZbhEu6HmdXV5oo23i2CxGejy
jlmJjl/NLWtlMIbdaUC+DNF03oPGt1mbPn1EUAtblZYjcFjZCYJ27hhg4t84qo16HsEFiHzV4CWS
9laCoDSTZEgooXpuVyKoWOLXEehyjgEhgoV7Y7pEuPZas1BZsH289QlmHDaib+ry39FF8RFSyxLN
mOplUMSJNA8bIRh3KQq1l1X/oCggXXW7al79NxKxuHrYqKg/HHCimq7UxAQVi+fw++JFRi66TsKL
WCtBpqzzfzepUFU0CqKhCOzk6CMntfyClIE2iHoz60eKRJq26CAEbJaQPciSxxn6Xk368iL/ajLG
9kz3niarrdpIbgNdP2gHAOtJ1EgMLSgqvIGuX3fh23i+nnFJa4zPRfvq34AYR41x2am6twJdi3BV
jNOK1BpoQz7g95D5zlxsTgE6BTUfuzgQkiunuYVweN7BmiEh0gHA7NU6G5dZv/TEAHwDnx66+GbF
HIt1EiyeQeeIT7xjyUt1j8Mr/IrZPoZn3afdkxwa/46nP6PXFLDEiWZaVTLJvdDNmxaYddEZAbHE
LSmoTwq5pf/lBpv+Bu0KBoPmPgnwmidX9+X3RHRlnXQj8MPLeEQRG1yoN8PAUcXMZfviMpY39N3O
mKmxiLRHzTtJHIwThSrJbFcd05XChv9n5obPGnhvlKQuWg7sCTbxxcIDxz2sh9Mr7C/x8Vgr2pbn
IqWLbUrgCiRetmx1Bg+5gVf7WzuzLizOaV0Np2OCWC2+u4Z17U5u45Dpmb6fmULKI3BG0PJrNxIo
L8+pdBaLPbT8eGb596XJGRuEcZT3kcaaPjxqpWycLCgI2p7SWsbkRkBBNn6658Ro8deHiTuVCw3w
eAqb/UJnQKcw2EBZO6BER2cXzIoQwEbCoOH0JNijCdmQNrpU6thsRk59qghYpMPg+ydn1B5PVnDf
TJN46euoL2i9u3vYt7dfq3aXYERBad71d0qRp5FwFXHrymim6lGXC1BLvpV5odrZX3MApd3Aq6/1
aDCG96z40GvCLLy4Ik7PPwRdGXMLiQ96UjpJgtrHQplgIvEeNFEztpxzR8JqGHvFiF7Dm7k3osXz
c+1MxXAleqM+z6dhjnZSiIO+kdEpU4isk0OzsmZ1iXyIeMd67YPWRtsix7QqdrtQCe7K6YdRdgXr
ZtmcuVol+T1wGthHnitoxI/K6gR6YjCNdfHJvT43lKBRXTeKvjerFcwkcCXgeOn5sGB0pZPmDHId
vnQhaJGU6rqnFo+mB0HHY/QnGzTm7UFQrv7tedTMnOdNH3sIUp3CQCfa6EZvSYmwq5ezQii/7Sob
M4W+olqsB7PFVvSo5+qIdoJxjTJCtFuAaJya9MptZRduzQesjbzSN6TDIm/ko6bw6IUzIj01rLGy
j45FaMNNWSP5uC+WGOAJ5nKMPp32Mq9TihZp805yM/hbE0y2bBrt+0NeenYS9SgahkkkSKj21yKY
DyWtR+bLREK6SiF8LIMny2HZJFb6NFThOQhaiTxdtQmPpHSzBPjt1ZmG6u7Q+VlV8ZPHvkH/cXGr
JIdWMqeveD+jam28X3Lt2TGqPCKJpaStmB1B/X9i41FwaBQBXVKy+NE6t2UnAkZRHUAVpjZwOfxA
EFiSjxmTsdW19m8LG+YKE/XFae8P53TxLq1ldmRXRdC2uXaemL9rXhSsj15I1fSWXNTLPwbPV4Cz
ZEVMNcAENV7XizjHREBSp3bQGCraFQkDh94YoWgPvpkXvtANFW5bYWKXvdebo4UPgHCZkhGNYjBB
Kea9KR8l+dJoaQT0amVPKYF6HcYVAj1lZRxZnSz6qDhca2qWUFaMhJ/no+uXUm9+k57ophwQ4nTa
0US4bfnqf7wqqzjH7dB5v4nCn0w2dddXU+Hjt+X2mizTdIhLXacQUCW5NlylUOuL9u6r+u+3TCPu
qCla5YFpN+SPUwoCR1dwss9wH3cgU0iEyWu7dIwD81JkPspzq8vB4hymIoCvkptNt5GQpNK08Q9z
LF4Vnt7Pe8suMMn1RNEP4HbKx04dvrghCkjNG1NzBqyY5ZQPUuNbHFRckH73rLw4XGbNtvt9+Pj1
JQU3/HIzkUI/Pl0awPUQZnpQ9a/CWAUzHyXkC7F+eUgi5L492Q3szFOYnGFNZ5CKvMuoj8op24Fp
5QSZrHSwrC6xYvckvxQ92kX80QVV5miqeGLc4fua51PAez/NZhv5C5PIrcVC9COacIZpt+igVto4
GZ4Xb/kHXj13Km9mH/P38RmFhr0lsELH6qFuaCm/CE9o+kVBQc4c90PgCq/LbDpozHkvNvrk0PpL
rexMHdtHkwzpZcajit3WAmtUy7FX0Hlzh2tycl7sbffF1Auahad04UDlnBzSN+XiGTFQiwg2mtlR
4dSl5zgI2rkd47nqUhtlbAVpe9wOtYOkjfR7CS7WYMBMDXJL88W2hMoVy/l5XthObvctCcf5fWlF
cQ+PtUmcnDtaa0CHurWPBA8Q++XP9Y4J9wNye1m4f442Htv61Asjvg+d8Kg1Mkbc5SKXjrULTv2F
losL71FBNewkRBkUj+gEif9gk7XcDIV95VgPkM5MvoIkOwWK+CS88YMXQN4s/XGtgbdyW1aRWwdz
xEaRYRhs/ZQW65VgWG3LpJAbZ05lOMQ0ktSesRtqtnNl/c8jdo46x5hJOcrGnXfFXjssgV2EaRiG
YGYdG/eXCnCxgXptLNz8eBFPTC/AbBZLb11JV+xMrDUYQNliFFYa/Z60dUKLLvqAE2uHycv9f2ZF
iaF5dCoGqUpw5AyAZuAoVUPO7ZQz5gCqrEP/OC1RXc+V1wseXMd4wD/pV2y2EOaVnQBhX9TtkdRp
yLyNRU2cn2WmCpQ3Vm2qdeWHGJNOk4fBhMiOCJfo0PouMb81b1MapZvTlRbUACzHBLMztH7ASiKY
eXkZ+Wa28ZBGSPbwIZcRP345KzPSa0LV2KqRyXvG6c1mRT723056odzXP30eObDfOvbth07OpO04
1cfyb99pky0LUIEYYQL/Kh0mnvYjG4QNZWw1UG6v5Ng53mdB19vfZ2nwwWdbxtbhwZgkttUoRik8
rjtpxMXR+rk21McDQ2JxDdbshJbDbJsWCndjg7XFYAXMazxDSpNcCZrVt1A/AaHUo3J7SwYa9HHr
XVYMkapEBbnD8F9tO+/7FMfaFecc7l6wqI1cEbXsrlYLo6WWEYwS+3AfJk+wHPvFq8UVK/jT9ekR
Br1TiyAebJDxA5Bqtz/AsipCPN6GtENTMLShIIgTfO+oYnzDMwnLuI1Gh4qD/6ZQvrRamk5KHPCh
Ymnj72ocsLcrcGwSONc4MTk0SF5XOhH8CWJzr2/7mg47N/7lt3jBk7jRmw8iJlgyb9Zzunla2A80
/5F3GxYW1inpo6X6zpIPZL5a8WQCwHy2xS4F/PqtYKJTfCmTpRaYGLusoNgai32RCypOwcdw+hCo
4VfVn+B93bk/zKreHcyBIrhUA15LclhVlgLojA/gJ5ioQEJqrj0i0vxSj1531/XOFPqJSaaRCRKg
joR5qc5dvysyQ0yfY4Lypw2D0otmw/JlSDNsUoleOx9twpXyelCUXVIOBLrNEXjPZw7FG9O1sXea
3tRlWgrAV4Q0/Lm3A6/KK0MdQmUROZbU/OsPGnI5EqF3VWQt/3bcE3nqu2W0JfENtlxiVpkr4126
+lnKIh3+w/CEcHSUlDSEqKptNEwt2vl7Tweyq5tzbY0iE3LL9CK/RXSdyHzaSovpj7kxB42rqy9c
79+t1/cx4b/DNVZGNTL9C+ak3UXho16XZ0xW7RoBoW8hC7K+jdnUx/Ah7XfJ73lkgcIQ4Ag9ZjLM
3EQZT1RNPGMX5mRzFzASgrtg+r2SFMR9awffobBI5ZhxuAsuXAnWl/qF+zFpKFkuj/Jjs6M3igdO
pD79uW2i12fSA0zB7SjEnDNq2zU+ztglelEKr/0hnlXWPZNvkW9SEpGPvWJxGa6I3v1ISRmj+l0l
18dxxEb8M9eKWAIV+c0eH1WvUIQVUDZUPMfuUXwg64ld5U0MSSiFJEzLqOlmawsp/f6jAGDKEm/X
Ho/ukD9TP21bAkbum38ShdH431sZ6NiKKUTT0NujuK6FL2cUpMzwghaHsjhFGzcDNDKWfqCmM3YG
FLs+L6r224mC5KKDs36QBS0J5TzEHmk4Obb8UgZH/aM8w5y0M1IlLyOBcrWQl8GaL59bJy6JBDd4
ed9DH8ZLq6qdskk0tLyYLD6CZ6OsuJpLYJh3KHwBYTw1ih8qpQVFA3+78GiKO7wUemUyk1LwUsqq
3cEx+lSzrHvA0f9+6aS1z6q/KuBsBwRuAEA57QNxltHrTAYl4pRHpqbjyIScmYPQ6yv/zTFnjbW4
S0BahoMq/5mUleWCS/w8zI9rfV3gF6noc75xli8Dwh4bEuxyxduhGO0no6zXiJTJKbS5aBPd5xdJ
QEv0zcWudcogHHCk9v2RN5AiQ21K859EjGWyu2yj0o4BTZEXf5Hj2fwxXb5mu1ENqm3xdgFfBEZ5
tUg0ggj5ZKhz9PyUSyy2ejX5SzX2f00GlWlUprky+HPKzFs+F6JDzhFrYLrZg9DWP7T0j/1dZPY6
V3Sn0vHdcgIyXLSdfZJ8JhLaLQflF2+lx2AsJ9rQDkYkDB/4HRNjzkNBP60xvp+qbrI/tgFJygug
Xhqj4a0OnisiXpkB6PP6WCPlvoer60T5NXUENMBmYyp0u2K33TyIV/CkL4W7P4uZCIOz55DjaUz/
8BRbABl0O92B7jFKgFyoq9uidkj+V0po2Yyp1R+syYQ3ESb+JMoYwP9AJC+S+BMCSVQIoHrbB+qr
GZwiEQ7WtOB0gXiqBfm2UWEFClTFESb8wKsa9AEw+joBBe69rCOZyO1QGQtr8PItL6PhWtM9eEct
69qvoyfATIg2yhHWKNspZABG3QzZtzR/3jP74LAUrtE18a1RcJqJXn92iNQ1sRibOfb85cPUOUiM
xIOSJjIxNCb5dTWmRhic86Ld/Wmfv1364F4S4UksIFtX6uw1ts5oOgUDkl7KOYL9ystBiIvts8Zy
uVG+TBXxp3X5lTx8QlLMmsAnbRfL+3Qq/4754CcPAC7fNZqEMomhtQUDpLqfuKRoB98wfIMd3tMU
ZNdcew/Olt9LIh6Ruc2R3AQ0mz9zRz8GazI6h91P89VID3AFyT4GqDtzC3tNpo1PPHXqbvwMUM/e
b9MXyLvc2HV+psQYuHxBqy6yTK8hcv0+nqPlOIrFSOMbAGC+xnDOUwIboMnnPcEK/WLZs7wBTEj7
6lhqvPAEMFprHFWf0/Zw2Jg7WxkuG0yjQ1cu9/fIE1bxa5aDL7DubLJ+9etfnQMxZIBMfFdYK8CV
Mcpbir4Si1nTsIJ+X9F4KsWHquw1aMVrWm/9jnB1VYZoVV4OL9RVQqVLfLHkmia5uCfT78KIoW7P
UgPXZhm87mKpUBAZBY1Eyb6rNIZ7Q1D93wb2KUxvXTdqmKYkz5zNIV09C/9cZ84HGmA8IpC1EUa0
Mql3xqL+eu8z0EoJin+DXnLtttMVHbAgwz+P2LSnXyvrBfkPvbsPTRrNOwi9uRlotWs0eafN3Tgo
jkpyWorCvbfRtJEHbLPGHOWHnMzYM0UltjGhJBaB4Tsrsisn2w/ZNQRP/wvFFf9I4JcX+n0y1Cyj
12TAQ5otewRfrCkllkkJUsWgQEdzvXAe6pYzPFAjA1vZuYe/2hj7dzsnfcpXh1/HRNv9z45CfuTd
hgCGA6/+xAekaalXLUYMqm7DC4ktYuds407NB0OD4BGOLSKCJXTeooA8hqJIub+2ffPrHsVvLm/o
AAL6gLlZ3EnLDMXoUbgmfc7LQdvj/XpXOmZYFRR87DPoNa5n2wYcSXHAcFUWfx4TNYiiKpXKiXop
qZb3Qt8GMdDK0BBgrWtVqdeyq9rfJO+AFOxihaQu7/PYz/nQ5qdU+WfGZOB2B9OXbCipS1oxFxm4
+W0Df0kSHfYPLJBKRt7kN+jmapbd3y098xKRyAfCLRGzfNCqPZBJD68Pe6tlrY/rPoZx3Nz1T8No
CaLo5d0aLXubLfqlZs0HCkGUOfR7CgG7CWlPvoNi0xFziVswa9eVXQ4LTvmPPlI5CMkYHOjOELKe
cNVdkXAdthdXbTJ05PqjJ/dvFoii7ToN/DkgxC7yyKr9JGbSepZptt2wF1N8ZnElTBD7W6aGSTLj
UbgBjd9fvAGR5HRdMSpUFiN/rcNaY5x2ZbbPLoNCNOwSyGy1knY/r7Pv/BUsT2+118TLJ/ukFBt8
YL8+I6k2LRO4r9sFGn9iagwxXmKrUUlK8DwshcsyOKWeMcrKfrBh3WvOrkzZ2PU3vIw7Wfi1uRSG
Hv8pQfSkQY9fK5X9lJLnzG0A+kUrDwZ+WYkkayorDtjWEzx8jut5Vml4Q3tqAlSX+1SqvcLglz5G
8Pfw6VC+iTaDmuuN+IaVfHPAgswymfCHFir3vrP2weYSYT6RG3VPM4I7uy7X/XnCmEMm2LbqaUr+
/zVvMiNJ5gNr6fkDJ/Es9E/RWehyHk7xYUIuilX7Svz+UPdAtQtDPmv8xrWk8siSd9FTTtkK3TXS
NpeqOEcqUmixEji1OtI/CtCf2LcXibDYjSo/ccnxZJkYYcOzQHLWExN7RNvdQMJ0EEYKRHXVdw8C
mIwarOogGV+10wQ+ZumgUevx6cwKQ6ZmRxyma/d68Py6k4tTa+jdw7qx9awi/ByTr/6mnV0ZxTJO
XXJwuxCmu/KJYUk5/V9DmEtrREzJDGKUL7SzlAZn3GR8Mempzo8Lz1KVCuvnxqjczGUWGrDOwRMT
VQYTBpyI3CVp+OKk2vWifOjFR7Y7Ccl6ZSOD1xHePUyEk1CZosLX43e9ortFRGkUmz+TJJYiFmqQ
MOYecYQJtmgsBDc+CtTlk8vz4s3n0iLI8oc4zS6l1raKjdi0DW21ZJ5Nm7LkZ41J8oIHE0QkjUFc
PqzpUQDJgYPLthb8ADAQWC61jzNGMpdp0wwWBNc8jcJxYixyl7IApIPBtpa+GcnbLIZzZHChwDG9
fWnxLpx4V4voB3bWBIfeZFc5szK9qpnwDO7mfP9OQF989GABG99qKIrn3f9KEIJVf0n2O53epooD
aS0RFCt2hoPQq+vyc8Ab8H0wq3i5/WgFq/fsWmEADiVJliq2EN9kPdkqCCfPCb2rxGOmAt9w4UC6
GtZTU3luv/E7/qlb6Xr7MZpUVq89lU6V9Ki5pu1hCVRoC/GEaRS4UMIdZ7KN5xXWGq4ywM47T1NR
zprfnf4oKiKm6lUDznkgZGsMrVQPDTjV+3pdw9LAIi14/wx5gM/mSzIFGY93DZTmkhIbN18Xo0lF
71Cfjjsaku+Aqi9zd6lCo60H0fRpi3n3l0/nm41blxIyfwmR+RuegIhBPL1rGXH8Jm4PcSloi4II
v+xgnsg3nxX2IgCT1YdjLaN72moQRC5FnWpukSOxotP8qGHDu1p1CULOBYUQ8Mxvm1NnMHt3FWeE
w+x8fBOL6g1anMVOpPpoVSnksxTZsl2qnKsk/WN3KuDfbx/iaYtc9I8a6hHLmebFSytr4E29Zcmv
DBn90nahx7Ha85EIfjtLOf+ml+tG3QjuSGdx+1Ifh8YGl0TX0FvZYqGTM89Ucv67AmdoI0mVMxVP
Gt99GNzAzgzzAzkn2pXDIwx5mIUVN5vJoduCMVzpsNVeLWJcWGj/6rNKuNW5w6+eEKAu8yU/o3cN
sKYz1F9eI9DbWtFMYJkucq7tn46FYjN9kJePbI0XglNVprycxhmXd4OH7YoRWa6YlBqXQmiDeE34
VWQfNTcXXmGThg8kqJd0ju+BERqUvp74nsBzN04zMlpkxqFt0gxAw0Yld4BLV9VwAqSnDQ14xw0O
eVRtiqGpsgZfSWCxrRYb2hvw8krhKHVCG9qhKiKbB2FWiXhU2e900+fsqQRLGKRGXZVWXV4dXBPC
GRwdEfDPCyTGj4tPn2yzl8B+byb8FEF7l1tQTPcVJPJfEGC4eqjsqvoecrZmVDMWBEUt8qqLvj7w
XxaR28WVjibLmeRH/UE3EmD09ZPwVZKAeiP+k/ggXpP3bBXoGyXpZOVuM7JiyyRO2skxkRIAhafS
nklehLY7OBQ4iXryXVoGU2B8ocS7Y4LGjLdzgZaCJmhmHnifBJ4l3g2Eg8MBrkbHMBo8/gD4uWfS
W+q9MxXma2KhH2d99CJRmNxJF70d9aCZQW+M9I9zZ1F4vtxhCeyLfXndO+gsleH/9kBskHrU+UmO
/TxpZxUNB6ca1LDkFGVx+oBSTxdq2nze/nV0I8f5jJlnuWhYkuiRC+85hdGyrt8cseGTAGvunjUi
I9L6xtnuwxLOjQ1iC5zk8oO09IctddBK9XGKAV2fhFxGd4APOuE7Yb12rOZf2GnZFFk8Il61mKE8
wD50fu2/lZT8rDcIHRm8E/vGRn6fMoeYx5ioOSV5I6BxPdAaCJqVXEtbUSy554k1cfOAqNjGlt+P
ILSp74hpI4x1t6HpgxgqFAnGBvK2Bboc3P7OjgvLG+j8qM1fyeWziHgVohS0G73JY2O7HYalgI4E
EEnPdDBRhqJ98S2+dmtXSHQdyh/2L6hqajUdsqZUgnt+T+TakaEcmNuEZsLh0e/ABZajdj+jlTpX
GYZVlcjw18gPUv9R1riy2d23bYycGtWdslMU4NwpgkbdADXtVT8dUAEyh6JXovu/QxWg2ut4W6rK
NrrGwuCf56ygNOj7vPDWsgaCG/TYQmwiDIR0RAt47kAEwwKXZhxgo5f578iWFRqk+0lhu6ZS0Ld1
j4aVgbSfydqhAAcD+0l1JxZYdRW43J1YSV354DVlOIzkirw7fL/bhW+TZs5C3pusahsl20uaN9fx
m/GQQZP1DCjREpqbQrY/wHvhOp4wEcRNNyz7Et8WsWoHdCW4hTMpGusU2I2ieQyMKz1bazZRL5aS
7HyYihfyR/ki8ORfetssAVd8swHJCWYbxO2N6U9cCVp1OpG5lr/yk1Bq6FITEblBDNONw5nADEdg
+3A3H72/WL8XHcvsomqbW5do2hsE0wycCclHFKXURJTuTKpTz6NcUd6cS75cjF7MTxr4aC3MRqco
sdKpiitHUsCD6kKJva51/ET2ABki3Ze3J02H0/zhXXkE6dsB9ZxyW+grNf5G9bgR5ld+kJmuYDXm
yafirGgC/uN7+5OUOWnl9lQ6bxl1yim3On7bXEfutxciuML+sA0jpBP37hyHQIhFBiz18F7wIqWi
tGxL44tnyzv0NjbVfwXX1Wvjtzewe0YVsisqaE7tR3mNB5vdb3YMRWgl19plE9vjddzqfBmRivkh
M9OgMLw3VHWJosaNx1yg5j6g6hnu0xMMzbUe/pCcYRFy8kH1mZBxtAqt2s/dgqzmWraFoDcrX9un
2lU8Q7NZe/GI/p1vvBjoOaj/u0Tsfpb5X7YTk4wP0eEmMEPCCU1WTPS25xUcBmyyIbI6cR+b1v2C
ZK1Ujm/7c9IsSFVtdNR+0a4QmsmdJC3aIWEYDwIDgotJyEfS8+W9Wloe5alSW3rF6rukxjibwSgz
i6aL1Dveuc1fnCxEOsimKdVJ4/rOuv6q9kxmVmkfGrUuTM+oUa0iEHpJ7iEF0+Sk41i31G1AzSqz
BBQS53pV3j7V2UZUrUI7WNe2QbMGXKyiuGXriOCoycyc6V1rgVnpPXYqjV8VziQlm+6qY3y2hMr1
SUumnvklKDsHCqYcb/1oHLVm+IzsO42XXMuFMKyCYioswhmMBuet7z36YRjBlHBFAgDJh6KiuPlh
W6e0d+ltknuHOGqwoEMOkrMfarc2TabCs1FA4Zkoi1yZ2wpIcXXjKK+ghpEgAFMxfCFbg3q5CQF7
YbvjwjUEgQlLylh6GsgvEJg3EJqUyFvJSJuTc1xNfoc9e0+vEjuypEsfUz1tLC1HJW5nuZ9YnGHW
TvD207NmJsx9hh1hnzkgSnVFH2IimAx5U5IsgU1V0StNJ2/IQbFKTkcQ6kFEEbTo0x39yesR3dj1
GqyESov55UoPGawdm4lD60rq0Os9w3Tm5I84ZTiAUaMeQCsNbQ/Ch5Wu9VlS98Gg6yLjcIVe3TUK
KX1PRW0ucch0TQgjAn6Opjnr+05JRk3lKW3AbHESx6QIf+C898O2QRfYngQ9JV+i7OWP+YDMRt9q
d2fxi4VjgsJU2TJ5rIccRoLnaJBa23fIcrfJtW1NdVrmym1hUEUMKY0iKWKG5XLV7vrZQaRhdf92
oQMp79IK5iRYZEdGlMPx0tS1h97IzEap91z+dso0i2Rx8YDeW07wWKoOwjX2W05s3kMGuMzKL9/N
3gD3y873eRmSUSrRAOjPNwLThAj5gUjsHvPGMrNuEwy18fOPaivtI8QBPUgNjCOZjuTZRY/1apfJ
0yHasr19vgoMIll5oQlMWXA+HFS7natD9pAY3KzKslaNs9esuqK4PZ3Jox1XpSWTmQ+Z39RE3WRA
2WvBHSOikubnM6UF1kMAX7XnNwwmXDQPWZFQRzisjMPgZaMKXTDRyTDJKIyJ9uD2Bo5yCFXGNfIh
NNWKHCPR/sVcZNaVlwumBbRbXJxwGGCInEoe29lMY9W1QKSxI9x1A2u1kVyIIG6c2pJI2urHQwC7
nO6rzIVwHTKJ16yIg/8w+tc9uTuG30kq5yqnn4rLNEt16CrDHYE+O5q+kzndFboizcYqvvWpkclf
1eGQid8yEuOw6rahHPze7mrKEGDe2H0xZcEIVYetKjMPK2ukCd18S9FIUO2tf0anJi9GJq/DbAY2
FNNNH5R3jt0sgYHu5noX8U3DMTZ0Li/pIasqYXWzShwfD+vWYxtgaDJzNn+aTdJmaYtgGgnoa5QI
6ZPVg0a3MhK3asyk9ekn6zcXWVH0NFuBa1ZgTqlY/vGXTUEuRXkGVd5kg92Oe+VsQGHcRI2Sf2r0
PBao9o0m5dFuN881Eb9LWvOn5GwnCRKOx/DxvBiCmX1M31sBV6fNmwKh+Bz5RVN2WSbpqPOKWmeU
zLmBlWdl/Y17Cb6/d57s5QQ74G1nX0AI5MPby06DqesPIdOmYBP43yjzbn+VXom3GePkxjTFk3gw
QuMASOimjyqpAXS6Qu6z3ski0A3IUiMXCMd6M6IXCNEpDf6/u3lHGnsVwMQB5v2Sa25ug2iKt8zF
P2EHeOBOB7EZ/RY4QUj0uH5xbtFtw9nRovncx6kSbMUe/Xw+5N6WGjQKxoE8elmTpi7RTWJULOlH
xiZZj0h5m1ePAjc9XVOnCeVuLsJQsdPys3Dwim4nmP2GH4rjrqOA2wRFNmTC3OdRm9BpPdTYEx00
6NTLzJqkL9UCY9GsQ2QM1M28GeFglzA//0fw9MCKgudLXjxMS0RxFrgLNaJeidyXBdULQi60uFBr
UYNuPaw+dvghsznKHnjOxBWyFJWXZtMpcPbRO1hcwf42yPzVGZNqaG5pUxtigCVs1q3ey2uU2488
Y7eVhJ9onbkayghoBnhH7tpVqVIurazUQqFt/U7pEjdkriEhssNdrCaxO5tsbOXyLiQGfDTgVBBD
BOoiYfi0JM2REq2SQjkPMc5C8CidqtCa9lZhotsjBJ/XR52bQPMOvrr/nAEqSwvlqNd2VdusHpFo
GLk5lLTGpAFVjTJn+oZXDzUpPi9c12KtjvVGaCt9qU26K25l3S19VZ8IsTiQRPtiHYzHuw080OOa
frOim+9pjcK/tce0o9HfVHoP+wMUWR7R5gwk/MQ1ZaE69csvcdVygWlmRcl3jdUyQaHJJpf81CoY
hrnMQpTxCMkp01pen8IKMlv1bmRhYv8m1b6tGyvUo8MnWfVxBJQaTjkbAb3vswbSffAgPNTVkALY
oP5Fz8PFKY71Faf3leSvGy2DeDQDNY9h8ZYfkGqe0q9bum0t/OjYaVIjPxAqtZiXiCmFtuMzd9gI
wkV1gkQCBMkDfm3vsMsEuy6w+39VxBBWuTr6T9p4NQHitifQlc3XCufhcjC50U0IoX6xt7BoqeEi
r+FenGn13vBSYQPpNrej76ZmW+c4Q7M6ieqpEavEDcKaVpPxJ479gaeiLzcNniAQRBV8sv0u8L4E
MlgZFCITbQw7BSq6B8r1aW8Svc3PgMO7OPWJxTjcF+UDkePH6kh8B0kYJUItShsyDkVUpPnqYHXG
w4xnQNBmGkoiLaJ63ywMAVTqsC3Upb/pnFSa6lTeRwHwVyemU9MWTVx4mT+KxGFfClcGKdkYzp06
RpYvijVWYHE1Ti1p02OQ83kDh4qV6WnFEntMUZipMRy7B9Vhq3ydMOIeom+HAYza/vwcYPK4aoHG
wNWrMrWqC9byn2/I63wg+bXOo7E6YpefghCI/jWq2+slgd3GJ6kWOZmbFTg/Mc33kJNl9uo6nLOw
rdjZyb4KGHn3NQt7ANiu5LDD7JrgN8r2t2eC9ZaRp07adSbls08iE+KFiWOgJAa34NwKVTfuzE0F
0gf8jV0ssegyoFzlcJ9W4mr6porGSllNSntOcinc1zgA/t4f8SjXX1NvnOSPRQ0PKlfG29Zg9uaU
iabqOtcPxz2zCnKJwvAbpt4TGnxH7T/5j113beelGcaYWpY/RtuEie178PmSZ+k/kVRhZS5hkbuq
qvBCzYb8luHo2pgIhNGg+bb3ELmzyPV0IdhYKccK6ZKphja7f56yGhAgun956MaQviHG/2VQK/gW
zFGb6/Wh6buxrYHCBLg4VzuKsLwPbyCk8PlluvMQ2pe10MYroQjXLijQgGYWH4qdSAT5iXrp3j4L
MCQ9KPGBshYtdPfwil8FFnH6suNoesMPlOL9BfPvTjfAzGoWsrYm+UIIAglMzrwG71s+ZubZXzz1
4NqaD5xnalSXc++/SvcaENAW9qdwxz5EXRF38Zb1MoISb+q/CA5XwFc7QgBPL/Z1peU2auZQO3OH
16jIN+EOfHYcx4RKBICfEHx9unod33v9fGK18FHk53U13Wwmk1RrQSF4fd3aTmJvE/O96LfPfBYc
+QbNp1c4nsmWTz3oTOAETXkf/q4uiHYxQ64S/Ruk8ICEUJAZNTIYxkSGVqTAbpTN4AhNkCOdk5Pr
fy4+ZMVByLlnhA+BeB1EDS47EeUKUpND3jTCQiGU2AJRU8yhGC279cAjmGR+NT18/jj8dLSgPCKw
RyNV4sVyyDt21alTNbXPk6b1JbBwXXpQwMoOe92Tf7tLTQmv4egPaXEnTdNoJ8FyfEBsevQfgrBO
f6lJuXOzvtSolQ/YSRzJ2YMxT03FMOWPnSZ97J0+4+6O3o3ZORShZZpVQorufbdMpLA/zGl5xEax
34azgHcLD0Sfj8d9g3bfZCDJptlrDCJTMq5iUwFEL38vfajhDPCxdQSqwvwFQSQ7KJi8AiQZCDpM
BbyR5+L+7U/ijSk1TOgp1mmgJ17v1dZMWhY4ck+UAGvAJELdN71CemBKlx0pLTlW0crDH1YPzwTz
vHJzlgo+vFDFajjFDymPhSl29EI0fdnrNEq94PVKDzKG1Qha0F8qB7gCbfR8Rp0WJeH6q7OgTf/l
nPNxtJZzTvMHng/nPszfiaOxg7QEeyGUpNQt95I5vsfKTqt9731OlrR/9JoWsQeGppjceE5PO0td
vYBgr2X2/6m+8mkFIiXNlhVKLpswXJYJ8AAZqjYz2fiv9T0ko3jTIcW0+TMq0ziNXrp8FaFh54aS
GX+R3D5kevI4xCskupjuX8a4RMSxvvDqiV/GK3ZQap/mDYfcERlND0BOs1kVK1V6il7+sGpvz2Vq
jSP+NSjSal+VhaQWoqgOAlkFnhOTl+jw5tdD67uWAiMt/Erm0tcFmGB/m0SKLWGNCWE0lTDMEnq4
/kHQJxIQ6gI8vfIoMhA/qy+nZF93Fc3r0sUyR7OY/ePDGOmuiQNtnMksgEDpj32UQc/C6LZnJKhV
kcvu0mSRP85yb2w+secusUrGJNLZq+xxU24ygkIYwwjHVp01EzpbU3kZxItU/82rgGZB+jwMEtvI
JrQmTHPDnTehzQ7K7dCbnoG2F78oj7etQCJ++9eC2LvpVYMHcBVTHQ1l3Rne5HmPDb6q5W/rCVPI
fX14NkQzaXMRBDh8odcQ1u64gf/dnkOrnoUtS3LCfs00lEDCbaeun2uYzlWnVinQAYiymj9yydDl
70D6NG/Z3UMIOwM5Dw3kLrjMQzkh8BsEl0N+36qLVxedHre+xQLKa2smwDhnu9K7K386emcFlAry
ogxL8OuJnygyT8UOx6GGagtNCvwwxE/wq+osrUmvUQKQvZYcq13nY2XlPXjNlOaLeIuIOx7WxU7c
hs8n8CKTNbACxd6QbMkHWOPDmQgT5g4mnmUAkDsQmC48G8RSGYeGwlh+o/bnyc1yWVximVXfv8nQ
yfUQSo0Innet6w8CsJIcDBJm+idiqfVdlptYWwRwjocK1nSXVAqvBuqypYxSqPO9/pyhlcoblX1j
Ib1pw8OlwoK/M4ZuRSXO+CLHvyVWATZKYn5+9IP2chNfkWvFmC2QQNjvJd1n+yaEo03ab6jRIPta
AnDsVWba8LYIY9zoaU+x3pmwOBaKsDAD+88JjKbKOq9Q1GP9FTbUXj9WPinaqI1mDPxU4PiiLqxd
7Y/0IV2UnFGyZ8mgdLA8rYOstljcxeR71Lpn/oKfr90xfhIJE0aP9zQd8ifFiG0uXvIT8Kt8fJHE
7XlEnXfUBxRR+GOtj45A4Z3QiV0P0Wy9lEqfRPItWwg/YZOPmRLMvPtB8ntezIX8uo3tREq9z/gY
eBk0fAm2y+tQ1r7ZDHduI3etdNFEsZOUl8rJ4Sdq7d0g1vvWL1i+1wq+kFBJ417Pq8whkEVIAQL1
IiwW+oZQMfINshiRjv9e6a0mFCF0t2fichUmrAjTGi1QlaG5Qe0CbomJ6eJQ3ueQZce6fhwTV1cp
CCqZ0IUjNQXTTfTekXZPu88795B+9hGYUfeBfAmIR5hjZeGGt28Odr1TmvMnLrSNBFlXhNJRpA12
Yr0L9OJ6ttdeKMczMTEvCgwwLk7JKi9Y3HEMYVeTG1JP5Go9+ZZtx1AR4ylqEjXOfAqXBq4fntTe
lWYeIYi7d0oVGjQUy0aPH+mBAQ313SUpWU1hKIB65XZj2sekS2fpLCBFMsZQ+HnKQNaK658aFHQW
1gzBth6UDuakQszATfHA/xFzsUISehjSiPm/LVNPelUV1Gnx8uWy0myjm+DVFI8uy2V2Dy+TlWlA
jEj3NpK8hg8L93t+qCRu0OIKXMwavJXbc3DgsbnClhSzRGADTfyOIT2wEi2z7DKEr8aRnwJpCnM8
J27M9Du1QdS/zllNq9zizU/I9cvc14YO9NQdK2vkK8vWUceEFsZsUGp810j56pnXlYOhJ6d1rFDn
DK9aKXZV0xd1ocCpeyTqTznMc2NIlSl2pcCr2aMfKAusEKZwwBi0tFY7gxbQgrjxGfeb0kuC4cul
2CKIunbBhhF7dSY1sM8fo0ofb6f8P2BMYz6IomE68vE4ZvIijpH9FpQrBf5YI4AoZ6f1SvZHhNMZ
YDYfonDEBB9qtuDSYdrkXtODY1EHB9ddgbpsfa7KKaeQOchArX8fCnIL2Z0fsM5q6qYzieulcW0e
uQ6TKkcASyqu8K4OHetDEtOyk3vBZtwVQwWGn/yd0nXnVRqTkw/eqWocRkp2DNFpMZ0LFQ8icnKd
WkxZ+x1IQGIDPbOv/WFgOranUbM2ht+bVqq834UES6GFrq/brumSqHWk2qAeOdeE1cvolI7M1cY4
iCbAZDRIQIRXL/8V6BD3lCIub5azds5rx0gjKsxH1o/2GD1obvN2XlKWmA9aMdnerLwNdinu7Gdb
lC1yTip+rfapIjcXpdUbCO0n0Lg2LgYH0tDcvi0i7VaA8zSS2rX2DfNQBk9O8GOqpjTiSNVhmeJ4
9ZcfATQ1YX7OxZuBebZeedy6anvnv60F+RKdDhj/z6J96tUPyWqigkaZ0jpnOMilOwv/dgmNkKSb
eQEbxDJfkQhD3S0gTXFPkmZBV0nHymTf3Z4iptPuPPktaWmOLg1bNh4pKQXCj+c255p/0X3kNEpR
rUsmpwueux/NQ2+dEnLdEsM9ENWLOHYic+nV6GNPCXSs33+WNKixpkg8lLS+XUHaAKAXWybzBPdo
2+sHroWX2WIzx8VRDmqFLKtwCSM/HXbsWCCIxPGPUidOsvTFiH19RaxeBF99oQ/QypqiUPnIG4NP
rM56xTvtciwAVFj1Vkux6pAWY7lmT5ujY8PbfJS2My0I2++kffQo6sPiFEGl/LReXthjIzPix5QT
O013fH2OTldcGAoBRSvyuoCpNDsNJp8MRVkfqWpO2pds+EfLB1+im3xkA2N9JMYpybE14ZuFeLxq
2gptJatGUYlcp5p+qhhvWfb4+XcuZbmzqH9oL58Jnt10TjYBAVR+OAZ6ereEmxySFvwe7D4YFVsR
9j/C25Jg090wr3jdkeAz4uetbsrHAn6MJ1gHWIne0BrjBTpIUWDhyb6btDuZjdRUlZFBJ4p1QZ5w
bOEuSSB2XiD6kJCj0j3h5nZ90ABFOa1cK6WRp2+K6VSiEPeNRDgt+55Y3gkIYppz4O+S2S9F8s7l
mJ/WCgz24OS9Kf19zBT87UZkPH+1ntxv4yxHtpAT/fWOYHLsT3OUCCKQsPn/crL50BC4tJpb2k7Z
ZosIdb8PHKsbPerzd/MR98fKV8H1Y9VprXM+9RkJBgfjFlf73JXv+DodvQDvrugo8tdbhsHbYXn6
9N7Wn7POjB1fgtS3im1gjGiNDdpnlTR6AVnxIt6/FE7sT/raguSC2lUo4WYlE71uH5PjHSMhbtH7
8EKOgZlyF8XRHi4bjiQUyIFBWA7xjxeEWBbdYe6/LdWTtf7MtalnckHo3z968AgfJspe2UsHRsQ7
BUu+nFp3/dVqi3B70bUPZuoQVH0yzVtIQgV1jsEsCoREVj5l7tRHjHPWlTEnVy28qu74NgX0/qQZ
kyy2Jjn81sasG/IE4QAVK5RUvu1GxHeUwtayCWx9cH49nkWLQpA9dxi3KJ/zfpBg1SSL0mtlfM6z
Z9ji+S/Spk6njv7wSRAO89P6TNhdVp4j5hN/p88kOicp8U9vTcD1L28RVju6HmDXc0U1HQo9HuDQ
lV7cm6x09dAKLYuScPnfQsyVhop1YKusDdzMeYqtyeyUw/h5/ejAkoekzsz5MBwv7WnKGBEcW1bU
jr3U/02JdVrnYkcazaIDvlv6h/Lr7ognvnClB+q6+zBVNMKGTKRoB0pyvJj5pJJ4Il/7b3dcCY7g
NtyHuMC1XFE+Fe8QhpagwqXTRb1lUc/oG9JJXsD4coha3+xCuIFEmUfncIAhxrpnmQ28fiwEsQkP
GefVJVvY/3fJQVOspX4DOGpwmxB69VeV/Sp5YxwHW1ngBS/J29tOFWS2zQayNlY6T5QmQ5qQlzeM
q/io7VjXKOkZza66+fPTKPeWiWdIJOU8zXMYsupklD1QAdvxUmFGKWqiSUiANMKHaGj2YqVaLfzC
5LfZE5nDHJRATdWfch4d+EoEQceueFsZYsH8yAcfa4h7dTTB2ES3aoWKuxB3P9F1E5TJ11cJDHkS
07ZKl1w97ev3CLJBeXj9ro91L9iEswtFH4ULKokkWacTijV6msJSAK9N6RdLxFUlhgFyIOXTK7PR
xfnj6EAQOBNBDTEgMfMtiM/MrRY/VAGyFrVNyS8CeOWRni7Svbc3q9d8LullWY3gIN1vU+ACIwhV
c40BwjazVFz47iQPyioOwufhdIUkgytWQH5IxfnBhD+0MdY/C7/AnukFfauZKSBIYQeDFSBQfq4t
QHWLURs0Nma9xBH/qcPtU4egE4/BfnI5FwFFRj158DxOpx0IFPIwMgKn/gIO7cDibWDfU38f38Ar
cxxlpB9S23A9SQJbSZPf0TpHkpwQLLqAt8Ab2baBYUvnNP+ZiPKESCjQe/m4G2KZTLCnX+BWuXLK
+v603+CSTWC+U2/bJMsofYpedkg+vYYVCnjIZbRfXgVJMIFEl6hcOUs58+ogVFqxToqZ/8MmCEy7
BHfvIKgsMvBTthQ4Vjpbx/UBU/KsMLI8trKthkp54NM1UWlkNkuI/P6wGAvcA0AIl72f+TAPazbn
3N8SifUT1IWPhhU6rKkvZJq4X1+/4FbEtTOMrZm3i5Vwvai6Op53u0KpSTNedi9bEJbvstJHWy2T
hPuyq8InDukBX3+a3YhkROL9ud6YsJ5kqTvTW8exKHxtjJciN2p3WdaAsKKta4dOdrqgS4jNw/Wy
6fDibv2Y0lm8mTV8dJZT9bB2DguJFy9R9yBr53IrTEvpO7lnRCUElyV6k3O6V7lAmJyvR45SEOLB
YuTKh/a0NcNws9QtQX7R4KpaxyQad1n15x7Isp/ajyRRv/mZ+E++TeYCLUXBvtkLGz2LIt/Zs2GE
bSTeiIvuwE2L7C2Dcg3m/WtPE2fPMwASTOINa/G/8aoGJiNe4dF25CEv112OMxHHldrO/6LXUzzN
LKWvImG3s7qpJgOkBoOGJlkkDU+t1VEPoc6qqkXwWnyD8S8N7DU4iwDek8eeMvOWgXK66rU6z0Nu
yXm3mksh4NeRn4pp56rNL4Nl6zLf4kvxYqvhmFAAeGo4nNi4lSWNwMoPjZUzGN6Q2L2RcLf4cY+T
dYIMU7s0Bo5DuHBiopJVslgyO3inNfyJsOuAg7kzneZ8jaoIvfIPTSOR6k8ptYkR3UpN9e9uMP1X
oi9P6DkCYEWTbTQrjaTW5bS43qt/I1/ploVleJ5k/BATZGiD0nltzrEHQqLIpJwaDN3uludoQkfc
MMTyBuFu80GmMHBbTMtZ5lqMCBHlFZEIvnq0VZLX5QICUxpoY9eL0s1gXQC459nc79FmrAI79XNu
WDldNmDoPzJoBgU03WxxqRe7YUdjV29qqmm6D3eLWVuqK1ryUPDoes5O0qbFdkoT4U/1fYu7eWhw
O3iDpC5w5vJwGug4pNW8dmR2wwzWh7LFmUob6gsezR5GL0sYc5MRjuKbvZ6gzEM/HenmHP1iAqLW
9BovEhHiJYl+KqPugfBKqdN2aY5O1VkA+XeeW1W4aaH39aZqQLR2iot2eqL2SLqRC1ilXc9ZLtKd
NEKjJVbFzIGhS8treM5IM5wYSMARy4srB/wycqHRi9qia19H3vS+SAw7Cuc09NayDfPu7oV757wT
HdJxUEHPwXrb3mtUizwnYMqdjr7ZCq7VyJIIX7CkTTrKbNUoytXgyA6+5+513GZ6gTGsVHIXDsL2
KM8zi0FYzruT9Ve4UzXki1vSEoUvCOBbNzsoS2+KvJ6q/T/qdqhF3+Ed1ORKWHG/FjzY+yoiXz2K
I7ubSHxBOMj6rXyNj/CYijWrCkBpBnot6vOS6sGuCN6MxYndBh8mqHnTHGZbo9qkCzKOmMNbejm+
+rVJh60lQf1mHFAxET7KSyRvzCaIS+lmOhBxgaS1LRGuVPZDyJ3jm4Uay8mOPp0y/H3gV4VmL3k7
DDOmzKHcBmRWUWcvoBVdK7fgqLRL3ZBWHs1BRgic8gkgCkS/RXluss5lpyFG0UFiTkD5aV/VL7VW
6IbnsNAVZQH94LxKrj4oAqBt2S6V9PIndf0rq3hwAmgqtEFTsl6fBY3bRK8OUV8XTK2wvDk/spqP
dyyNpQCvGVRaU4mhRChS/d8YnfizvYaGr3RClKGnjZ8sx4q8YYQm2OHoh7eYMoDahJM5Be53XgOv
06hwOZDYXnSD70LXdD+yVowBpbv6p2UYWnNaSjwQlmysDlUABw51Id4wKkyP/q/PXTpT9ch8vAyZ
xlW6w5hIviscNU0DZ2wYly/sE1I6Ir+2IqRA1JivztgHINyZMhes6FgZevBkiBpsv4w+37mavags
X22HGCpPEt7KOA7NJ7Y+7TZ72daeBHAalMfeaEY8EGHQ3qQm/meHBQ/Ljv/brk/zvltUn8BATwcO
CqBy+2j23mvAFbrpFCQZvnixNQMmpjV+C161k/xw5ojwUxt21DJO1iEGXHcraTr18P5+pJF16CCB
gvImzd5u+cvGiwUVEne59dSx91Uk5wBrKlnmWU2dBc+lzwtvjT+YAhmq8gj3cScfbI8IjHoHS08r
SWqeTaRs9HStPRoc+SbgT47r3W9L4FRr9WMYE+bPnapHcZFzs+j4j+bKXQAtECD3iLEIwylKyI5M
dRFX0vS94y/O+1piG7AiYQvYJwhwUSCnbI2m2LQn3JwV+fl69bvE8wxVBUTopialLx0M1RIjg/5t
2Ap9YKHWK/IcYieWwwyxvdEA9JCe9DFADTUyf+HuYSKENcRRp75ojpTpSeXx93Xo7PZsaj5PnHo1
p7HPCtAia5u0+UvARoy88Z7TVZ0GT9lN84VD4xI7gH4mqUd6Xbeo+SzydSxi1QCBQKwzYdUxyCSN
ZpCoY705iZSXXkTUitshTjSO5oUYrF4dfHqwciYvkTHyWKnV7nXMIQTZRellAhzxvNxquYgFTyb5
iL1YICkXoDjs0T1t69sLQGoe3HZPBpGOP6gt+9X8UOYJVRZrlcbQVf9VkvJmMRiQsGKlRP30KE3A
5mOWb1yF266XvSD/37ksEGSU8fwVwtVyYdtEarPJ8vI8xduBP8pBTYapvI2JcPnf06i3TRA1u+xs
1/RpaQFCQmJ6TV2LfqRV4wvtiYtyLo37ncX7/eRi4iY+FE3x6UgqfzFkbNpfNQUsWY29ykGYgem5
EtPbicw9Gxi/asQJ3azaguqVaq9LYkTl+qS2/8Z6Esx4Ef/wgeak2JAETiBOVYetwLYMLV5u2nNL
ZWqYmPynyM/tPyArs+GftYqPCDemHdBcUDYVz+Xqluevp7S7fZUOytV/Labe2FWnlOeQXjXrTBGH
sDlTTOc+uGVVkibpGOOFEE+RjwMEu0m2bzown+TFa6OHdV38ObeVYaGrBO9kg7wZaItCoIupyPH6
Ms5XqNcmraTCdZbBr4tDXj1ANwWECmaCNMEFmQ3kaev+QFtFkhKzCt9Zbo2CgEyPKzUQFH4BEIPa
gnTIXrgthR35amgZwhk7QLev9sKuwADjJqfiJg9y3DI5Xa0ym1P5bl5b+LAAygQmZnWEPtK62FBR
IypWN3l/WlaBhLfzpKF+/S1Rm2lmyC2YFvbyC+jKC23Qwarc2TyA+qmK5lf/2VeuyVu8DdplWzmd
pFwTzKxCk1xSWdLK0/fzlisCsQVy6mn6Faba/F0tF3t2g6bWV2RNj6aLlyIW2xoon8238xIo2M2k
1is+W0ZskQ0oqaHpRqx42LqHOgbwM/BvJWBXvU7SHboLr2hhgpEQLYIKNur93+H/Nid/XrUCRTpM
EQ9ttUfBGrvhYR7xmwbKKTxsVV1mRSxfN5OyrZ3j4Aye+6ufb8ScuZsl8j/jsMyHWDl/lDLHRwcn
MLHMItroV8nQaqoHXRlLvX9r0imlsfaU+6OTP2uL0uE5jWp0usS3mXG+7e7SvfRd6Eql31bkFpT9
4d9WLt2lBkUWIa7ajIgHnoyls5ufnlg0gLsMhUp8ccMJaO1+PP1nbbFJMBNbclcMjxJW4gJ9U3nm
TtEE0j0FeeIh+p1dbYAGFhSjPGd5aPq41/mykIzGwv2g7pweI2liO/+TWpTGz64ikBA+H0fNYspT
reZV56BRmdjRzZyDUMViSxOaVTWQP4bGa4x0j5ZFeD2wsxVsPyG0YyxRPsw/fhMrEITtjWm54YbU
HKm9HYLwP4M6AD0bolO5RpdaKHWKdOf69vuRQ0eTWh367VncbcXf0/6GbqH3K6qHbZXMY13Sk5Y0
UikzpfPzzf2lvHvefl2cOuATXRlxp6eDXPCsuibgIFXarboPox+Dtec8e51uwvZpA/Xsm5F+x/A5
H34+N2yKV1SMJVfuIEA7mlNnixaFz+hJxLnxr2Felp3Qt11y3cH4twCZakjc+5RG+a6fcDm7RWuN
ipayzA+rXMQyD9A+axMniJ8RnavUauEK0d3V885mRnHgv6Hgu14dr0l4Z9olQlHSqQ3zZg9h71P3
w9Y9bvSxlZsXW4oFJokZ3/eNkbBfMZQEQEpI185brC5wfBC7Dkt6E2wUSvUxjbQrkxU1kEd4x+dX
6rj/FBE7EcRT+c6QZ1hV4gX9gJXRMg6pI3WX4tyVswPRZnz2d5tutmnyc0FEN4DvH5wuurJuvQQC
1odLu+NTuwCEw1FC4xOjww5knn6xCigVPf87C4cbxUYIsGhrJMO2jXtM2Pt37nfcLNATcL0XskA0
h5jFRha+XfCQD+IkssgWNlv8UNXeDCpBL5G9++gsT/PM+cquypMPaxy2+4GT4SpI7cv7kBr48fDa
2Xhwklp2tEySk0t4llOmFkGrrSlJmJSxJdTEyTqFLNl6IXel2InQRthlEP+xrAJxG7KyMUiSTcCg
ITBOYZTpQyKq5BGYe7DlO9g18iJTdis8ulYfb4EhK1BgLsiZtUn4d0c0IBX0+gQ/UHghzeqNG2/P
dujeho2UVM717i0Q9fH0cODPZ0Nz8NwW7ID2jSQD+K3QBBZGgiGRunzOtSFkTwsn7Tw6lJkGmlUw
8RX5q2HHflHwYVITSNhOEI2dcPdg93dPJOgIsToN2AWSvc5bZyTa9FEfTo6RUVD7a+NcmxcE3sFV
6q+XPO2mXsTpN/z4n1UdonZLleNGe+Ku1M6Tqv8G/DVTEpotx20OVT6R4AarKooDd10dwuS/vmIL
mg2OJQqv5Ih9IBQlJ7ZyBPAKzR/Q7wFp0/fItyyjoU8M2U746o4ksF3fwn9aM0WPYOsT0Ovwkabp
tTv6zrr6/1dX6cQgfRrj3mabBe7fFw/BZ6sCJNNAAiETK3vh1zuxQRU0m/qZwH1x60xOzJ2fg4Ck
NO2h9l6TMR5Lv6dQnVzgXx41ZfBwqeySMD25vOpkbJIr8T8SjhB1k5r5T0tqLCIk1sQ3b0RxANiN
cd5i1b/fyMh84ZpJBFxVVJHLuuCa93+xVOPdYCmW2Vqyx5mhPCTzvyZ0Nk6v0EXCxnbeaOxMSnks
OWDik0AqzD7Z82z/mrICZRdODcGpxMUBgq8rPeYabJWIg5Ubja4uKErJKhO4HKD+R8a/HyOLQh55
c3g2zu4jrzf21qdTEFOjoLSsW7eyIDNLyTs9bbEtw5SLVMU3AzzcYQIjleiUF3wZVy4OZ2bnY5Ln
h5Vw8q6e1xPCCJYcr+AC/CQ1H7Dp5QrGlrrYF8dJ5cfx7Fa5qQJyGX0QO8WmGzNdFxBiK/cx5SVG
RQK4md/IgMhbRxfcY7/229DpWn3iDqA17VIxAljV6gDdJz7/mtOpLTg8grQNoNP0Pg354VSFh+on
3WVJCIWs+2285Cydwy/fqTZC4SppUWCCUxXR1KwEvjT7PfiaZZBVGpUY1VJiWU3Mu7rht7c7gDuU
Jq5ErMKjLsP5GtGBSZhciowWzmqZZHeIdGId3Dq1cZY41twT78QM3UI7u5ay0cNH0h9n8tY0QgvF
+ofCxCgvqzWjzHIEZUiZpDTN6Cfd/o9ygWyNnBHYbOgyyHWwUMSXKiVjmvbn/E5UITYEQppCet98
Hld2kOuqDmCo5CMivtw6iXcBOlx7eMex8SMWWRKCs+Fz1EcLlSGOkxyUdZxJtieNOf8jN4m4fEcY
Yg+L+VmrQ25yuvZK1ZCglJai9tWtIPbDZ9MQhE4DA3bIyp1xHznmctetudtMDleL6Uu3CU/WbsyP
uqSG8oPS2kPHlRTWrWDwKaUcf+iFSi5GxopbXaacFApRnL9qDiz9HfMpL4Zk8x55wRmS0gax6rJ8
J2Ee8rQKLRTTXPS4TEb4cJvBk5MVC4H9ynVZl8sbSEN3egPmUDvEaVrkrSgodal2tpNaWm8X7iB1
sZ3ZxQlDxw4qiFxSfutH+0iZGVAHiZ2pyzmineHHunyhI2HrrIdepM+mtXXDYWWDosIRXoYkIzcf
WUxGs4msWIkOJJxnV78f1//gKC6SW+mlIp2DGBOY6KP2Np2Ue9p4C7vckOJ15pSRKbovjX1eLK64
ns0dDbWrWJTyst2/lYxBMXZCR6IzQHjjUiB0rpcIG3gv4duBUd99HYtsXSS9aK8yxlEmXd1q6M8G
O2FI2Xvec7gSECr9SttsifX4PWOhB2uLxabDrxaLF+qZyYi3fAZzJ0oJvlR05F2tHggIX/LdW9NV
qlGXJlJ85hFM6XoJDgwGlSwoeOhC7yY2AzR2b1oDkoh21QzhZPq2vetPhvs+rzde14xvyQMtLX40
Voy2gLj9edTebLPQo8PJo3lBtArOkYuBOot02WaHedc6F3roLrFUSn38ZshFl5MI3mN5OELZvNeR
UQ8eMxMGmdgxBye+qkONqiGrjmk1Wsvjg5d5wZ14SJElw1pLM4jzc82QPSNhwU96xmbv4qEfRMA3
z3iheobMKXzsly2NrAyeUzR6YLbz7ceAefuC9euWjZappr6uZxZtKxk2rcOE7XodaZ91JLnLUlkd
Ur1Du2++/HHPjSAEg4todZ+bYwvl9/h0xiL+BLoPjao5Ddky5pzwxeses8zRhFJagUX9oC2meDEg
DTCIIYuVgg2NW+3tYanJzsUIHU83dKl4/TukW+NN6zzKxytIZ58+cX7TuWFl9o4Gq7DFpHhWhaqE
E+Hd0hZmi4vB5GS74rKQ+MIckr8e9Lu2PwoXf4D2rrg9OTZYGiCln2gT6aRx0yfPyMa7bCKPDqSn
NKmlz9j08CTBUuzjlRx6xohgnpQyBRs4vMR/e0hsKJ5qol927yzZRyB0kUji6rN8k44UKXM7WPIJ
aKIeST0zzpMXQfQEnAKC3GaeJasZDacCkAVMOUSDuab/fzI+KqWO7uwMqhm/QZ7KqRXgyiBaC7Xx
gj+Yd45L0SwlHKgMnxxLINg3yGy+qu4jRBmCWw44uBNtZthYP5dPIlPcdc5oFEnFgaxSOGv95EfE
lTu7Khpo6rMI7J37nkwAftQmqW/+ph0gi2prGb8LeZlkoqtYnYfnsj5OEZSyVVJnNT0WsvzbzH0S
nxZ/TnhqinzW8QMIprnkpGn1uB8oqSUt6Cl158uRj1Sf4d8YkLwwDrn0jhIAo8MvAMIMr4zq3/6U
FmN7pp9mFPZML/FuYtTnNvTE8YKO98+fXZ4oF4QrqZzGdAC5cW08UvJnHQhGS1vy2q8VgSTzG0io
Lj6LvbEmjZnF13rzZMyxDDX7+T0V8MTYRIZub96Fc/b5vGvHoz54awpkzFnzrK86YPjEmowPfaFL
s6U6M36ph31qc8rPcFTZ3BZwUclbp9v9J6m9PQK5bj2KC5EfAkNhkOfE8xtRga6JYzk4cEFQryjy
RU/OJK/8I74/zdeg4BPvBO9o3aGHNeXoXoBUslHj9XdPI0aIi1GkXj0j04h03ywtKDu9ctPDslZZ
+lKcTSiiA6bD4AbxV624ivSW61m9nBi+wvPB8QHDpmLHUPzrnVqWyJdC+0VtBJKB2LzRkWvfWvRy
dbNWmbZxj8H8rBaQXXjVlFrNzrJmTjysFUCRY0AKXzl/vcxzGyeZ/tXK4Is0GvrQs6ghSEilFAS3
fPFGoREkYtmdgaouojDdkU+ZF5NcsxVALUix4uCIv2NQwPhuSk7r5a/hi4efl9232JScGPlCOk90
Kg3DMmHbKYASDGUYpL17Ie8pxxy8Bin5OpKL/UiQEfcpQqxhyCBg6J0IHoH5ZNM+3Y1g73I0XuT9
XQ9gLGXRyUsXASewbD66RWGCHF0yezZ9bBvzNT6PopqB0QNdYOuB4typQiNzLCmoD1yrREM9wS3Q
qJA+Y3ZKn8vWl54YK/gGHT11Lz5dFugGFvkPuSmw/k2BNnXsB9nD8ZF4oLT4G0YqFYEyOigTIko/
l8C370vIATpJ1wh/AQS6OnLANaJcqfwW7ctyz2St8wHKv28b17KNYgz6YdBw3rTc7dCCEkGUxwj+
pqOjPaV/k/wfo1OeAbLi2GlPfB4ifhqYVFf7x0WcwCu09kNPxdrFHwJlemRUJvz1QsiVkZIlE+04
sVoIGCzeQFBzphlSc1VBJ7XaeRfy9xa+mHJqsjlnC+eyBm9vBpiq3ryaJxYRw1RbpB5aezAO9Xcl
ITdddruQvkAFD5hx8cNy5VZ4MqgEdQooLC6q18BfbgY7CHXzM0oz6Mt0k8vZl/Tj98X1oS9oaQJi
5GN8MDYoKpaVwiJn/SiZrVe5jRxUSTjhNGkDqKO9I0GkRBdXn7M2HOx10AHlFJDzEopWoyCsF+kC
Itm3JZzeRGqphvyU8nWF9kEPwi3GK8elpw2jBi1gSynLYc0GDC+0D+rIZcypyCk+KxqF+mftcWRd
FDcDMBnw4L3t54EUcbXFwljASS9BrmZ0h0qOdtCsQ6r0z5G5vo8qbaRWz8svPux+r23DlM3SrS+w
E5T2fNgOZfl8ipUFO3GCB/BW5rPoWv1LytGx/LyQ11RdZ/ABOwnbBo+Q5bzbUParma9A1ttiUtwZ
nGUAH2RPhmFJxtZlk/r9bmLbaR2r8iing24ulPdTJUYtMD5sj75Sw64VqI+9VtSBdi5IstwRm+jE
H8COYKhBJFnf1ZjGqKI7xbR+yGY5vkVC4nDKODNGfGMCP1RlSSghVsscfk+0VqbARAWJ/zgY3ocl
YeIHBaI7NKS703OJb206jdwBz56XckBZ0NUhcZKjAvoz14YqWNF06Dx6KrAbbDbhQ6BMxILOH5rE
yFzS4HVIYQYUqIqF0NxVUOABRg7ay4jsQ31DF778/UiBietwIuOOAQ3/LHFEK+aAakEazr63cmDD
ovL/r6MlBJSZj5vOl2of2cHrHEl3HF96I9BWOIfg1sWMeGwby4rUKoW8UrTWpNdNb00YECEL5ohO
hJpZTQVVf5L09xcLGTB87Cy4Dy2ILEemNha2JJ47ouLlOO9J6D8SVkEsw6M5nbQwqkg6RNJLVbZ/
UqQ6xyCC2DXpeeOjYLE3Jb5GMMNKQaXnPT2dRD+t+FD9DcbcukDoAlzUUg4gHhuK1239DLCCBUL4
a3Td1nCthMuY9VweH9nTsXolSflM4TlME9wprfLugQ2YN/hr1jIHjS4UiKB+y/1+cdCQsQEaC/Zb
vhFHxflbGqqDFt1Sc8bu6fl0ftlv725+u/Rwx1Y5+/SRn6rZ13htOBAVX1/YXq61ZzH1ya8+NaEm
/W/ZZ/eoiOqdUTp/4matvVd3SiHCa9XzHInQ87FN+esRGuDrwRlqEP2RWPxLALqySjlbGvTMd2qz
epC3DXYcITQ3qOz3dOfcyYQ4xhIlXqPhYHtw70mpdseSL6iiF9KYymX26EjORFdBhSXhiy2cx8X6
NBgb/NKQ3DLkoSc5Ar+pmMYkv8rW0tQpT+1wae1BqGyjpi+0g3vka7xpq81VBWYTUmzORdm8UXhK
n/Nsqe9aVg6Wa0fLtQs8NLJg4mFoB13jgP4Zo8yTf5HeA76N0xgMpi0MZ54SCNzUlV3qA3Y4TIJO
yHUQB32HHy01YwSwPHOwoL+xiQtM2ewG61VSv2wvU0h8OLRI4ci3UOX6VUchQJsY8lFkjwlJPaLZ
TQPoh8Q68LTcsU7bmb5gXln50+iulMfSIbglvspqAjcUASeA4SCB3OYnRAtzrdU6ZWSE30gV2x/2
+4FIsz83AxreN/oHcKBzWkRSpms+1p4IgCwOExk1+s2T1RRauaO7/05/UpRPIImmpr3aCtPAhUbW
qiCB1Ik4+lCOTx5q4Ii+pgULKKgfJ765YpfNqn87Lu+WqFEE25STIvX5Aci3GDLFjhk37lZJ9XRk
Vrv3rNn3Lv4HijYC8ExSq1Mx/uV4qji01+EFxOlOhDAHG20E6jYaRpyv/bLAdHh9+F6g/zW0F0pr
oXUsT8YGe88nvGyf/fOmVb/ZKyxpBo3oawi7Vyo0mfOxmyRK88oc1kAtAAgoAiIcaWys1+ypSxw0
wpxqjAN0AC3eJXW3P7NZq4lvOX1CjIU/Asqux5sOlhX+Vjsww2+jRY6HE8Qv45Ap7rQaO5YEiHYs
vlZjiGWUXkm/3wV7TXEqe5f5a8Pgq6PQSiy5R8AvWtbvEEqiWd5XjKmyxg883gGsdMxAsijLI/Vl
vdtPiC97O38EBBksxTECzlAk4eEHZRH4dSEuezwQ3Sg4BOKJY5EcvTeA/5X/LNlMNXuGdXy1FhWA
VxD+Ew0j5iIVEiFVw1W6nryKIsZ0s0APLsHZPdbAtkmF1gBzDuBVMP2Tle1iIeNy1LrqpyFrE4iO
IjTBG8ZvHHu2h/uKImW1ymRl8TAhPCGTpAAVMsY+4eu0lFiuEIC73+vkEQNweO3PiwjMQ1NBkSQA
cczPPcO0AJnKdpNXyfYgz637m0pXJMiQVQXnSla8lzWFbrk5u30MbSBpqAdHEeZCxrPfFmQuSGXN
5CMMfMS3e7ChSEXgawwBpxPgQfYn/HG2IICtDmW7d2HFWePmYdgJV88Xi9mKSOrR8kT3XhyTbhTw
UWE3uL5rdZ7gwmehR2OMEZNHavtqhGXeCoBgaCLIVLzCYWfeXbQ8NngAz/fZCg/gNvhqfwXPg8KM
CEI6CcrNu2yUMwtaPpvbzIG/UZ9k0coQwmVFiEgSh6wGUiy15Ibn3zyNCs7qkRnS4xPufYjwucGG
LkcwNS+A3JyNJf9cq/Thgq9WOSwulHZ0h/dbxDs8XiPkPWSbL/kI09vPOGwe9KEcDofhX5I2Q9n1
lbhP9A8qmxbpYblsFUXe4izuHmqDeQu/3SU5ZLNDU+eA7AA2zfGu5m0Ia+Dj+b+rImnD7ipRpWNW
1X7WJtsfqw9gsyeHMmbRXZPOAi3MJHuW1l9zWJUZqXbkY59uf9xXdO2/r9ch8o8flWu3atNPt5WC
R4lwoXzVAyP3rbdPLlHP+K1N49GMC3trkp6dlAuMNjs9QmnoLyvvEEBqHJIFEMGC8E2bspDVQADD
SkgA1G52b5y0iFzRbBMpC9FfeWv99UJvlQWwZE5ng4j4PaaIH9Oz7sgyGBIPn64dRMHZ8vvqvcqR
jEwZt+w5R0y6l0ayszl4bgDJI/810c8k6e7C8X91hfg8GAGK2PP3T/hSv8ieGzuhBbwDqgFVSCn4
Fb06a10Cd0VUsnR7bAmCiX1yPxGwBt79YXrtrJ0uJlZs8HDo/zDyjhT8kIESQ7hx8IBuOpODYfsC
uVTjgmY7jF7HbxFo7wgw81J2hfbGezYhv1hMTImwcICIDumOfTpn9bsRw+mniVk264SWMO0Npgyc
u9dO/30CRSq39IHlKb2qh1G7ot+X9Ox0bKl9Dszue5rD63ZT4wlWob9RiaZouExFUIKOu87ExCHG
b+DyNALoGl7R1DFSSDWvcFXyRQB31lLvSrhqdQrFcPh25ejCTGHcntCdvqhP+VgzdA3GXcSDpdDV
eH7PZ1/bZ/WmFY9pbBlXM800mrWS3dMAj4DrfOZw7sOU5TpadFrql6jSnhBiwoxgkzuVrMHJsJOb
oG+/VXQ9qyejCV8kBGuv6+hx8DsTtGZjPRL39O+3ecNW+XosxzAofY8BDGKTFExnOvsqikVwK+Fx
upsBOaSEct+/oiZFnWv3AVTBMaGD5ksuRjt8TvUbqwgjT+Yxli+g1p2k4qxEiaSJlIXR/OlmpO1q
3TDO5RP4zzoYaYXQr662wJ6jmspfcfypl44CW2f0X12zYfUhXec0jTh+RPpln+e78Zuhxa+pLBJG
ZvWzSe40EtRxfVFoELwnkZjobMVQ7hffWO2VWEMcwTxShdsueh0H21hCoqHsmbEYTU/CO6UC506e
n3AtP/lBDCOtmhrDtjDy5YvKZAS2hcpxpEwV0r07sgvJuyPCu5e9Ib2lP8TAfpWYFVVqnuBENqzB
z95KNpl/vXpvc6G2G5cWeHPRukdsPJCXUsdNO14f+rUFuh6t+8USZ6HwJ7G8+Yclc9BAvgRTka1m
tTrWRakWFspT1ryGMAjMkuUajcW6K2yIAq+uZqEqGbP652Wal1RsY/MeoJURxUQMoinCY6c0g6SF
l7B/Qy6N4MR5YTlhvSNPqwJrD5sSqUjEps7IXZadgoShHQRyfFznWVjWznlAdyvjuGsVhDlQL4BQ
oPQL1Jlem1IWEcN9X73fRBlVJCr72pW4kI/DaYHKJ5s0d2xGaTdMf3BBHqH0X2SEbdLMbha9uaFO
mE0wjsLe5FBDVIAvseMCAxNmWcAx4kjCqG693gv0QqqrRuheW6s/OI5hFm8EGKto7meFLdcPB6Ph
qLs1rbQ6IJw+Kk6RT61rAmMhiZEhgbCwnEI5PzKOl48fJU/ymj6zAWhALJf1x+DVspMNV9T+krZy
uIM4z2UenEJgwxLbZLcz042RDHuCRK1NnZ/jhLn7u5WY3KSAwt2Ea3j0T0LZrgsBEO8xDjA7McXb
mdvRoF5ZDAAmpHolxWEQnccDoIlnu+/vBNRZLCchftTDRmkfNZfN1laPX/Llzc6yvjNnUePtiPnL
YehQGB7gme4DcX12Yq0P4RGNxvit1q5zj3fwc/GmWFtqw1dSZUYy2zzNIu0dfIZtLvdeKp0rHuSo
PX77ZMeHr0pp8AZNJnruMi7Qya+XLu9ADzbTIB9dTdXsM1Xmge6sUhAz0h1Fl6yallwxP7FLEz35
TacTW9Nk3cL6x3OkyGmnXuoan5l7FSNNE92K6/74Ux9srdq/Kld8jXyGRtxA5GBNXnTGcR9ddgU8
j1iLRIrVmMtOUkOOtEbKhX3inHz9jBuZa5FxX2lr8F4nTSwwE3SJuj8E53pWIEfPe9/fECWe+Blr
MhJRCA2niHGgL2iYrAJXfijAFirxPW6XCU2mtjmzHGY3fpsLvvteA1i6FYGa8+6iJgwudnDx0IMZ
ilkNXlMYJIKM3MokM344d14gLykJ5D2uvIjEySrYpVhxWybDfqdp7cG3i8dFw6P/s5RVANTaPafi
THj1iEjWTj3EfQdOFU1kBWo0L+5jEK6j6DY1ubPXWIxZWL/uWBFoxB1lJ6aorYt/9XMWfOosO4lw
FL4A08qrfi7w3f9F3SrKeUO4NodD1tlR4i09McXShShnrBGQ0eLuuFQDUL5Oq240Vqm4cimiNMa8
8gMqKr1cv6FJ20I8n2CovS+lFUk8UkiWegZFI3/QFfZolnsCm+KM0RDTaYzLRRqmW9J307rccKbX
nXsXZkmDkEetvyvwrKjc9EkMbGVZqLbWz/kjp+dJR9bueaKDqE6WEJdbyuUVlMkTmPHYOB8G3sOn
QCRO+CafS953uP0h4XUH1JC2LwCUBl3fS+pPHmN29gwJkmlBZ3nltOIPZejqwmVd3nPpn7IK+xO5
XeqPLpouM77FhsJVQgp+HuqcS+MZZdRIB40EH2a+4jSw5gI0a9oDntmk4Oxlqn9WwcPzX2QXsiap
v4x5EZp5QavNx+EhBwTkuCrzqaZdU/wNe8FmdSARBBB0HVKmzeHTQ3gFxSVo7kvRcmigGWnc0RPR
uAQ1i9pgs6ZF3pkqrDwbUc3/jaS0HHdcElfrGVvdBe57Lk1r1LqqlZBDCLb8uujYm2OGwQ1QTwY7
UwC+/2E258ABx3TeqPq9aBZqKPOpg5Am60WnoHeopweT/DnNFw9dzx8DBi10fjiODO10IkSa8RMU
1yBfSs9bZJz9KIfuNZXxCL6TeaLgZb3jh6RpXJ0vtxkH2ZlboJBAP0qQuiuMVfeOUgfH57aWTHhM
MRc6b2BYlsQnzyXXfgxXJcwEQOLiLJTFIPCjm2thhouM/z4gD43SaCn8DwjzHAJRAWBszoJ3488H
QjquSuQ3EJ96fbO0koiaxZv2zYSV5Ehg0CnzZ/FhFnUCTcpC5+4h2P8l5uYrmz2g6mT6/VgT8PEE
fGgOWPtk2/0xi6pCy5KnQb3yfAMfU+Nz0fR96xsj/47Xk11kO+fFVrnjrByDF0BScLkLPzcE3w9G
UUFrneN6X/HXx+mCKN2O0s0bJHbbuM8UpHSVvegXo59DT1eUsUa8dxXuK/vsZF2xXnplYUeLsEot
reNoBqIzrQWF0/fQg7cy194aEQ3Q4/m/Pu7Bpd6N49n/uL+GNtV6dZjXW0vbvSWjc2MqDuYsoCY8
TuD7O2vr3MQLiWkkKF20qfEIOGwQw6ct0Bb18UKtPPmncZ2WxB3g5G3aJjEoRf1xLzZ4IENMdatu
mLxJreJ6hvBV/Q9WcdE/6Z+OopZp1cKeCWngeioWR/rxLMcd0j26jBQ1kpedNUt8eYOug4gLX2bc
iGyruLZtrpWAYY9DuOo7/v6XWO9luq+f/z71svogBnZI9B2PBy9sMtCskltQB57qT9PINOGMRfeV
gV+tSOw++DCeP2Fp6panWlMY5nVbGoe94IVKFJS8JUrp27i/13Yj9LaA9bZ5Cb4ZjB3b5h/MGEz0
dBUENs5Tvf94R7CNPM4Iyq+aZroccmBxoDSV9LT44TJgSBB9lM3XHQQXAloq1Jx4Ql+Lw+t4p/T6
E9ytdstqNtiepzzHkdpzLn57bUxXhr8K02p+0Xg+xQwKl/dp+CV21E9kaxhhvlT4wIUg01zesRP4
Xn2Ua6f2mFk4dV8+zYa5wQE8XNzvDz8DzS98qBlwXbeIy5ogH2uubyZvTv4P3EZ2mR6XGXHut28A
+GmhsKARMLZGpHPRI1Pcmv8aj6xdiJcteY60srC7N0xrFVLTKXzrcgN2kaPpz8dBpWBssaLmTsUG
HHh8h5RWyA/RpVmlOo7Gfcy90a6cQaVuvKX4/qW0yGWEMDfcAMgz71irPVOcchDEXPMEljIcDr1R
d3rRlnounRYMhhsP/UoTlaEbeW+OX8S5tsdfGl/oRMRKzOe1+OMvG7Qvdo22LTzLFde1EW2ubUZM
Smg26h5qka9zhFNZs11I9S/ExG787i5LTB3efRO4dtPFDOwlpJd9ptWjDWOsZ0vxJ/wiYHJ1JnaW
Rrpp4T7cFpG7dkI9C6lYDDUR9O56NEDIPbSiUEF8trjXmQTCEz6yiLuI7ANdpu1NdlJJg+1MfIbc
HRPk0ldyu/zxuUjB0Yc6bGFpfrNrRVC0sWmCdxrazc8AtjknhjnY/t2ChfzajhiywiggTUL2hNUl
ThlYF+aLE7ZDzF0dqI0cCUyQfDHU6yKPb7mRN144LdXO56K8FwbVygwd2PHqquVEXmiTltaY6p5m
SU92cJqQPaFlt3k5YpyxfG1Nv6jLFukTIlZ8wdGKjC6eR3JQ/qZgkBzPYQXF1vxG/02EFIE/1eQW
DfKWZPpKDfoveX3Os7AHZ9v2HqEqTCJ/zCEjmC2QFhv8XGb6KcsYLzAThMdcqNXVBboyLWc9qd7D
vhB6iEqRSVdDTl5zVEAIubfFVZg0GbiZ1JBbUksVwv4TEFQX0yzcv9LvOhLJuPcMNm/UxFw9CYM0
63zVycMZ/vqDWiDoWQjcRy9o8GXwgqlU+pzxQyBbVbPGRr/zSM0708WUiEe8c2xNv8oni/TxLUun
STaQH1PSro/nqgYKVM488/t75wTqWU4fh1ZAjVTLU2kTrO9qPrMuTLgj8F6YdxUgrLm7p1r5FPof
kqCRvJ5Z4pd+d9KfZY19dn5jXZmqtbOz5Rwc9x0PZn4aTTheaX62w2lMEs7LH+BRDARKm1yyUae5
mxrqB+slCpi3oJRklItiH3KDP20HQYwEC6aLOyv2JOViVRfFyMicO9KIasLUw9BZ39nwyUtS4ywr
wN/E+nRB4PnU7WCRHqvZ8fjq5+nzZ/a4idE0xh0LhVASa0nSRidnanE4nPVjbJtjBbtvTsbAlyjj
qI1UGmsLQpr6z0DCK6epqbnltck45aioAyRh7WagUroTKzfI3FXdMNgE7dpiberMY4jD5SAktiK0
ivZNCSp6kBrNbut0MNvpi4B7erI04OUxUnUwW+CQkgj7azd3k0+4pGGSrg8g1xeDQYvfsgVyPC8x
mRfG6kH9+Ufj+nV1HRhmKkQZs9Mze7lid4akBRqCJpHmP3r1sCBjnvu3u/TelpHvtG4+ZQLuSqd4
xwJc0mfDT4Xix4ONUGg9jl5ZNbElQxhwwsk5c/bqY+EQ8C1R5RxM4J3fS5u2Elat2onnAk42S3hu
WAJrCxzSHr8ZA/ucUmefHbT48Xrp75ckV5jHBUBhLDFV68NsrJOIQjSp5BaASiwXc9xxpq8/KNcR
st1EZdd44+veUXMcB9N19eMiGakfEavD2rAr0QJo+yQOpjnD+HfYAvYsCzCcozo1+L/Uq5ks/ZKe
e/QpdDYaCMOZENO5OV9y0jAbvuyRCfDIXCaOQyv77X00RS/5USf3ceA1buYYrk8GascM3wQri6Ix
tv1v2UDvr8pJiFeFrVLP2iOdyjXOQzjx16ctPkXmXFIHpE09KBtpblg9Bf7TG4MYXuGxcBNeFPV2
rvR9tdqjJCEqOb1he4+c19upvE43lYPhkqaig2SmdWRvyqdQbGC/FjNmrY3BngtVd42SWCcA+hTt
utEGQms1jeIYbQ+Uxl0yLiNgvFuERYPk11f3jlhXt338QpIFgB2GS+iptLqvm0848BJErhTQsaLu
0Alh2tDwdugAoYhogfnCDK4TeCQYzucl6FUVeJY6r7nPqNqsC30gu5pJLjBuB2GHEsJ5doPZBYrV
T6PDSXV/80upaAJua6feuVY1Xv+DGK4FdhvHaRdvaHlVub0q0Oj+mrj1SL4+JRDYFx4Uc29eE8pN
0V12i7rC0LbXasVwLLwx+dWndjYvO9QkHTsHV6uJMQg2QIvDab/7TASJKM4890d6EoI8iPppnMCl
6vHiKH96S2+PwvdfxSJKVS+2yEeK0gkICxZtN957MbxIHr/6JVKVrwHCoVzOBhfX7xnS9YNqAzU0
eM+QZmHao9nio/djFg2jVF8EtlB242qB44CzXX9vl0quK688F9oNfCnet0ub7QNukqPw8/QTfMOW
Ek31O+JQ7x5MLOxGxc/NgDTJ9YOS9ZlnuHlMZgnlf8rMuo6KxGvyqbp3JWiP9as//113DcdLk8cW
UEQsHcP1e+3O4QXHvUX1p5KnWo9JlVSDUELWp3xD/WODTKGANOOiu8BIvereqt80tbBLqLNqgt0p
bzCVcng/j6Ikwl9KXvNW7RvPFSPvgRQoOI47iZhoGvGXpljjUChnw33PbzlcG2c0PpJl7cYKqNRD
E1UiAcEJWLjbwdFFQ8TwKpLjE4All5KFFgj0jTIYad1AbChzdDZZMwdHb4e0nqNgsgiP5eAq7fSU
CnD2890I7ta2As8aMUuoULmrjDwWaTzSyh+Zsu0J/0rFS/w+bmnxAj8IBNG7yhnKEsCiyunbBZOf
TR0W2G1IyXq3UvkJVM7MAA5k8jGE2l0A4cLlNhFllombk7q0hLnbkAl/vPTKVwXxmzbrYjuWvH24
XojYhsMJSbPV4Jt2NjFpZyvvBpEm4ULZkdPyfVG9gFca03f6Q9ndA08qMvNUU5NQs60X6LQJw/GQ
Dj3ix+o4Z36afdVFv1ZoS1tBhpC4W8hMEFLqsJpRpT4q3gSAqIAStc6WujhA0+w8YPuf7/w99xuc
8phlFFNilJWKpp8eon1c2T6J1vYg2T+gd5AjNa6JDAHJAzuHOq+6Zz5R5uRkd2l/Q8RuBVBEVIi7
2uYDEY3JL/xxM+Dwu5ArMFA0nTL0p6j0CgcfoREfJ47AQO7vR0N2J5r2bq6uEct6f2iA9FOYtxtS
Dl5gtVf7UaAM+nf4LtRiQIA73pgeSA0vpp7m56bWdU/RHc9l3Nie2KacmZ26X6w2RlCKOaB1AWgS
HlIjxNgk23yN93Y5WnBpjJDIXUWAoHGORHtyL6ORjchT+fPaIXM4Pb6FJl4w/smzf/Qq85q0lwo4
i6Rr6f73pB7me22uytmYxMw476jzWI83ZcWyzONDpaqAAF5P3+DTH60eIAYXL4I9ELZgIt+Cx7zg
sSELWig4Q4engKpJ2BThEaAGCjVCTHUTNDIoB9na7jUy1jV4nJXkhGzHSppeuAwXntkPJc8IlTf0
Xzx4ZfnAec5A+OMVk/F9V2AqKgrM9ZK9rf8MDDCJbWe+vfLfcYq+iZDt4oRgUx9LE2FiiuH6x7P2
9TUH28SELeZ6FKiAJGqr2Q2Upl/dm/hZqgbQsAc584gPebN9pMc2sY4zri627rS1BO6ksXSQ7Jkg
/wf9g7M8+V8dLrtXqRruS/B4M/8CKKihiium50Sr8IBkNEC1VfSwkkEomC758oSI8Jo7S4QhYtEn
Y11rkCsVM/cSxKD7AjjCWi6o8ksnGP/LZ6dGGJHl4OU2fM93L3IDOt/e7BBuXCf/HRyNX5yKFVsE
VoIgVhRhL1+rfxsAFKbQwhU2xOVINhXsMyvmdLPW3jceLUKqlw0w3qPgqG7eJLek9HEvuqJPSGAN
6uAcfwA2YQ9CfZCV6dtgfQHas78GoLWQcF5ylkV0RFh9b6CNbHbKfHRQDb1WHP9x3NNl5pdCeNFM
EdZp/Iz8M7ndrRoDbZ52aNz9BQuHmJW5+gOkCifFyI3pz8bVqCH8WZwrzYLT9Fsq0KVhl375aaPp
MsAk1DsfQp8DQZC9EpsOdPfXaGa49PYDTNm1yY9lOVPY2hZvxlsiMTC31dMrGibBhWJ/+umuxdb3
Xxeime5ShaLK+h8ZIDFbTW/OR6BxvBSP/dqFpyonXDByhrVcbN9JpGWOVLL4UGPcpsD9+CaeQAKC
7BjwmAWgBECpM0TW5RytUiENysd5mQ1fyBSg5hKeK1W5MvFo+3elYRvcf7V2QHrdcAgBMPfLKh6Y
AFz+BqVoeE6onIkgdqk1bDbXREj5PZk8P9Owxmu9jOd+mQ3HnGy0SdJZGuSsX/FHSdaDDDdpTYpj
Abz5XpPXOjIlORr8tjwuTzxCN8PeV8afg2oukGlYl9RHGVLHfqK1ebdx+GmjEICos530rwpS77aM
gwA+KiXk1it1B2pv7R8E/PiGpxWPw4H6vvXo8iy2BFGKJGHh2FSJO9PEcS2IIgv1b6X4jXLUaEa9
IYPawEDs+WyeRx0TMUBJcXDcuMavWHTRSKrW3SjvE7BAuAWpBkZaKAdcnuzvM3PyRKVIwDtGJ0xk
JnpQhEh1LrUFiE951LZtqItXhUnbiG6s8yJXUIC9Bd7smUzk5SA3IzQwSXYpsfI/lVR9JzTDG8eo
k5HIuFThZJclfJKFF9k4WVa8V9BgtC2+95kQ83JdF5da7g7bo/Q8rHOrMH64eURp7vOL2WvldeVq
h5r5jYKx9KqzLZhu1gd1pXoycUGkrMEGJmOEAwAIKTfsjNN2P9pfQd4CRpQsBv9hVQa8GA078Gy+
tErys80Wtn5vRRcGAe06bztUbhY1PAX+8HB04UzIHQHttNDZSJJQuMGvFLUFnzhHjIpf4yORy/+J
/G2KxE1tPIU1ZhuFJImmP3l7hUiClXW9AQQN5oennaWSKKETyeRgZDYQjBs8czuBn9Kud1iyx0U7
f27geg5ZkWRWWx/q9SWr63WCtpiyQ2/N5bOR3JfXGaN9Bk8O50OP7/xoV1yF5pfgT7EsEcN+eSL5
qjY5KVOT/odRwIlaJ+uILRb0XfPVq0YySGkHyNo79jsBoMIL1lhuHQ4cg8oG+tCFTCZEkGJz4/1A
Hb/48eyp741i+GGfbhPLlL8m6fL4rL41PduCQR2QXMJpkLr4Hco3Hh3jGPnrcgYin9ewElXr6gUF
w+dJTkLReo7J2ulIGYqWGfViD6e3h4/bBqBz1ZxO/DeTunZy5CO1qV48xzLFrWHSqSfLA+qFbDqo
Nxxb1Qk7rZgfSr5cxEgPzXnCdt2rLvAUq4rDOQIrnloW3XTh9Vjhq/q7VFAgwNRqTf8iXnlvINo+
e3r6jM/Y+VadlczFiwV5aRoWyDLaNvhVAEHa5tlbClSkjZBtd1nJdLgmR8QDt26lJouhKynKEce0
LwHDMeQJdFJFCaM7V5DWY6XHJBuAKHVuYkfDsfo6inG/Ikf48xUCUY2A42frYG8oCu4BFLeGUg3G
Hf4C+G5fwAuX4xQR6wesWnflPLkqN9N4vy9MvP1OtC+X/FKz6wa2vsdkJDoPmq0E6Wwk9KVAdk+G
SUFXBtx1OYpvVRaa2Z/hXW8cfZEIFtznZL6OwNLyAvOT+niYv5VobM6+6e4wcjoEekcRebc0GuR0
VzUTMB4RHZ9v3r382LbzSD1JtFtHs6M5bmEzeVzNKFMNRkI7mqU+4wkFlXaOlrYFBhePTc/Hi73+
FcTYRyEG62w0lT/YXSPBJ2qNIN5Wj0qTYFozwxBG/GzBWjpqfFjtMzZZbnX9i4rQ09fDN62u2Cyi
ZMAs8WHbJ/i2BOLT3YoJLKOMto3v0N25tkxx1OZqisbNW+GbFO/KViChojFYbF433macDRr3zn4z
ClXXxxQv5jcFM8ef4x5aIBLaJeqXfZUpg6E0NJn7IcKaJkdnMoliNRDlu6mKoxkDusdk7xhDKNQX
H2KD80HlgKl6WLFK/g9GdAsg5eTJAwBYukeF0ZanNJGTK7ibFuCe+hBDYKCQ+Y7pJO839ES7lQTH
Notfx18SvHqiMlth9PBEy1UCyKeIomgIGNKIZQI1ldr1/ffi6nJr1qjYM0jE0UtYFQIFZqhIK8tk
Um+OPwZl6/BYFC6jz73v/SLh3mS5WLGowmVcpGcrc2ID3GU18GPzn37SAYIgovLiS5BPcL/BzFFR
Qi/ddfvoqYbgtj5ghHj1M1/9tnBfiQUJs46L9zpryAML+sDugNY5EOkYVPJa9u5uIOVGnnWhUdI3
QDW8ihToVsJuGp0BAJoanLtdb5oFK5iDm4SvlL55tCtiBNUsL15oqO7sEG7O2I67lOmU3puvuBdR
AiiRynJoXxLrfj0cbIsrDlbLVg8dHbhf2H3WHUPvfe4yfqozXCxyPj8EMfIxDXLwfqkLXQzvtMxh
6MTYcSbQC5EZ/mbbzxBTbnUmEQHP6tVgUuhaSIZzYHmrsG+bdrSGSRRb2EP7mTSexjnmYXNgc1Mk
ARTPl2FluJbj8q463xRyaAe/rjmeZiinNVtKouSpzA/C/JPpXhmFrMio87v2KtkBdUeCpqGysr/K
t73YEgXOzSl2wZ5WlRYDdv0QHpBPwAfIuJifqJucyFCrxPJupIJzIlGhxqv/+8tEhC9tz3Yu9II6
UE9xJEWY7+LnpKd60rphHtM18EkOemsFuQ6vo4fKpXFcOf1NK+rIflukDkXA7rErxMJci3b/iLKh
IkknnQkOrXlnW897HLyKAi6mn4aMAnmFDi8rNik1Hxbn7OLTYBg+8MDTx1fgAEw7jpaH4qYPLq0h
n4wQbgQPJnmLKrrlrYotHlOxFgNz0SNn6IDxzHg/h5sEmsdIJGSBBCwoRNY5RHdEcPBean1dPfH5
fu1jjKbfXZoymPWIyItqH9IfM5UPUPojatTk27kSC0z8rrXUNPHJKBAUaPFQHU7xSssejIXfZ44i
HCDBTKzhGCQwOyuI099i1vh3j2zI5vYNu9zUqeNSX0QhWaE0CDyqk2W1uBRDaS9Kr1yrXle/7v27
3cSlCyRT9W51nDJMGF+jFIFc8hMRm466Xcl8VAPw3jUSfQFH3awNxaQn85AmRkLg9wuMfu7oBWgF
E8zAbKm8RBVL90nGVF+YlvLWxj4p6BG5qOiv9pD3dyLyZMflzTNQC+MMMOW8bbSupRurIvswBKrn
299qvSm/MKHM9O1Saajm/kIlxWhKme4w/bxUHF44f1O0aITQdKVi66QZAhpiGVCwvf+G8RjnLXOc
9dSDiY3jlvW3oo0yvyAuc7ssw6dcDmjrMAHypiLn2NekhJVjt4adYOdfkQcchelN+ZN7angyhR0k
+UXcXRmiK5m4rKqf7qgDn1ubwvvgqpOiIoyd8WS/SYyfbldBvj7WHEx05WFXrssqKM1YWIwpuzr8
f+RSuI459JJaHd4vgykYtcQQJD6plCzcYDFLoYzpZyclpcUZvDWdYvTIP+RsiiU4NysiDfYPLGsq
Vzd67ciNN5FM49m/kM9dgGtXi7ZXc0s2N7iMkKGMATey66946IXtCPWz1pY1M/zf+AS86QdxEPj3
tAUZXmDftXZ2U3RBtt7xPGzccAdT9fwKWAI4fuDbCqLs7MNEBe0sPpAY0bMp5Gz5Wap7d/i+nJhN
3WdHL1eXCNnI6rP7TbeK+GYyBdY6F6bYyfV1dZqsvijU9sPPcjHi2eylcSiGRBTsjeF7axrz4X8N
yTJ9FVheu/QXA4QBHw9YX1aqDKDPviAxiXSGJwKqoNtRbiF1RicOeyG1AR8xVgtElvmpQgN9WJX3
KT7UpDeZk6Z7nW+Oswh2TzFpXhXf+jC2I2F+GDyFH+kgZuhqDkA/MIK0aCJlSrIzF6OeLZ7yJwZ7
1VVEzRcsvlvXw2a6w4pKjgIEbFKct7uxQKkiuLud/KYvmnruj6Nd3/tcWGEImINpyX8FDyLIWVCv
u1SxXwiB7eTv1BgTWym8/LMnEec//EMNbsKg8MPf0D/dimBhk83NmInnFrx+VTZ/g2jkUEc47Luo
XRP/qFLoWp79mkDQ4MckqrKmh3zCQ7X2GDYbEDikMagF0xadSBvF4peGaFS3DA5E5Ebjj/mRIFSg
5GKU0Ogv4cd13SMtKY5mxgQYB+bPY9V9H//mzeimBlp0ijlM2QPGQAOvNluTgZfm5EOma9mQp3M+
i/s07P+a6LM9lGA4lF7hg8tZ9ffDZC4Vg44ExW7lmKy4XsGi4Vbbz/GSYkVT0ePLgGxbEvjryhFr
oFPIuRqtWO1VAGNP8sXswkf8SnffGBepqMEN6clrSTeuVrfYix965+C8yt6uodjDMGcnSYCwe+Q7
qKYAOPCZYv1a9jsuTqTj480jZc+incnYEoJ1uHmnV1UxQ0kZcIwMxiBO/TKHjZY/Fq+tDDJpJ5Gd
QG6GxyAz5XjtWJEhTGzwYc5QVAjtJ8XBS2kbMEsuXxjjhx2PFgqLc+pH6Tk8y5OVLSVPufnCmX57
KUje7Hm+5WN5T0v7TNysysFHHMzH2IjjV8RPcSL6M5P40AyeVlJaw4Lghw2iszRp8GhN4odt8ALZ
ixyf758qEH+n0ZDxhc/FXXlnONqaEX1nHzwr5BzRMoPDdxLZKGAbp5CktgcNc8/a3oBYBkJ03HeQ
q8P+UsvIzxRCGh+9dZBVafnVfGOfWfrp7nHFw2/EHJOi9eSRJgrr9Z+2P7Qab5/hOQoz06nGhcqL
8IhcLrZrIA8nHtjfmulEHZzE59Ej2Zobksq73ahNIQmy/tSn5/R5DoODjyglodrQzTEG1FhKlnXp
z+TPz2mQyVWsHHVTHx1nxBBgxFaWJ1pWLr+sp9ofXd+wj6ngJxMmgIf3JvBPVK59p0dAOpC3u9Gk
K4w+5VK4Z1nchXl3yaZPrmlJ2n5wUwXz4LH2WdOZDGxle95u7bTncJsNw9tlVrF8Sd34t3XazMgX
oFs0HUNFGf7/KxPjzqHFCBqxrZpXmKgrUWt6gs8VFNMFW6A4bplJ6XdplkgW29s01cM8wQ2I94dM
NYvOls1/nPiUGWUp7adHzrbpxI9LK/RHXoAl9BuHA4juWv58+Iw3T26WJFtZ633mVRAcLF32GqrT
mPQcdG204muTH9c/r7VJItTj9TxdhzO19mVEnUFwOwUMs9vjtuv22hdBO88Aa79qmiIrpFyNusxq
fj26p2H7pDqgLLsjGEeAwI/htAgOBrPMpOT7HT9TLrYKyPZdM2GXlg9gPZpSCNs2UFRY7TI5kjrt
G4X3/SFfnbLY4ED+cqRcHUPx2neNYK9j8/I9HJuEDioO/OWnw0jJ/4v+Nmo06y99gMNv7dX7b58z
c30IlJio9YALwWpMvPfDXM/nE6i2Atn4Ge5UAh9VPY147FclvhgpAjkABDjpdkjHqJvpaEs4ahLA
vPwSAHbvVUCIDF/qiAaaFnJXLFIaCRRtQIFfWqn5TxwnQK20VfmAMksqALni6WcWQwiFlPiUa5hN
ZtzgWMfECHUf5SGhRfA8upuAF3zue2VRiXYyluEL2pHRSDvGm3n0e04rP+odkE2/B0eJrJAaO0eI
/HPczNzPThW/s1N66OdzMfE0DMlljjbnXtf76VOtozD9dP7gkBoRjef/iShQLzbxoiHV6VV89tdz
JLcQ5YSyutM1qk0NeTM4h1t/2HhVkHVzJEzi4gUMgi7pmeHbGT1EgWx2958HjdR+bg9QTU2gP7eq
QsyNAQ0OpNtuf+sblX/hgWDnn+au+HO3SryHkOr1/ViaW3Q7PEbRaWqZT9YdF74J7ak1N2KoLNxU
PNgKIlBZgKNmG/BnVQnEuQeFueEhUD4bUIxLWtgri4ZUHRBZeYP6IjX0uZMPPirNAlRfAwUxQHXp
NBUpgWzad+zTD/2tUjd//J5YiGlryqGQHoyELt0M67BJ+C5r04LQscdLX7lzfdIkez1LdnCfZm8U
UuGc+sDrG3uTiPirY36GTtVJDx2piezMCr/DHcUT1YLzN6uCTrpGd5nNOvMPS/RFy3SxeoN49Iml
W7hLCP9RwjQNErShXjUKzw56iB9N+BqKpjRdGoFoHf7tHFN/OCQxwlMaLDyUMKGj0wGXM7bl8Twi
wBWhQsz+QPII8neJf912pPhbQw6146fcfipL3yM9OQdMJDeAeYIn4pV4hgYanndbcXFpCnB2/TDJ
/X2y2zXtKXbHXCaHdW87ld+oIxhaW3zuIRjS8qmOWeZeaYXpoQJwjrZUGKJStLzOzROwg0xLmez5
2h07ZwmYLpw7rUmmOSZx9rAHI2B1L+yr7RDJwaOnDgnxE9f/NYhlUvYhSBNy/58bq0n4O1MUldKf
PWH2Poa5+U2xLlSguUEeTYPqeRlqvV0CorOriZ3wzbP3NStngdQGSpj/pQnFOnZgSczJP053g0io
N2H9VMipBRBMUYPx9hfDmkRp4brrgUYsFkWUOMFquFATnoUw9lvr4IObw/m10pCDCWDiOpq/RLoX
/qfjlVpsYD5SqNHOX+8xfm1EQXIyaZmNKYgxDujwqMtbct8S38xNC5MoWLwCkfvOZr3BtkYXGYhJ
0Cznhmpc+8b5mVNyIF/z25GivJeJTQZUdwbYMdMIW7gG1WdUZm9/mdwH2km2kLUaVDe1XSoxK71H
G2ZsX3ZJZlMsCFJ+PwbhYFG5ppz4zz8jN2CxJmdjddvBWayPzGTlEAvZwNdInrNAbKMege9ODEst
ZF+VKnjM/A456i6szNgYvzq+alnCLGjqUOI1Jw5oYPvwgBYMyVI8TLZv0rlJgPA/GcwFi+kgw7q3
TaMa/AWZDjJPYB9SCf3shxczHOW4zYmaHVrGlpQDxjR8INnZbZKn3SfrJdLBR9b3XTpyIvPbySQi
r12IGMuCXSOJbenTIBg/7iVY27nI16EytSrCGN+0V9Ka/AzcuXKd5upuLD+Ex63YJL01xnITfilP
H8gh1oJ91M9bsHiB7VZbIqn0JxcTPNZJnsFCu3ZXKxZe6tMbFcDcxYz8q9JkiUZuIJzufuYvtqdv
gfomOZOIP62/BBDYW3Vl3uoyarEXmyXh9MOcOre5mgZ2mc5H/ylCTTb35ikbP9dR58zS1tPqJ2Ox
fJrs1fpXIMN4Er/PlGM3CcFgwqg5WTXC9Y48mZhRHWfS3xGvuZbxXfnSjImthZ81gsROz567clUe
1+6y4DD66duUnL3ibKzt6gCNSIetOG9vVsxz6072YnMXCjWi271sgnaydkRhdXAe4D14le60gvqL
wspIF2RCLjbC2SSOi8emz1KrmLRPYn5mMFsitdpO+C2TCKDLGyjzMU31SEhSrHkTne8bVO3km6RK
MUmZA2M6M8BwolYY/JJbfGjMWKvzuc/MH6dLx4zDSVJIW3oTI3If0acaXoSuX25MKrK4OlS0leuU
BuQHJPYj0Tkcvy3AlVpvvTKExC0Hrxlx6VZkR2rrJwj+cqZNpf/qBfmGcZBNFfUUXKA7ur4Ac005
pW4f3GYIpcKuCeVlROgqOyqzHqwYSzaMG3I9CPjBgP2Ckcd9QO7JpciKcF1eicDHxDZbbZpCTN+4
vJfpiCMQWJV/iN1ekTnVYKpj8vcp/AbJoz1geF2c7mlO6YdHBY3WHXZOBnKxYQyOAldIWUNHjC/5
UiB+Vy4svQQX3iXRHEBsqKKoSuY8pBSbBEls3Izhyb1Ltu4L8kPhfWi2wRx4VmVmLsOFE3ZNf8jL
PJ1JeNPJltu/BiLvhTrP9rdRtikCl4yg6PXtWl1o+0BmUwO7WhOlh6suMPiGcFpDxFbkOE89ZVeB
4qeSYFNYshDOeNIpeyYGTlgSPeLJ34HiaE1gX0BMBkBvCFT+l3JmJrLEiSnVDgN4AxVBPENIG5cx
e2mLPOEAEY4NXhWzRMcI0+sbEw5pd9YcgQyvQib+WztzXoOuEBvKIV4mjWG9ey5JYxl5L+LjDlBZ
2heu8rgsJ7KkZreiap16+pNgtj3m6hdUjZcbU6oafKutzuWJdGXrzpLbbv7MNkYmTJwxyUdYeL4z
SNV2GlLFYg5LpXy5Y2x8pIc35VijrswjWcJ+gw3KDmvtvNlwdIADa1IUZZThTeTTz6RE+4UCzCCt
sXCxAPZkBtWv20cHL5j1RkaKQceupoRfDk1bUL593wUrB+Fe4JtIf3mAWh+p0BJ5MgYXMBXJFsk9
bMViOYqZeWvuQo+TQgZNJad7oJG/9iuvWJhksbs8hVy4RRqcYjgAIh4n3JaDN9Uo2rT8B4nUSvrz
V5B2fARkNp90DmMcDvJvFtDu/vQuT/kRhaqopaYezNGE0P08zAESgpPpQst8RvhrvdiBzHTT1b6P
VehPBVtATG8k7yX2PzImkVZJvOpnbxvxSOns4Zd2vr13ovg0VuEQHzIfVaEGuwy5zOCr7B9lIQ4l
PNzMZQOhnExnyGMv65I6kym8paE+SjRwqrG+I/FsjR+jV3X3HJqZpLabdSQCENHhzN99au2leEAS
Iczc1cZHxGWdas5xQVs+3+CmpCIlKG7JAB6j60Nm7FYi6/i7+E/K2Vmf552s9M0iMAXZFJbC1+mz
cGRBqrcUxYvF1Poe598sg9Efq1rIjcn2F2fpD2IP6zf7T4lHY7+YXcZw0W4KFh+ehfVLvkfU2w9I
cd+EQKnEhlM2mTG8IZete+ubTQsk5dqZ7U2yxYlqOGz/wmOChMweglYITpyb4HiCE1MhKveDFoHV
sIP+C70FEkv3Sd78kvNKpOT9JOEClxo8migGuUm+ltKFnfnT1JzAVY0JytveXZ2qhWcT8wohy1E1
xuHcqX2NQs3BuAS43AnhkPGVss5pjpgwsv85LX0RAAqLG07ZoYwNLzocD77IdEF3HmQ5NLLXmhp/
8DdQ7BQAOUDvizbTucoAwRj5uqNufiF+prITR6DxSAo88Y7neawX5sk5bZg8ULdq/arPTWXFP6Bj
sdl0F0JF2VWeT/zLwmhFTNh+48OT2AH33gwLItOuNGaoIGYOqDCXxEYFax8lbdR1cI19OzlC+mYW
KYCz7BAIN5HaHGwgWCxcTBNoJGiW4dyOm8lqrjuB5cAPdwTMw4fK+hhQ8cS/aGWfAoqXenxZ1yla
neHtSiuLAn48X7Hlum1YpWTYf8+9bfCUmGaQWPgT4tD4uc85A7Wln0cFpRz2zIjUgW/pJf4skFMR
R61T2si39CUFiji8CYuQR224UWGu8gchI8OU+sjobdw4+WG8j9v8gSWO9AOZ2NjQcMyeufAhJWuN
nMI9+ZKpJicHWas9a6tZQRqyuPgkILM+Sq19p1GAeR0a0Ztd6B8i5rj6J7aKII68cvViRswrtLLl
Wl9ttHzeddNc5GKi79SC5+0bsP+0EoPBoKw6khDL1lh79oxX5vzU9owXTx9sxEp2f+5dvRv4EHIb
FFjvwfhsfks0QDTUxodjhyMyGFez4URjn3ian8EOq5BJCU8PfzRL0CLBRfb7Vl+n3MM19cEt+9mI
V6iNIV/8F8auPqzdx7inBdfhJX1R5jdNXflEXA8nk/ky+KSOwL/+zeXz23oZk7LH7+PyUEOmkX9T
EKScvbbtyqO9AGA+lkzbzecG8hlYAFcEfD0KE2UdMDDzEP8F38tFZDnyiD2udZSplCELfP2M9K6Y
kk6hX8JVVY29swWzqgr9j137REoMcyYvfdCkXL731nvc3B5LlcD0oty8W4v/J7q81o7EakOZVRGk
rPntzzH7wwnVTA7FpqZ0Xg63qaq/2TQS357o+KhBGPP/mjWDaO3PILG5x4xqE/GIqnntGkqaU6uQ
xQchBJ7T1DZGcirO9mizaFkNHahzfk4s9uVRx+6hXjUwZGhf3QIakhnpljwGvg9gTk9Z4DayTe27
A3kg6M2qaGdz2zbomXNNMMIKZDjuZo2ZR0nyc3uGAnrgs/PTD1ToOHzaEc2jcGuYBYjhcT6TWQud
cxNUdkTYN4/8BM1SuFkhwFiQWqHDvUDmPxz7dHhO71AxzkkbMYsEhc5rvyUhPK6DV/qLHL9gK8du
RZHOL5qcFSjvqLzOLp3UvVOFwHJhL057xNrOhRWZ3FaVlg21A4uCRibaMapjPESKZFgRsl/EIFFO
BYoBuDkxnTUY1fDg/gz9K01XqNmBCHTD+uoI9QI2KruCfn7v+ODk5VQHH+srsHBaxhdchgfUZjV5
xCfnJIsq+q6glcu1fk63K3jiR7VyFpKlTeHYR2l6XJl2mx+q5IlEnH5UnElX3gWJ3XAOalB5RIN2
oD4t8Q+uHPPCKLiY7iEfy7X7MYhZpgKhELBebkGBU6J+7PLSTAUc0lMRGmWzrNKGht/zJIJB11Qb
V4RHRnIo5A2DisAX9lGTK1oFrVGIQAu4GcqugVXzNUUaI3GYecITFLlWhadk/3dT36k7jsXKXjam
cfYKG8KM6F8hcTBM8one5HemFCl1d/EKKa/zNKj7SZdM1jP5clibqvwO0YvtZJoi0EVM08RkKEXZ
0pUjRHhdiTAWT4qks5YGVn4H8dWe5LhufYkvyw+gyqGWStpY9DkO1qbbBMc6xq7/YFthhMFVSrPe
EWNYRcFjK0wedueKYEC6hJQONoqm0gG+cHG81f+EHjR9QZ2HtnyQNCoK2xu6KRCK0p3pVShbe5ua
gydxbOh1M1i+xXHjVDEXJUheB1s6gDqMvGSNo7c9rhzH+hZXocWFMiXVXl5Gw4oYhNu7AneJL7lP
jhCxJHEv1x+zEyT93DQPXWnXc9qthK+QD7puWAlW+/1NoiXlmewn3ZfxOpahXaUDihgIcNpWvGSx
8C3Jpx/zXFq9DxVUf1sv+vs6bCILde2rG6Hgmi0z8vo6XweZzgBBcBuQpKf+2BCFE1Be9hcX8ukJ
jC9kID3+jrgEDEjIClFk6legm/YjddVNo1Zbddrcq7TfJN6RDuAO0/zpVByml9iHn7CKSiypsTZE
3L4dX0mnY3iWLXZUtT3DnXErJAdgUoLDKlK80RL4WP/XBnPD3n5CiuAFrw48r2IBseC9exgs1Lxw
rR0StuPk2gvsgkIUPzpxNVcqFu8KU+vZZmpgpO7f481i9+7Z7FZfmOCt6dsRTheZ9y12mFle4Js6
DTR/LF2hKnjKNJ+XJc6x+Q8tJxaKKotilACIEjA82lFNwylkBPR4VHqY9vN4cDbaCWViHpR3osLP
mv1MMkLnLx92cXGH4GKl89SVcp2crsG8/h5uxkTf1vfKOoE40ZCaZeYZVbCES5dfycv/A8pfpueA
vYOwxwpMpKaUEbFyvXwd1Cvy67YYlqFV4pWPaK3LoV6DyegZ9gX3rdfqv1eKpWEJEhSEtrOUPaSz
VUzP5EIODbcxcehTuempTgZUWfDLBidU7V6qn5iyfdahaZMSOKX/IRyOWerlcKj+CbyXd7TrcOER
F8GSAgyarURZIU2yJX9klMApJ28pUdxmcGsqw3TkK+wZpgGrG+TVMxdtODbBFCUFsa0PCMY77pXV
WSf9v98pU61LESKFciJrGv4c0NcZkQsTZ8uBqyfmUxadPl/whz7Qy7bm00kDWyDpaxsGKy/2lGuf
tDr5c1e/bQFHCozywG8I23f+Y/l73CuP+Vome6dR2229DZiIqdPyyr2boZXlYXphZtOIMni/X/4G
kA0lXAfD7XLdQSm+IcDtFBPysB35SONBgpkXNLSOGZxOVnxwPHuEWwwpN8cBzScfqtjZAX+hmo3d
AYlFv412073EqEEQYJ1SiHYGA9etJMhhEN9aB8P1XkUQ11XJbH9q5FebOKVx3s7rdCpy+TbPshiF
nD40U+v5lABRoLEM6qMwHi6UFm7Tq6WltWIlLB1PVT3fQuLRI/u4Cy6lX1AQ8S2GHDU6Wq30YFB8
c7JQFS4JVnss6bmeKL1FoCH4GzUt4QdKwFVg1sFnzm0ow5b7TB1I9FRM5j7K4SW7NsOQCfxa/k8Q
BZj9hFi0oNHr5bKEGvvFHqoA0G6p3rmdCkkysFwpGwvaqTHogx7hzPvpQsQ/PNHcd57EEHESjsZ0
MRJCL75fHKvhfPFfjISb6zYNHRk5Bn1fVuQ3kBH4MFNzX9XQxpA5L3qTy4J+Jbn/YdRNVMctCyf6
qOOY1ufninKQbk0wYIAytMO59QC3SCWFe90vJq+6WDHT+7wNNy/8ioeFyQgVO94zq7Oj+vkNjTwk
Xn9prRKsRlQI0yO8Fp3TWYydhiX1RhzaN46x9XK7yUXs7ESOH0KuKkQ+940ol5m1GU1m4h4A+++U
pC1mMBAdIAf/ra9o/+wl7xtZAVg47wNRVU5DO5HCpmorM36Z6mMr8OH132SrGNqLYTqc5rp032qW
2EpxwrfM+OoVS84/bDFEN0pC7slaTSERK9K2k24Rh7KB82kwmIP0mkEENi8mno7tiX0M8GCe067L
/QwkCa7o8XCjg6yvT9MnrbKcdLH0CQo3KPtGv8mAr/v4xzZ+FpNFNeZb3pHvOeackMOoyXk95EIg
v5va01ia1jeR0Q8zx5aSB4Ecv8ErXDhvCH+G9mrI8jPOOl1SIUPZ9C/I8YE/nAkpgBBOBAxwhVsw
DDMnG+jx52Esb/5HOfKm299LOhpXSirDYefOa8Q8Rcfw3fZVAfFvGyO5tbW9DS2DmYVjoR0VrvP8
k2VwAuhEAYHoqX+E0GxVOuSm7oYzN7XtkKGIqf5qd2Hy2SgpmoCt2W7miGWcSTkpXgdMdxUsIws0
I2X/hjfvpAYB5Cc88wEX9t9rv9QoYOd6QWAFJFDeN5Gpwu90+Rp7NImTogmLB/jwMkmb+KLKIsYF
9Z7MkRpGK2CL1A5H6fzte6xkqFU7xrEV6170GcEWGbVHm7ab5sxT9YY2rZ4a9JrrB3a0yDavur/u
08qyiRmydVag6q8hoctmffnFAP9ZwdX0Z3kzYgtWDBgFMd0Ia91lYZmqlfNM3WZac1ukMz87TWiB
GMQdiPo+LRzMJkO4vAGxrU/gAd2sBLRpRG1EczBn4M8zVsgqC71hDu5AFSOhsunz+nCSZfrJoit2
etn+33Dp8HLzwxt416tdRaoIi2isgBBBlk2iNwghfw8Qk9UgF3uakqa3p8f0gdBvxkD9XwISHm0o
sQUcpiNa7OzM5SoyjhWTAGgjefaKwjPLx/g3nfBvRV8mgsbaeDoL8a1t3/nkDfJwpaFgF0l4+gRi
3osREplmHm0CMUowW8m3h9VtktrpSNOJe2gl8LRa27X3iUcyALb/wk+WHxFGGbV3FNaGUMh0Vtwi
sfMmEWHPPqrYnWFI8MmQodCAoCouAkHnu9u+PquA6sGOpMRfohfoBlmB3czOteQhqP6xrUo2ZMwu
0HPA+SCoijLSUKa4MyqDSZbjULrFcqmQMom1SaVIB8XJbyn/acqlgdJdNlNvOn7XonQCWJMxik0n
KT7qfbl4DBGKa9XHafj5y57CyE53VV//FCutG2um+qJrfQV83gFKBVyH1y901pBwdx4Z9sHZegp6
Q84A3GEyzyBpgMTNh3ew2u667epJkI6xZPJ5TBs11DkI7bvLIvJh6oUclCjztOYRgLwqle+D4js9
Js/W4T5DI3mNo9Kew/DMmVBhJHaDmU0i0m4Y3mo2B7qrcwbWfsrmIViQEaHICgGLGqPFC4zTNwCb
P/0Oz6Po309Si29QZ6qL9ICGTfQ68MSluZ0edqiG+6Xj1U1N/Bv9sj53xzSII33IO1rEj0W2iVZc
eENDLB/xBBQJ+34ZCewuXcxVi+73HEWsHW4UlK5Wpg85mY9cj2kM3I22pedHtGD/lreUMUVvwsBX
D00G0mF5s3WrV5qWpATJSzcQjycV15QkfBA+rKMj9onPsUBbnPowzZDxSv/TajifrQUqagatvWvh
PugjYTuVhlPtKiWPJubfv3qa6CUN78j2IVJNRefMPUMaLeWK6bltFrRHfLkb3xiYCIPMdB7Yku9O
ngl/NzH3Fm7zI8ATCO1DF1RQpdg17fuAIGKsyzBw5mHQgrP6NljOanNuEUH1YCAX6YlJ3PcOCig9
gFhpjS7ZQtjudwQ0jCVMJoTAiutukRrt51qthwDDfkbWtOJ4uyioRDIE6BBLDMYfDvmnFSYeWils
eHb/5fhnXx8mNx6CKnsI9PoykAcSKuRaHdVtjjhKQZKveqSs6/dBdLueY34lQvF6VfPeTopTEzr4
XiIgtIBEwLJCqLSa5mhPwJ+r1kHiGyoEi0s586OF7x+T0gSTBcrcnCTKW85Fxb6/ND2oXduurz7z
yjsW9aO6BLa20o3oVXQXBkWhxbWNZQtBL2twmZ/y4GV1LpBImYQ0Qjb2mfA7A6KT6zEmv3E8b+NL
/N+wy6xeAJFXSoXmSesQ2yMajw27R+0aCZ7mWxihOcpzvcoXcgXAGGgbmumYXf9E05uxABg33IqT
JrCMCrdAJyDe4el3jYl9EO8VbdKvjWJEx852MTvn0tp61m/jfFveQHMYuGTO2glo5WjySy2RK683
W8k3pCHPEVHrJMYrzzffvjtZ8y7RfNz7CWPFWNqnlovqpyJYvNAC7/Ksw907BcM8z5rKAfLEftC9
Qk5QdT3OjsQ6EQhD7IQZXulzxtzkLC/2sZQEyoUbuQXKDoUb4MO+ZG6nkw3plDIbf4t3Vr0rt/Xw
jzdIV3zV8nh2v7R+EQbW/4HfZYAbskTv5WE2GPY0kzYoL6ykm3Mvt8Su+Cnj0jGB5kRNY5uNhlyv
OOZKyobu+54C65FC0TAVRFpD00VzOh4NiqdnAF/ud5rc4d6p6SPqrfM7VMZ08BsaZi1j/IALlZdl
vuANpwNN8LdKs1aTEh2qHB392r08LOITtwLJHD1XGtnkLjNm7owFZgJyXbSoWuqxHfOakMfoez4B
zbIgDsvXuRYkmI5bMzB+/rDHszpbHYPkhrMXs2vBsVDiZ2aiJ5gPBDKknLTH3IdG0zVNrFTwVx4N
tAO8PKJxivVGphQF1DuE6H0wZtyMciL1U+mhDgnudYYbN/sFMapz+Bcakcox+VC0GEK3HTlNEjC4
XBDjPYv4dwT/O/tU1369h4bSYWg3rE5n8aeU28FPdOJamDPixT3LHLmdfnI4H2XJz646Y76vDemE
b9cKH5mrNXj3N1cIWfPXzf6M4oZEeGtIpkXoMT8LVgYSRd3WEOIINGBvRtCHc+5a7ZzUH+VQL/X8
J+1t1OZUtOx5KRHAfTYgXowD9n6f/OK9Ijvy8SaRlM7LlyiwHSZEyxkbyePLTmOegdI2JkyIDIhS
zCQT0ReBLJYP+VFu/qIvoGnudbBJ3TezYMR9H7FKw8UoktNlJuMVKHXLNzVxcF5jrv0jCd4HvmtT
ndX21YfzrfdDyguSjSMW7TdNyxB3VyYHcRqMyp6KNA2gL0YN9uC7ExCqwRAZ2/wlra15dTn5c0PQ
O5C7//ecBdydE1QxGzdpyqvDxPUs1xpG3hPsZpJDErbDD2voKESXYP3mZI4bfH3gDraBU3FLH7QY
4OqF/ZpCEDn3wPhOiUoKnQ6V3AQDoapP2r3m3sDaxJo0hKHpnqQMUj55yOKPQE0bQp2RssziM5b2
OIiHWZUpAqFw6f7tuJxQauvkFml3MsQ86NvysXbTVPgZ1syVG3IHKMkuK6Ii/hF0XOdycWQE3j2s
ccdOBfs5g1UKPNtOWLnJGOcrgwrWvzdP3+tx9QONGaE61fSVVX2E/wxPxEv+wIjVQhz8p2by9+O2
oxiaQLXALXtluYkooOzUuAzMfGPTb/0HLTUoqIzKk6eNcumki4qr+t3SSVLQbdZSdyXi3R+LFDnQ
24pKmFgKC1YxHeP7wdh1FgqRyVt2nuZQFQkTdVIi41X8lgDdtLUVcalxS3ZSUjePfgzomwWMOOhP
mzbdX/GlXgCK1yr1gseYcnZ+U9vUaJxMJPboWaKhNTk3k2UseXVsrtRagwNHAEJbSZ8IA71kUZs/
hZqh42B7y4KrIt1x61GPMp3KbXE9UFrOUGgs/sNWFNNSPAU8bdpG5RL9BOr6hZQYGz5wzBrK6XgZ
pHyiB4PXtBiF646rziEh+SVZ9iVOYgyzUSDTGb4op8OSg0mOeFnnMjtZjtoBhZERgZx6un+oB6N8
jLKUM4LZxji0zuwhhELVJrQahvUVAXyNJQ+8EsBDMeXdeR1E4AF8amoKBvGPsA0KwZGJs6ITW1S9
MOieh/Am1UeupF667W0ODvTEXghHuKgJwkuN2/+wP+EEWdaV/9+pAFNjnJ9VbufjKZUzK58uc6E/
8BmQ61JGU+d/MSYKncyZkiUY7UAkHICsLMHhCCpTIHdsRK2G8bIBDwZkyCcNdc30CD3KLutYPVYb
FQjRTZLCLbvaWAVqKbdhxrtPOjNk/V965jo7XXolvmk97JzU2OUH4M+QcxwebEjLgUQ8/N8ZW8MJ
aAGkzX0lZmlhe+AIl+nDlZfD/hnVqZSXNqsQRKHcKEnL/khzPeRB/s3xOy+l3Njw8QK2R4DMhA+u
Rpw+s6IXaIXLpnB5pS5t0xGMnFWM0jqRaa6Rx+sqpQeO/dbumXEOq/6YcuXbarpYrv92R812dny5
w5rVqfZgA/FALa64B0bRthcapV2YajCNpqSE/zfhghuSBfNJ1ulDxtdAEGu5N/3X10Qs6GFpCAiC
AG6D5aBdSiKUJhtzRDEwPU7B5aEoaIjccAFh5+LK8/qdma83zgT4pJTJPJipuauUWJeityrz+4yk
G8++QeVrU7WkDZdSa7ijDibqfZPcDT0TP58QwYfKwaajAZ0GsZU1F2bOE12wsHG0Xx47RyLPfaK1
f8O/gTT05hSlOdQkM73oI7O/zxwcptXXc4UQUFkq/aHeIUVUCmlKOwPltPoZ1ybl9Lpfq8L3uBtz
1JA4qzVekp8x22xT427Xk/btRDf0BO0GFWbO476loEslTEeY6I4Kz+qQec4JKMtTLx3MUUIecGuS
f20B8obgAvZjPl46C6ntQDZ/mQkeD7mLZGKZkXw1dCWCh2ahuF3m0EHdTD/dTLpUBubCvV02grSw
/M2jx0fl5FSxvNfwqBNS2oGSCK1Vr/UdSyQWlYE+9y+Txon44BvEbB0fqerIh8idVlaX39bKh8YH
2xMcVvM9tmC75MPftDQ8CLPyfX/PtMDfKNjl0dVD/Zqn6REwy+O24P5mU+EYQqH1JqDcP5wrU29j
ywNSFG+1t9KH4uA9zYl1qB0ogwf6GdOWkx10gZNGXXrdLLmD3LB7c2tX+eM3BWWJ8LP8gtsw0ksb
Orh8s7ZYejTSxgba3PbSUSnmsMQ3x12Pa0HgF83o3XnE29S94UuCbeaL7CKkVaTrFzTCw1UHtVWn
D1PQIPOaemEuo0Ie6/01xYBsQmwy3rLy3G7edfZoD25pMFP6nKjS/8CTM/CiuDQ0MAks/0DYtRsi
qTMSu1p16xFCP/abYz1vvP3Kz8Eqb0FugVX/Ldc9zxP56tK+GNuV2FcyeSAfehzTE+RMrrUItU5w
qctC6L17tm75c+y67+xhmvxEv7KXBG72Y/K3tYI8W+NQo6tOU8AMAp3ngBcaJKNXGo/r6M5vdSJW
ST+rIl1YZkYaMk+8BBQ1QpX7czQxYU81l2Twc8bosrGtKYiwUjSyyLq75dwTDYNvHpHjvEvqi7XK
0ge8VghynfVhU/uxRx45OzECrq9zlS+fOZ3kdh36ybumz/qAuQkvFpVlVhHGU4ZFxSKya176mK8U
6DO05/sI1aQE5nPbu4mRbCpWaonOMxO/IF6k4A/7edik0pu2g1dMNzWAAGCA9TY7j8mpSUUkFBaW
PKtGnHSBtdsgWI3GxPguAcuR66KDGb7Pm92LmF8QjTYe1oOVFUMww8fZBtXqxqH4M7Suuhzwt7yi
OHZMa1yfcxCEy3wnhyIooNRdN921zvqWzk7DXftYHsilcLY1mEiGSl2QRszTbhrjP78g1lM7CR97
Ec3nao6w3mYltCxDqRq8uV/2OGOR0OiQSiNjNgSo3ldlikYrmEDqhFCefaHcehNNc+XJTpJnV0hY
rPsQFDL82w9aa9FVRxjmw4kHmWeyBRBV3/3uHpKBtx23806TNOQr+f8FVGF6VHnDm66P7iJB93LC
O99mSdvTV0CBH8zNfI/mOZgIYuYuNAcJWFalQ2dFcIXuq3ZC6OdIoec3loRFpKexToRs16CDQKZO
1MGwecAPNN5QtYSTVbQ7ONKDn/byFbo6Z8WG0iZ49pyNTjLdt4JJYyO+x57+p40DuK5A08WXFpi+
Mpz679sj7I4ec7buO5+Fd5bAQYzxaFmH6CROpCCw8BTNrBgG57DkGymvuw/VW8wb29fVClu0/Nbi
hoi5I0dlbIRwiN593Kop0PndAekiWsvJlzwkYyURJ/QBNZfk1RA2QbnlRx5TI5I8feOyrs7AOFwd
oRQhBr4f6KoAgtQZN7U7BO4hFnsb3YocEaIIECc9X0R5p3OfXtdyYQlUMfE5JYQ356IvAmyG0UPO
XE3WBYdTyMdUmRd9TV68mVlOyC3Uz9b8Dj2MN//OmdzvUgixXrQz4ROkF0RPe8lTu7XKs5LupsrZ
3Jmhz1Eg5gKn8TxdSZQbp0d+Ls6uJyYd5Ku0t1RvNtzdOd2zX6yTuAMXRVlG00DLfRxbc8hLCsHs
V3wSRZNvuKqXRHPdM2Zz0yscdInQWTBP4B5T5ci8lqDqtKowBVAtsL48zFCneB2I4O/6wSvD2jsL
WLCVkz27cMw/dHLDcAyX8qWEGaPCqubYYGXjOMhAWG70QVmQYv61PF+845IQkfKShksUMbXj66Xz
g5P+YrA7+TdioQTkea0zrOvgSARLtTv4NTUqjtgwxhY1v1noAfmSgR183Qde//HweL5xUUiytdZG
0EKKxApFOt97AA2qgwx4QVyv/KuxqS6Av5Vr25vIJyhG8WB0LhG5xdQDjq9dYxuzoXUddk4mO4se
Mcpeu+cmMeaLoEJsFjZklth0xpWCV2on1TWhpYKWJzZ7mLdfS0y+eOAsaeznYxgpc9BUYV5y6Hlu
2MEKKDaHJcEVfe/LfJ6jk2mHBIxiYcpM/PP+0jLw+VTubRLa+fcb83BjWBTvB2IJxQWLAtHIpkDy
gpiPmQ8jBot1eQQMlkJ2IsXzhyzDXkOmJOXsqX527yOnZsT5uRWfBA2xo9AUKfXWNiiqEyjfA4eS
Ai8W43yO94J0HMzzh3HtHe5T1TYFs0QbcDOX8HrbRiSUWW29K2bEsklP4H8NQfNHY8SBXMeC9D1K
R4Wx/WCF8nLG/I2aacDeIU/CGscIwq1IQVUO7zkf1EbqBF/WDMNJ4X33oGl39tIEhmm6cUrVyeJU
QNAx2lj5OtUp7FePwwYlXPxX5T2YGrNJjkm3HU3opMnDnE+AmkdatcNQWkVTFHZd5yvsbKZ6H8/l
nCSR0H20tk/UzQ2tNJbwt1INdO0tOHmGU1iuIktVmcfcVKQyTRfVWa1vIJ7bNYH5muJpibpEVQLY
+Nfz7UkR0HGyu2VoMj1E+8qO+yzkYJileDnF8/qA8RAIZZ7/0AYoiyyzccu6wsclRgfnleS0rEPG
I6jdYxmTOsINNAX5jS2jUn54QhnmbXq7qFraQkP+M/Ij05VjTdFOUNih+ecZN/yBJf1XMcJZ8SUB
q/vO0OIcXi6YkjA9HQWg3G7FKdOpX2af8u/quu7UDaEEplkZgPTXY4bvnDnbn1CiwoDceXHTLa+g
4EBeRRp1tmUA/9LbkBRnQsWUptZ36r86LRSgZTmuomcwpu5hNZR4Y9HYMyT07dYV+DCmt+1OyjP6
cWhc153XDOjd7Kfbl51ACknGpbtJ6c96v/+u36LkB7AWk6lKgR1Aat76pvJ3fkkM2/R/mSeFoDXE
85c2yaGVkXwCa2Bgfd77XMS7531S6IBLg52gcdttLSzVsr6cltRKL3qzjza8sXGlF/Z0qK/Ruftv
9GACAkZKEvumpEvW6EGHz+QYmr9Enf1PJB/rBQNGRsEr4lr3TMNLIDhOc02DguPJZ8A8SjzvmQPm
aQiFFkAuBhw9XSN3SNS0jEANibck+eFp67323mf4a305BjJAtGi4AGdGGT7g4Y8Ui2osvyDiH9LT
zVdkYcrTNUBBbpfzRn1K4QUvAPnrY9xjp2ucMjg21YasHXGCfTNgbSz+lvS5rj/tvHuqJ1HgtJCm
h4WvFtnGtcDOz8O5F0G7k2ZjGSYPdsIfqi5KwVo27pq5M/0L4TRefjpeDQwLYowu4nfAs0ZUenSH
dgyITXD9hz65lBuwcNuL5scAZLLNZHb8ZvNpBxeFEJk45EYWG0omWneuC4Yuul/VtF5wbqf4UHvP
8MCQGES0CHg6rfVAogLFmhk3mzaORZvhSQfjoxOE+5azhLPVO5hZnS4KPdIjkcpOTxIQBJBCA2sS
O/RSZDFbASzkQ9ydt0vopFmdCFxk3HVi+Elm2wxiDdPIb+lA40Ww9YbYiaDbDX8UOSRTzNZVrKLy
Qg9cUoE8XNidN6wyO8QFnUrrR/7tl6ZKMjN6M05ASwQlBkvFv+jVQ+MJfk3Y7fF5naykEZV5wEZQ
N0c9rIeGnsSpt2n61Zzk53CbmL4g8+RtcsV7qoZHUkRZOY+wXyEX6nSjI/uFsxXesY7h+FgZRaUe
SHc3HPKMDWUJOtGdyyFGeBclPWeTLocaYHIzYO3Kne+c96kyEFCxapcFXSvbbClvTiHECFSdDZG/
Qi2/TidwWb1G+KFHlLT/X+GE40pfTkbliUlNMfBtQ2j9zSIQvn0LBRgTJE6CJjoQEgfAAAoP0oav
ZDJV3Tr7u4oTW1AsqWv4ecC0DJpWjfLgw8qdSY4HABBG8R2SJu6Qc+thdPMHJrbYykKsXeHG6l6r
3DAcg7+Q0IW2hXpDeBBQ9d8D6vlHGR1o4s1llzBBoJAfr31WcROlQtQnXimCZCb77VvhpVe+iwfM
RdRgAIip5DXIBQPXoanNABuOKa1AKGZSGEph4Q/9io1jHpKag3/heXEzhKp8yuNZDwf/vwwwWcpg
jKe4I2VZWYJxVXoegPQhgIK80nEeSinVJLjIeTWPPvoIcDRIulwQd2vV1mvkL7ZIDyUpz555hOMi
A7p22iZis9uCV1g6Z74jhskkBCSYrDkA6YyprWpT8SmMAknFI4TPEkIdDTdXG8aqmt7fJykxNXRQ
yLIS4eOAh2uwWPJXL7RXse8fXP0XfLYIUeIKRS85XCNBCB7C44KK80WYoQbiFgJRI83ec0mX+rnB
OzXxQRncYVjVh+Y7RsKlcg1gy8kWyEfUEyL/fKEDA2gWZtCTF1pXkCKEVqcNIh1QlHDy0PvZQWGa
nc2ov8ydvFfEcyMT0JuCiyGOYAmrJ17S/NLYnnOiiv+aiaBN5uBcyzr3oq0Oe5ELgZdMIBelLSeu
GQxpdYw4AJaDQMAphktJzD7Gmu4kehJPTfs+TGqz98c3gMnQW+1vVan3M7QMgAu30PcM52cTZxDs
0FRym83f717sZdu6rMG6kcVVHqqIAM3CIEchi6zi9mN3K1839BXhDYgTORpL3BFmGeCyLHoFEQRN
VQOccZStmkyoltno/SrlsChSzWP5B5zrGmuzkbJqeBxuMpoentjKiQ0MjHLPfhJqREtF+8IPm83/
2/EPNTbOh9ta/04XBAurh37tHmr3D89wFG9PMQhAyiNbWZ8DnoLs57rIU9uiZZycAIDdCH+tV4UR
m3A+S0KqeKXnM3Rcg6vO40piDZh546Eo2NCsiYUrPANpnqxbdc18x91WjDNTQprXVWXRbEzRthp0
+sDBrQvjWPvdNiIhqzA9Du6SW1uTwjTU6UhmV7YlfW6CQctD4EXxgpqFFa7sHqITDkG+mfE88RIE
2H50pfQ6JciQUfOjGKi05m1v5xVcGmQ0YOXj8hyt/0ekQlv9QUuqgUgRpGo2AWMiXxKcJKJaHI2o
KdTtOd/FyLYg7bU0hj1wncwGbIaMRH81aH85gcCV1zelSbfUqXr/QkXQTinxlz3GXDATMiWK8g0o
fa20/kE6evYrFhn/aRKIi5lmJowZ7vSEBYnjnb4QbO9T/yEWsFX6R8OJQpsoMo52Pi8NW9VYd9zQ
1XrDpQ5/K2VUJWqZncbrcFuS1E0vGWJjoSO3DeGZwYsJ3aLkcQkYk0h/FkQEdK/H5J+i+7lK47kI
TTCqgV4nuJ3yWSw11t6/T1xXMeE7Hrhr8mCCV4INCO9QcxboV2+/jz8MgikUTfbCQQe6brf9sAU5
yvbHwkTOPIHzIbm7/r/pe/Sk4tMjWPnSLfqifjcwwzRFBPSMwacUJuoUOpxA1XDhVVSRo59WDEtq
O3EEF5bV3iIcGC3Zzy9aDnjSSx4/a6E0VGKIHeJqhDyXHhQxbh3fqQ6ElzK6H+c7ZHaHVy6LJAeO
5/hu6I4Eiv1DiXI0+g97VHaNDIs+4Pbdqtq+iu9IxAWEvrNWDHeqbADFuf0iDMfp1VKUhHvMkt9G
EtklIaPkD29ILlocMoHBk8c9RVBixmc36ArZWW5hYGSC6caZ59t+CNbN0bSZGYRx8cG++5A4pn75
3UJW7UsnizHDDnVRwHxk/8O1Gmq2VaWJgab5Jg5YF8chNNPNjVvkKnKQt+XE5q6o5PINS7l4erRN
JgFlxasbmxfHkNZExQBS97P4mRyII20m8BpxechYlMSL+J6I6k761EdgBkmxj9bE9gXAE0MlKT8m
8NDPpwOio6x5KdxeNMVIGf1HqvxFqFLTreLPtyHblF7zEvdDoM/zI9xyNqVqBVy0TDpBIwAvQ4Qg
eWele9PxiC0bZ3wivXwjiILyzcYCitemwKQ9AX9o+oCqOwakwdR9J872yuDZu4WdmbA4vcSquauG
WYg/5g36252hbFwncP67H1mqdGYLAWNhooQ2vf3eCKrgRwIPSaImiUV99zDZR4imjJe3hrCW6Jvo
w+q9QVoeoWHwdtMCCGHfddq3lsEcTcwmI1kC/mZbM4Upq/Od3FUuKA2Yur1ydBO8igLZfoEHQL9k
1LL2a9tMv8PAMW01H0Vl4Q9WltDD6YcrBNWCr5dTbXeMU6UnQBoImlDOcE6XyUAvlHlbZIa5HQgW
UWPUDBel4Ow5AsfAU5C5lZ80efVdqX3MShi0zh63YVO/Mrecn+P7Ft2yhP/ItHU3towaZm4m8hPv
y7CoHcP2cgtC8ls90dhX3kD7AIdSMtGVxfne4cViTdFpv+ZWpkDW4bxoeoup8u/gkE8ysIA78IQP
BOsXqfujuEyhgkDiZW13ngzdAumSgmHCNEvfAFfGMrvFjeaLGHAIezpj/tHlyabCp5bGGtSxbVqF
vyxXp9a0mefzXE1Ko30TPjG6h6Mk4hYvOdlbq0gmI4dU3YIrAb3aAIgfNNLOoThdlXllnCXJezd1
QtcqtfmFUjnde9Hl3YazBsNJ54wZ6wpaCbtBn6+o+hdsGzzmyh1Lhah3ouzWAAL0hg0nPSUT8X9j
HuhbTTabTHnVf/jmcDvKIjk9dKNc8ezWXfqRwH5fDYo1dUikA52e4Hg24it4ZTyyeSM3s1xbsk66
8dr38uoDVlo35l1EqBghBo/d7pUQRlobYM2TKCuXN7J32YdLhBbWUxQEJtzri3w80uw5M+ohiHXz
SGVYc38IEsLVeKJ/E0FLrpn7ocwtySy8+2CVa+MXjmUrIo0O0JtgtZJ57os5Ho6JwwkBX/L6xRXL
u0vVl+Zbe+ndCDfa5WCUOEA6VMXWPt4WZW7TQRaZh6cOM/dHSJ09yHwZVlWWY24PnHpHBM2fS62C
2aA2SsPuMH+6HiPiJe/vXvjAzbJLsXIxOIL42aDBy67xS3oQyOD7o+C2/vUL7DcOs4afbueTLyAL
5uQ5VWmED1PojvH7RqvF8fiLg2KhtJNy/M9Rit//fvYQcekwNsEt3T89WziFfP+GBZBHfwD+Sett
ZqYvUFasBaY8cCmZSPNmKCnGBtN41Cv8+5FlUbNy0aZ4oEVsk3L6XivrFLt+9CJNMBlPO+pAwlSG
pMOulb9E3e4lrwdGN5DeXfG+YSIe64fxzjIbwUpaE4jCU5Ud8epG7lcLzDCrBwXX66Lhd+iJoZ3+
cmmDR6RnC0RQB7OfhfLjPK91RabadvOYyc6dGi34WOe9OwrhmP988hHDdepVsBcmSVs1UBGT+ri7
WUOFOUgIXWe5gbeCvvHwFJU19sjrNSVNHEgoRJMT5ewkhhuNcbBgXgWhSWdkO8eZaWH4en+Fzw77
NLVazETYZGgn/RGqiahlQaE8AUdc9IHmaLumpCqiW/6P4bmw1poMNvMk1Fhsx3EK3U0X6DhK5Y8E
wyTJPBHKpVoD9v6KlKfVjoXRE/GUs53Pmpp56MW7vPerv0PoBj6z+4dU0PydKFjX6hzisOhbL6zj
huVjT8irNnfjnaJlyZpUSmaCQtv+AkDCZsNAWMclTL621gzXkROChGcUvncrcs0e6EHY32JAwAq0
sV6jDnMSAua5Hs9ZSdInjr/perMdiw4rkeCKVCvNS6YMtV5W226U+hJd9HMdLjGu8xrhNMprlcFO
xf+EeGdx9tldxcWY202Tbuk75UsbwxIklh4tcxDjnQOb6vFuIGoBKLp1GSWOr43ImBgUPBCABKYe
Sx0etoXH2KXONJQJGeJaDZr1XP8t8Pw44UiVGJ3tf7pL8GW9PZudXpIJUcfuucgHe1wJXNeWmn4I
js7JG8QwJDMojnmLSa22jSktxuV/dTfD4P0b0Smu0/uh1SMrbqoqWo+WH3m752foiULWX0HFJ5vz
KocDUqNL48mhs0ugXL/p/WOShRxNxdhOyKaBKPl1wJ4FVlBofwTgIKqeVJbnNcfCgD5/EdjYm9SG
W6p9LQadgFLZ42eyiqzaZijFdUKTno0NmWPMj1Te9MIH7Tb/OelokENBVco6NVSECISz3PvjmYBv
fegb333oArrcvFC5NkaXd0jyDTCDuITy+1wEUFbpXZtpWPvnEtMHXTQnEX/e+fjoneJF/bPEc1Hc
tlSBTg3XfzrQZwNBuK7bqCZyrQFBWNiRLHNFdhd3CQQntWo3xvn2PsmZKOe51tn/5pTGa+osHr+v
HE2RtWmac/mEmRHQQvEMypVblfu+GYJk57rSp8mwqYlLnveeQnQzr0sbO734v3hcJTzb3yjLtVb7
pBDln0wGF1WtDzVIienDo1ArlE/kYKJXkO6/LyVzpGXnqrQbnCA37p96gx1ciV1ijoYGiPghTnD/
mVwe7R7KBA+53b0/lfhSFVpDooesdygqw139c120xs3FYaceGeJ7HjRe4uVnUip+O+okHeYktB/i
j8DONPxV4f2x13WIIAW/e6isk6vzTwtQUH7kvvK/X09HwIbIM5QzA64w160JkIHO2DhRUR6mIrov
8aoG09A7+U8mxfJk4YiY52lZrQBcQDgj4whAjyitZUk8LN1ulr9UFFLtpbE9Icp6mpbjskVewwUp
NrcmjIw+iI8+6+6vvPFCVLjW379nWEHVBq+hkrn0Q/TbF5STfZ18yWIr7u6SIdK3/HCNQCiXZz/K
+j9H4C2Bxu81UYLDOh3JQKeedJUZLNhPxq5BeLAEGtbQYQsn+lIQW2qjP/ONVRkrqZrfWsAZ8Zo3
5JNv97/gCdiCeVrdA1Md4TXhmvM9OcA9rh8qyIjHJNFm4AoXsxaTjXyNVbobB+U1icFU2GXwZR7h
V/b7Te169hATO4FWmdG09irFIIDHtaG94ZjdSnBZeGyiNLqdp98fd6WyQvRaD2ACtBNfV5Hfypdt
8u5hp9Im0tXSiuvQezSgcx5BAMczJmKvb7I7lLDovH1NM87ZSZ+VQto1fEhC7JjU5YOYotJJ8RJp
I0ZedkLvjbb9GMmN+cIqT2+J/UrbfLhYoaGbyjZW8jb3fqqP1gSnvsUBp5lg5fDaWafq8+sCM2XB
hRi8c3AXRKEphufiwfMVZpdV9CP4vhE9Lcsw/C5bTfGSuxfngSuJzPTkAxP38v4FmFbuFkKkbKv0
AKroZkVGQPLPkuX926NxCaVUrzxS9lPvtE5p1FJc7AqeinMXQOcJsmg6lIrY3NaDytg4EXSi4jfk
sylMd5RYLbCAQ8doMtjs46wiioo1acGLj6fp1H3f574YnTUbfJZHHlmdpKmMOZWwgVV7snLP4Km9
1aanp/stmPNxHhwvb4vVjPBMYS2cgIvDCofY4LAAktF24iCQLrWJp/jKtEZYYklveIXM4GJ4iMGS
0xnPAjEJszIrUpx/U9fsKo7C8w8Ovygn6GZ4wNTrG8O9bmjy8MkbD3L1q/ihNWHxFmFsnZiXlClt
CSLG6r9oQbTtv4TGQmqtjZuhY4bjeaS7wa0OygDqAT5R3GHA0lf1qvIQPm2SJKfEQl9XjjubbhO7
B+moq/VXVBvJoo1gCUZP0kKBSxtOYI2hpquJTp1dWt2xEY4uC0OmOT3+2hwNgKo9V94dN5rW3bNM
bvuwnZ6VlAcMzLpOx3nABCkk2owbS9ZCFEW2JKN7FrLOevHkn3uG9BGTjz9vRcnfDbzT65p7SHmP
JcWl+w/nSB3QFW4Xtp6nQhf16eCLPoWaFrdy+bVW/4pV38uvJ4momedfJPmBJRzN3Fiv/Yeny3Lv
5vsOgWH2QZAi7dgNX/TCgn9fD0rl0xI6Q9vbO1DjbWNGOh4ddjvtryBPPiPvkV+FaXxVQx3uQo9a
MXv59+2PT9YntEpmiPHxi/i6xfnmBUE9hiqY2PUPC0rtGBG8WtilZP+qJejA53hWbJI8XevuQlzc
5kbxVtK81biAFAsHeymjQwrjqvEnc5jwQ8R2Q5uYIp0/Av9EiqKdaCEEkvb7YKD1UMSzHVNH9KML
znyMPW9dV1pN5OW63VCe5mIWraLW3T1Gk6NUGAIKVRfj8BNojdxeBlmjHfymFmh6oKENgVGq5Yij
p9FWtvPUDUzSO2mYYbfx3sPPfXyBF+XAjOyORlbno+oRupPYdGGPgSaNCaVJRikuu0Em0EisLk1r
CbdBJUoLnl+UBzhso1FOUezApsuUGZnqt/ioaTRYECVMcem1TI0l+XoJBEll3mtgZUictxk3PDTM
z9KE7h8114BkjkYgy1yQk+SA7yCUn37g6Dv06v68McwEkSjdegSXpHrgtBNYKRjxVcEcgze0KTwc
VaTZ8X8rHZ4ZuMMFvDHzARAznMpUaryEh/3No80h69ezI1cwrvcsRmBvqmBr/KG37N68wZQChvra
eFlGp1LNhysDoydECKOR9D2H0EpjVJJt7E2xSl0rxYx4QdUTT2JCeztvRnuhdtW/N53v8xxs8dPU
P0Xw37sWDWrtdAo8iz81Ef1Sk1MsjucKD8HV52JvKwFby3ZqaZ+f+TMb620VIQyKwhyQ29cF3aIr
O8HAWYwDof1HHd2cz8M520Q52OpUQKwGa/eLkeRtH7/5SjBgF03WnZ1KjGIoM02rH2NQhozsPXzz
zjNMAb/L4xY9d9Uhd0VNyQUYK8t1GngZmDiwn3PURsry3Iv5i9jJZaoYb5Ljq5TyMZ/Qvn9chuJT
wAtLTSFgE/6/Toq7LZcDZuvMdvalHOT8LwRN/BG61CQm97bnaUvV5dMvfgmgV+MV3jAt13Mb2MLv
ph3wShN+uJuVvZEW50UxAyTGqdCVpgHXRkOw8HZZFI4iaYzPvRXRkW+PqEGW3WPGGH4B1wSQW7KR
PH+/KAsUjuR/ds5n+O77Y2PsYJqsL2y0wBXnlkrNU/BhtqZD/vb3gEDwvFMqUkMY55thEM0fWED9
4G3YCiMQivrvkndmG7DPy2t8mfIKisYT3O2M6EGJb7CJcUxOILe+bI+jaU4vK9ZuCwOOJTHhGfs3
LCcvHQkpIqMSuvT8ojHf9od0rSHHw3Wq3W4UaEKMxDaeKoleGp/E/vabGP1oyoHrd1v/GfbR1CHh
j8Fxfk39B8AtH1JXvvNJIWNIqN2ZMvgLXx29tyo01J02vFBmkISyNi6iFsHUFD0bYsg2EMoA/HXG
ENFDDkKVJGr4bGKRzifI68B9i/1NOgRJKy4+gmUU1l8pAX7WhFmos2NvcPGRMyRgf7cvHX4VH4d0
xDJVi76rk5D2zSE0AZWiFnvhICNqUPcqkTDApMng9clUYGeur9+/xLqMMULZLdsYMb9q7SkxDwkD
yb7S4+HdZ7/AXIossLnXhA/yZ7fyEvjsxwa0f2YygRXUb23ksJxcUuiw6mwqN8eewbSHNPsUV2Ee
9ysWGMMaGgfgbCs0HtLOwJWsA5vbTv+AROFSV6tXyFx38x9Ol2WLSOBaxINaVEDjdaWdoONH+lY1
yEFkzFxsrbTrpcppukINgc5se2MSaiexAIBpzDjMt18jBV87KTT2FFTnDtyWpSDMcpqvNjDta5kD
DxvndPw5tJ5K/n5HxHsSENuWF1tJMmvSW+nQORZJUMQQgRoRbNzD8IfVPRcLpQ411vMaAhY1btza
qfRShp130J3Mxn7iLOPRTivdgBXr7L91kPN2OfYkBaefG21opNO2oiYUqh89ibo41e1oy37TM2xU
xJjtGD6gvRF7k+vjpvGwRETE6grFK33DwCLS3XC1iYPWXprYIcPii2SOcuclfgYJBwMUbhTq9K3h
b9V7kXlwj6Us1SIKRPMX7KS39ZdCx4hgsEBUE8U+YnDY+lKzZ2P7Ct6K+MtDkAJu3X3Y0pZibPRD
6tNq6OMOv8jQzHUjRVBeyBcsQyxaNmWT2p4oi3VH6/wDSLdJGi6CDLUmQWfkzlHxdkTXC2WjRxur
ojfGqQ0uJZ5FmKdqbtBP1Rm5XfAd0VSI0XCeLTHsOIrQaStJIzHZbJlYK9xTk0iifKj6WcNYpuv+
LYIqnZXDYTHQw2Ju1085uX+Tf15m1xKQXGjkpTPQjR2PExm2NM/h7tYwH5i1A84PJuDSN60Pofde
BfSnA8cbmnmAcBJZ8darxfayq4jaPWT4kHr38OquPbcVYK+Dlg6lGFxy7GXjNb41jrpAocAIUgSz
6aQB6dEO6exXKMIrq46RldYhLfRPgOXjMdYudQ9AntP6sb2NFNvxsQNVDNEBSvjS9PAtcdwujHIY
x8Hg/dVTbfGQ9DK5ZLtLrZ4uGMTSN4jDAEFUuJxJPvIWF3ZJ5eDnBXzG9EOHHvr97jgoL6tAkrOR
524yFgJwf2YYtxL3mBHZbcStNlso8+Uh2M8xnf2z+ljR5cFT3PxRE6RHfWxrVx3Rnpjl4WRLM023
7Q8w3C3zetheae6tC9bIZgIoRJ92tOzVo40W1oP8d9HD7wEPbZA3peP31c6JJe9XN/5/KazKHszS
h6Nq3lEi3bnN/dcqUnt1X3wjvq9V+AmZ/KVlz8YnOo4pHGJvvpO5Nk085GWjJWISK1c757yb/lEO
izbqxBYoOGa2In86HCWsSJ3WG8tixaSJPLHmZlul9LjRgY4wl83kXOfPzk4U5nlDCam9UKON/P0G
W+ndvgDh2ARQDzGeuUn+Z9hdwJMU32wKaemVzBrLZMc+WZ5R9+l0aQ8UQkQwaf8j9U2CHjD/+T+9
0tMDHnpJyFtf1aibHZDoDtcSeho6OEfSITcf6Ykbnq8hygBAT1b714bhAU6auDRpT/Np++3QrLBR
b3+WjWM8DOvFtIP0mT0/LGgF/mPH4yvzW0wtHaGsMPCsemgY5dKWVb4KDoF5tk6WJl/sWMKzLouJ
AS8RAz7ZJwBnYfY2wpWKivuIFZQ4YKgrvfDkW2R6Dt0e1K63+X9XeMHpCTg6Ex1MVBM5unfXlR+K
zuCSQcB/6bHiNeHAVho5UZgfJY5s4SzihFMCIKN2B5xy9ifdtfSXNUaJp7XSI+DKPHRpmOsn15l3
fBtYOBMY7XnzSLhX2fiDgTDKK7y2j1eenynkKZFg+hFMk+q8TXwfmWKQKtJpdCpmTkR3FkceW8VQ
gz1EZ2DFzjIilIiqefjyPqlxEWwD5DM0E4yBygqX+7ZFaUg0jjVjY9GlTsXxZPuK1PBihyHpQ5gS
fpl9qg3PqteVwrkw/UfxzON0cS8of38L/ycb9374g9QJokYLNaS4htM0cEXdohqcxTm7fQA2ASJu
TAr7737K1r2GwFCp2wcKPWpoi+q/5JHS3KtOHWcBdR/pVzcKw9dbF6dIBpt1DAnG9ZYl5sMLiSGN
nZIKI3dtSSD9usyT5zDgFPyZTfQVFh0Oqpd4Ev00ReFz9ejlnQc2m3Qc5/YWpDk9iPkXofEO7rAa
PCSmTf+M8WfXsVS4RgECD+bGst+0sPG6Id1EiKXHwFu6MIacPjaYgtaDRh1xkoF+XYLGzHep2m3h
KXsXaOU8uWQyo3Qn4s3tBff/HhSsCAeexXN7y2JnzGI9X8RfQRUMwwGb0xwHp6945XwCCwAXChnH
lifhI3upcm6b5jfF/1fVSeUPigLle3j6S+1sjB39dH1p6502BRpMYXjkXT95jhj+Tt/7VUDP20wY
4dGFKrjL8AY7+sfDDGHyyz3reSA5gMIkNTqQ/1Aq9zyCM6N+Hin6KNwVMj1CWEq2obHLH3ZK1A9O
OrVb1g2ycIj8EaHvC/ryxWU5ywubnd6fr5BP0JursJNMyn8CkDbhqp+HMSSrKZrTg+WMJGT7GFH+
oLrwG27qld105NuONdL4W/BFDb9NEj/6zfaR8sK1IwqY7xmkxDRlnPvn7ONyUlIn3UCmziNWqH5w
lwqfJbSqmc+eW00tKqpqYiplX3yxwe6maULpXqFFbPEe2HfSdZ0622LUhZjuJbHxJQG9JDPSy6wf
yiMwhpVFBhyMGO4VSOcdJ449vbIKwFSNkyXmXEqYGZr058n08RIHIdWQc0ws77aFJYRN37bCn4uy
wBFSgxR5Gonk3zKCwXZEcj1oNDA4llkvrtDwhYp3ihx798j6SC8Ifypn0XuvmouY9tGagAHPH7FQ
8jsuI0a1pOXqC9qZ8iEk/0EEg5+gkDDqzaPVJ9997NVZI/OCiPi+jO798Hsoy/r55jgw6kbd+GE3
p51a8d53/y1Goctx3x8cYfiOQyPjVQEXqOK0zXDaM74OMw9s/wviUkf6RH7TlT66Q/4o0Z4Jp5QL
8TXnkLOHovGYyGSNvo4D8pbRL3YAs9ckwEdE55MRQcg/R0K5DIXgNU8YNxNEyzo8JpFAOrX8HJYj
1XqKxV2eJ14WlEJDM0tTIrcfHqJ8IT+8N8hZo7kdr3us7CgG/7h0zE+kUCjE6T+Tds2nhy8KE3IX
41AqQS4CL8FpMKTfHIVFCIHQlUXtVdEvr/KdWaIcgkKkfdkiJ9e91NJcNIxYADRlCRRjHDBlQTAf
4eIuhLiKzXnHcCPtQo/x2Ieup2mgxD2VTwxLWftvYUqYoErJTWm5InZA0qpkV1Z2W49UnqOq6DVL
VF5YANkk7TsJ14Kgum8kjTCJoNGLk4+28IwvlviG10dvzB0O4qqB4pnvyUBetO3K7CNYU1klkmZJ
3W4OcW6r54zeOcPIk+6ia2ZY4jLwX1OCHAZ+DAbVruhQebUTPgpsuK271bBk8UhJq6r2b4Ty5H5o
b4m5v7qx4TRg8ownj381lXYtfzhd8Q+5wWBlw2rXSQ4N1iQjCRfdqL4IOPlkiPO/WJ4iYgfI3N0B
Hlds3IAorNbZUlWr9S41sfNRnaUeX8ZumIyq1qyilQbRGKt2LitzQsgjdMAiC8R4JstrVEiYB6Ve
KzgMkhz5gxZMmknX3DS12uWQD65UvqIAUohVQWt7xHQ/iSSjMOJrFbFjmNUxRnSsCabTHd3aspfv
ez+YI1DiVKdxMXQYRwnH48U1aZVCkJf/6yW9fqU7Zurs9KKEbAqgqB2cX4K6nh2UU10pNdcPafvV
foCqUm4CzyAfADY60J0MgeNj1JGOdrM1vNSD3Kq3iTb0XdueeBibi3LkfxA9T6I9IZ9od94UVPkx
Mt2gjEyJckX17fKiGDL3ojjE10g659xwTDswAX28PVMgkzubVfCtsKi2Es2rXgw2oAh9fdEKEV5j
nO2+0in9ZoG8IgLY74ftcpHBNZZREhcz0KUgeI1JJMG5LBjoE2D4evHDQ30Kej9menn7+VsgL64B
XnbA99jOsO29l23aRPWFunvhtSucZjigWGlga1r6bNOxEUkbYQV9K0nYDgvwokuVqm4AwGIjku7q
rWwJ7l/YwfMWfwgX+Y3rJb+su9Bb1crsTlJzhn6lAppbVlNIg7XDyYxhGihtV0aJai1RtU1v9Lu+
YfpP1WMP5OFDMWHmwSv6aOBKidCS4JvpntIcwMIs2/bD4et+B0KISSlQJnMnvzMRyBoj6ySsQvUV
38N7cx3uNyj6YmeCThO03lf82kuLHo+HqPnmE585HAMwS3Y8mhaNTjLtr9Dntx9PFzaP3hM8ibi0
JJ10AULheRlgZ9N5QehnfYvMBHDs8Od1ZZDXEA0lwEr52X5ZdoooARjZ0NFhSBHebjGwH5uTVJ3a
5+BEY4Xvdwcpo46v1Bv3A/Gu881fvjaoYGJaWVzQJBjOp70d3TrMgX4CNiF/2Z9V0x3J+vAmKcaQ
3ChhSE7gmQnDdrmeq3vprsrOcNNJ4Yh3HBFCx3fI4/OssoTWnEhD+5MAfzSUfmVR1HoaCdlnypcg
Eko/hV/7bZdtbh2dwFrxMUITnASTQa+WcQ64PXgClNrNDTEbE/8BGx86lFw4k7fCTwrCpy0Cj0dA
RBF0Hk4hyScj9V+Oy31NHBMx22mvdf9FQGcNcl3X668n0ISj76t3/tguldnjN/cbpg5OOA/2S4i7
VyniC6x7VTkoBb6qvgk0ztvCtGVlQyxjMCxY7qJ9vbVBpROQf/wao1kXbNJs8uy5sU6U1579hRFz
heUJxwUxLumhUHm9sjyy9ox2HcDuuaneTChsP1e/B5vcY9t+67h1MMsPVEshv6tdnLANKJQY5KPB
O0bajWrky8Nhd+LkoEwlisrAlweXomuoMwb+r6fMy/Rkm0RKwgWj0460nQ5EgDW1FoCzAy22QQLx
8LiiSdZ5pP47HMkVZCBDG3E562bbHOAnGoXusIvll79n4TlQ4gvrujrUyc8bHTvoTNw1rPBx1xRF
wAFNLOJmNHmxoQczyMgDrddYqV7T5RiBSfbhWsPqJl/YYX3cva4NJjN255DY93voAIxvdhdUeOzp
f+IaDoS0BG7xG/ixrE/YudcqEVQxVBFCaNaBxyc4U0Ur1Tbv+vLRMIZr+ay8p52uXRAv4hOtKlyK
LIE3hBWhNoYgIJydOudPtHEBuchxF0rAjVFLO0O16IfyL9/Q/WAfZhsLkh96DYFjikwnVBb5tqGT
BGKeAl0eKPXCf/cLpow8QT+4r5hOErOOzsSu1Zn0nma8MiVakPnyKTvgIayF9m2iEJ5VaHXZQtZO
jTd+V2K5mx7YFVDtCxXIaTJhMxpHgVl2COGWLOBHYNL7UKHSq+q9ZZH9JeTA5G1cV861bmRThcz4
AFoOGu38DLqVM/iNemmf8bYqAOVt46juZ40KoDenTgZts0LIaNUs27KffECwp2mlLE/2/4hQ/nRu
klP4eKjJtnR9dkhKn4OGRwK5n9Pva3vmL6NHVUPc6uvjGG99O2jRHIMUQYgcsvSEvDDVaCIbHxh1
NlLAK3AWKGTVx9Om8fP+m230aPkA5AEylRKa6tUx/y6Wzc5mO+O02JZZvPt89lvP+sM7RcCGkVqI
G7F2yqk8GpG3zMI1Sb1/j2bAj+xu5okJ0rYU8825nxaVDszLkjIXTkReGBV2UVVLDk/0ERaC38F9
YiboPTRUjX66QPLXqQvhnM3Qa2GVJT3WKobPZP9J6JlmfMFsomNPpZ9zq73VXtEfHH5dd8Ott6Vh
HMSOMzUgQ5glQyN4wVejjD+KwJf2GSQau9HNgml9tmOkOjB03JWuMIxIsrWNMDt4osP5Jb6dLwm8
SmgOue17zTsK4HwWdOH3ec++LasK3+JwZKnEDZSpg+FGB2n+QwlC2epHDK++rXM+RLN7+TEAn1Lx
XWjVCLU1EcH/84laWinfny9Hcrj2pzcwZ27vEbWzEzD25PCT0Bm6u3ShzKuLM50lTj4N2lyHGjpJ
BN1g48YudpsoB0pEYNbnd5YExOerQMzfkaSlEWON3sMQVIvsFCItpvpN16POWpTS0JDJi3m/aJ6s
Dajaq85VmXKMPXg4GLidu38RLqnoPIQYuJrTF9n/Azhku3KeKo8XBgxxfqeWVM0L0G0gkvQefJQb
6lroc0Ifs0jG3k685NFAIh1iLr3OVlmo/0mbU2hCntiPtTFDtJJ3qRN1O+MLFgUqMQgOxt/lDhrJ
BCkbywOYwqL20MlfCJewsly3LeqZePcNCFg33HARDStloSiPV7EQtxmEjf4fmtBhDzIfBeOPI3o5
1q5OFQor0R4ofGjwduynp2I+fsAPs8oNafDN94SeBfxUMORRBq4+dQDbsF39vGUgCtB9IyqwFXSW
4vFMtJ5fHqGlm8xAeu8E+j/E/xSuEeC/+Xy4RCizUECcRyahgbpMnoL7WdKveHHM+gSIKSLga18T
KMib0kURsTKCMxaMFqOKn0doTtIV2T7Agm4oHzV+TGxOMLccIvkZxQNM0aVCBUeG21jATcOrLuu5
LwOu/tp0E4Icw41IPIEaQLnPBy4cnGZSJE/hmTt1GMXTGiOOif0FxEUdzLvib8YovUWRYPP0mlry
Rvc9VWwW8JnawOxwJuU5vKVRr+y8VQGmaRDIvz7EFacPS5rhn9qmjGhcAa7Ut/hbbt2EB7dS1LKk
1S1mNivrkOtDnYw9hBjs1bf1b2He69wuS99ji13F98LoDsCjn7wyIFm2gxzcsEihe2DNeEZSdPnV
kiNfQgoyKtT0k/wlbfiaiF67c4aKOiDBMSqgaMwl7bnkzGVohf6Dsejl2REOptz4+LpJmCvfX5wB
d+rW9oLfaaYcUtXU340EPFmBRTA4tlEzMlD6CasyLjwHSot7DW/s27Z9DdoTGRfIG86pMvmpBHU1
NbVEn6Yeeh4skoj0Jw1+B4rwnbiQy5u1ZD/Q5D2VxbOePV8eNyhtzs4EJB0Txcqs4vAHT9EUljB5
YsvK/BfRUGWaTuh7OSAlGVjuBTKjZSafXW8ILBC378MksXeBKseNEPbmW90dKWLvRibkNvz423cJ
4UUF7WWThKZSFriftnhCBujzvlOKjvEaGYQCHAwqhKmzRF5EM5YxhJfiM2t367L3TlDI7Ay6Nm3H
8IG8tfQag7QeIJjC7re3JaZM821UUCJZysy6UPAjfzWHmKGUl5V+2IF3461Nzti1O3nC2XNxHSQ1
F12XkHDSYXIS4X9LycjWMRDadw/hKfmSJXw2XqgrpQH7lDIFhCOo0bWGZZ55eNlXoUMKaX7wHiU+
l3YSU06U2JxEZT+ixVqyfy5Yt5DSWSMonc+6fUYTmwHfrYpcxCTFlgUyogNtOp9QtXwI6dy0CR22
2mwqOjdeDStccGIN0i19i2sqN4yvg9Y5x7hb/zIz55mEcJ9DISErkcX6HdrUN3Eoh9J/wQI2eleX
a9MskCAvXW/AayFI6GTX+Pgs0AwLNgzvj/AlNqaCio+5z4wvM3coB7ZIQofWdIswg4VB18tAmkQR
6KT06ygAkE19x1RWG9+DxVgDPKyW3+N1n1LyUD+hc0T4Hpi8DY+cGXpsh+tTu5gmV5zw31KLK1+k
F5H3kdFsuYo8TB8E+ZD+Zy+Pp94i0c6yWbE2byZlv1+hM11QJBgA4uaGwpXlandMYbo6dh9pdJE/
CB3swr27brKUwq+J4nNz0q6iCL2SjCQpxzIs4LwhNf1YjvPs/Y/9F2IXN1+0bq1YHv4OteoMjFur
tm6bXG9NQVO2odGsVrDtfgnHZOMFtq2IxEpPUmd1adsm3RgSdPqC5QLO0xJt8OUBNXyQwNyx9uGV
6wQt5g+ePMWccITnF9TW5Eim3se1cxEyVgswuyOyxZUR4Zs/jnbPkJmxo9lW4JIU5+Cs/G1MnsTZ
o87pE5tB4NIiM+JkLJddtk//rJawcQRyLsVmAfQEtF0eufd2EHeOsRk2G/uyZy97SApJ5+sBtu9z
hljcymdsTLWjscCPWV9Gjc1NdFfy9Wu+xY7/ZrQFB56gRNB5Hu/2wtFIRP9+dEytMF91YUnQH1wc
NLsyFW9ipT4x64wvS8OinLzzaiBWJS/n5xUAq1MskqG+xNP5GP3IUUgQmVRkekNOSq6SJQAy1F0u
xBMEnGzf4LIxH4HzZ5dcKBP6Ux95odbUXC+eUnf4LNtaO3WNOB9jyCZHp5h791r1DOBpDkKBS9qh
lVlBwN+V+iPzIqE1RtN8xU66lWlaG5U3vYaLqK2wFFx96SIA5B0AweUENrPqEx6v5JrBRv3M4qyH
grGw/ZcDLrBYOp3wAaNfP5HzChyXh1J6H70+6K1e8j0E0TrYJm0j7fTPT4FAe6SfmJyQZxHC2Ds+
s7P9czCsq1FfJk68Oa0K4d0kA1Cz23JHNpK2DprEP4KKr+PKSBUzEgsHNlfho6O7pMeALkzelJ7y
8yHELPSfhTlL7DKO6h0dO0oL4mKPoWsL3K+fVV2InJP2BRBzmLcafDZa41dtfxm0UkiQoaIUcz/k
LJ4RUK1nQOnYxW0Q88uwC4J6EzVMuu3LLQup+547LoW9zwxemyNlZ4oQZ4mmL1UTx+Br/T+sAexD
mh5Z0gEGLMjlB28WxOIxrkxkyHmt6sGSCu+2xv2cwFYknf5adc7jAaGVUvCHc94gjTilpLsIGxzL
9zdv56Uk1dJe7VVY0Ahc9lI+7TsMeMhLlyysWwE+199DiHNg/kulM8cw5fufiL67pQfqR3qX7Mx0
8kCn0ur50EMdSxILbCyaBqawj+5gS7CKMphlRHzT7e6lfbdDDgCsiaI2HDKAbzh3w/gBAZLktrM7
HcT9RA5jbkYKPLmQZ4glBgOn9uqZ1oCmf52r93lA/y3hsdg+j2KfARWPAN6u9ZPE95W2SIv7EfBJ
gcKrzy0ezJ3JF17AaAegTiPMSE+Kccl5J7oRhNdtvONL7tvEMF/EXXBgp2XuO8CDjqj0sep94pcR
dCELkrFcuZHaicz6SUtyPoB4fVyK8CsG9yhRWaDQ4T8WUNttPbmxyAXTPk/OrQY6XEA5uNFlhv+c
vHlwn/PHYPS6FRYuMHItk/MS7pR+z4xuCaxNng5D8lfZT+/33MC6XJ1enagD+45Oif98LeCktJPF
hFaY5R3egAYF4ybozuFHoFwYlgqJXZRHLXp/iv9jIA6NAcFRchlfINjocv40xmNBiR/uZ/apB47X
JxUw5wi61mDiI/fbUacvNC3ueYxGE5Mheag98JsQYCK4DBdjzFUF2B4yueVQa/56iKDAT1PuhqG7
0QdN7YMNju9N5vx69yRDmJ1bBF4aqk4G+b54j4cDDgRY8inNVGIPFO6PFbKyHI4QKNAaDc2Y1qfU
IyZ5S7DsHBgPkuziERJtFZQx/Sg9t/YU2IDqzNys7z/XWJT/LSZFoJrASaKOw6yTg+f0oVTeQjnR
ivKQWLKEJIKLn70UnCK/UozSrQFp2wjPJX2BT9QKKweKt5075PkArSLOUc4eq2wWzQFqaLxO8uhQ
xoRwo0gN0GgNt3gEb5oAlGcHq4zR1fgx14M03foHmmdABzcRE+2MHLESJ5Icz+TnPAO5D4PljFMV
o/s+dDDtlvJ+U2nXIeuXC19xcnNg2V+bbMIQ0qo/k/ZrZbUPv49pLv++hphccV+69X9ZONBwHCUD
P+TOZH7rPHBui7TdeEYGbFPX1NTNfuGHLGYV0GovbWGssBGYsz2EJIkTZKgrHV5d0EFYxnI+SMzJ
UZLCm9qJTKs9L1Vf0ajLkRNOOAYXytMZm9nsSuf6P2pGTWND/lABrI2MQbxgdWINwzpz7gFZXbc8
2enMwUML1BbUdyHJ60mw5DcUp4Gae+0T+f8ClF4wUzTni6CKLezNPmF24zmOHn8ajX2IRZ7kIYUN
VGE4ALI7dWN2+sSgPKEuA+/5icKypAyB5GeBwZ9NHO5tshz6C0Z/ovuOavV799y3fT7XFBTDtuD+
4ne8OpYev06WOeSTselOAcJxKOhkgw4Q1BTAlaDSx7q8mD46YxjCNYpIwhdvuSB2u0I/hwvcnTmE
afX/0Dz/SW2sDIN1mB6AhR0eGOMhqwFWVXdtK1vT6bO1h7quZufg497rTyG96oMCihML8kGavS+3
6i+NeFoh3hTIdRPqP8Wpd8/QteBWijW55ZXIvW+9++jFKUXiTTku0tRktkiWOknTsJhZU3xFEEgk
vAK8kZF3bdYmvB29e2mvobD4d2Z249OieiSkdk8rdl8ppQ7snlNwU0rAZdVZoy9hk6JXxbQSfuCS
Zpy1PfpV/KKpXcW2Pmd/YB9JzBmvVENzPduJrg8oiPZKbfR/FAywOIoWLfxuVoO7T7Ri0d0XKond
5dW8B2IBmVvGRBUHupNYdK6ALvLrPMJz/S3vLwlTT7YdM5OZN2PxB4IB7m+ZajNq4rSXgrGt8ogZ
ln9C6gjZpXidP4lneIkskasiYlYNgTarpBKg3xIUl8RrRrAVG1hua7CdsSkafZUpo26FJ0KBNL+j
qYg1FixjoJ0p8PZxKmlh4YYLZylytIbwsRyCN7z59eiUwdtMzTuIYJ2BGYU4xRmGna3d7h++sQV/
YKYfgkfgMnfCYuG9ncfcLL1WoVKdcdZTGdE7aLzJBeMRA/IESUxs80UtgrHJiBUBQciWqBe+9KVp
2GjapaYtQfvOhoUTq/2x6b/3qqyjm9GpcSRO6peH4kt3/laRsXHWbd6p8wgFFkmumJeZ42VzUhq4
Te1o/zbsAqfdNe38WxS5h9YmCe9/MSe9xMqpz+QRgP6pv8bfFjuXZiflI4/aP/Hzm42TJMiFziJb
hx8pdlRxn4e+i2k1nwggW5LBHozPujmL2qJTWDmzyMoZ3GNYVEgNyYytIMQm6Kd5Ya1hVpZds5GF
EK5GTCsUrTpNzrs3eeug5pZR7tzqxWLCsKOCLCdUZjkVPvlgZje7Qw6LYD/E9juiC5St8zzkpvEq
DB9MmPVL76IlUGdEc9G0va4WMLe06r1nAg+aEyNhSbmauk/GAP2OkT0ZDwOEttPjILo5tWTqCm8D
rCDQux/LtrXqFC/QMZXyLGF9CiWpQA4ZpprAwURfg38ozUTFBxcHxqnqBxhau+kSn2xKKAug7OoU
UO7zrv4Fp9ddE3kTiZE1z9tigL01viVQFvtXNCr6Wcph3kocfJem5ookOmFxbcnBZxOCZOaTeAoL
lz0y6v7WRsI4qT2YXnUh7abgMnY+WwwgWahVVcdk3adM1EeDMRSlXzFmxqI8dr7O5n0gq48c0fPl
G6lD6kkfGHiJ2jz2c5VaNW6jB7fsGhbtS2HTnkipkhHRfdgoB1n4foyucMbZ6J/0AKSJFTzBZZi9
eDdzx5zNCOhW3wtZM+94sbxkqqS5UlRh+UFnnaR3Oh5K3rLRG/Wa+7dO/vROn0GECcGvSY2UYbxI
IZqDYSiRWz6wR9+SWy9Xsrpm/kU+CG3EYX7i8+h7iiobdioTx32k74v2rHo/3RArQJrpHN5ueeMp
OXRRn1Ncbo4GDqotWI1dfdYA2LKgRPF4RNkvxnyTHWF53f42sJBoNEtHrJIj8Dvvp0YZ1lS1Yvmt
qmWgJfxSGcoaTZTR9aHscBbfcR6Bb6y9Oq+9WPxcTnJjwA5rS/bpUh9pyOydUv6alyQsIkxPEHZ1
yuBCprk7lNhFO6GumloBHE2e6L/pNcmmnilp5hlpCGba1x6QvimYxuWwW7g8fiV8RwDBDAvIUEiF
GS2AHJiVsx3QsV11Q5UgFGWGWimvH0ZZOkADsi4nY44NidOm6cGsfP5pM9Mxhhnbnc4N8C1kWGHZ
cb3/LuikdzNl0PNI63BaiT1u4ZqdUQ32HCKZ7pZnEjpHrrexvoY+TW6epil0eLC1H+lFF9a+yW1y
wBVIukchkJXil6PVVBqIWU/TN5KMNtQR5LswA4bR7tVQoari86usfXy5SL+JBlNsSsc/MlNmComK
e+mQAvq22PftbEu4dM23LoTtQ3c58s4fVKpZbAabBxxRaUjUMEGhDgknjp1g6GwSZ5t8DbEpgaxv
N+LV5YqixdLCzGyaFDutyCUNXCdqj1KBmT1xCovdyNdGJ85zmTUctT9wXGuVm7+xdrAjn2ju9BjA
49+Nv49UHIJrFy2GJv8tMyTmuzknBIsZzOHWw8R/lw8hl9Oi/ZhoWmloPYXB2phEHB1w2JLN7qGP
RQjwTyM0i6EPpcfypJ3NCu7iKfHUs0yXI8XSmsiRgPpGEmeD0jz4f7oiFJy7xDNnPzNatkdCtLgk
H02R4zDH4OYMmzm8o/g7Xk37xTnylSPXzIF6x+HkfOM4j2b4BeM8T3Ll8Vb8KLHkc6G4nMptK8Z5
ElNTc6GP9WM+Q2L7gKoe0bmXBNIkXk5l36AvPCNbk3bfBXdvdRZEWsxgpMOa6SOIweJZsnLKYt7e
tZHo6SsDFEmxLMWYCgs/ritCiYeLEm580yDGkEMtHckQOU3kBn99rY5VLJSmVZQj2q2JHuGdnSXt
nvESF1FEFyrmIH31VuhmMIJ2G5Wygp+OhYgDxTbn2hpPLUtgwGQ1Xqb6an+z78WB2egP8rAxZSxZ
ADU1/lus43zRVwztkZhGUN2Z2aWwiB7rGUsoRy/dix6UNkYZVCN2xU9XXiqPj0wtIiTAacsX9QWY
ktkWZAGrajKhvh+Szv8ziyVPrUp6JAckY8oWAUY59dG6ksmMjEP4h8i2uCXo2RUcC3JlFBsIx4V4
TmOWm/Si/SYjY4a4eVvzNK/M3pYtYdDjLEEAdH08ZNoiXeETkFLS8mz604x25rXXtPRQd95a09Dk
Urz3admnrJvdIiOKamnNhQOJQyJE3Tf0tbz2LKNP7AYJJNZrw2lnxmMxNUZyfEmnmI5kTxJjBHNQ
QUcuJ9RBx2rhbmH9QTfkO3k23DATQkJ/wnbcSoO9b0UxIcFPkzriyGDAEDwCzh2cc/PkIbckUhk/
Eyso8HKIA7ftnWHmgTSDb9ex7uXRCUEIVTqlDDWJcN3cHj0eOAcz63we1kflGa49G022MxOgrsWW
5Lo5xCXqTSAc+Spgtat082nc38KriQ52Qp95l+qDBV+vcnOD0vQhll9dcA6SFLcAXysIjVUGmrVF
14gtBtFm9vJTwNSwu5+ftVoYBRql2eM77ra2D0lSYUitg0jN2gwfLCmEtpDlH0qq21YX7u0OPV25
NSBauw48iX4GYJ+n5ogF+bYSOTeW+vOlfUzhIIkykNJHILc3s/hQCpzrmwSauG4XXrCoXUVnLErZ
k4Rz94G2TGUqXz1Y7gPNWmJQAcGLrS/6FBbN0mMqkwYm6gE4UstqCRemyt7ty9RMaoglSYSuI4yb
K4AigY0Tcxoy6XbxJUmdMd/oqzAkkZkimDSALhsW1vKRBd4lEefnB72PfBdvE1uvdxh1nV8yjBa0
ONzFWQk2CGyuUDEnfWJ7epDTYwOxG8dpiGss8hO/2JcYbJjCdrAGmJIc9t+LTKx7MCkvU6nYu1sL
5OPDlgukO/vf5y731t6oN7Mbhbvi0fIDO6HY9IYbcXBvHkKhBb8IYEFBPDCi/21ASrEsnasQD7KU
Utxta4nZBfr0cc6D8CwclXcklzG6jAyxiltWzWrT+AE/TpWVs8175o3lvRtD9F1I/1ZvkjF6mO9N
N/0J1econTAElpssZkjqt/ZrMt01Wtw5gQzJf1xEg0zSTYkND78HVB8WTeAiIJIQiafm+nV6guOP
k7fDpJLHkMrHpWp9vKiTL0jKeh/HP+G0Rcv3ylypr6d0ie/UD8xVwYx29tofsn+FZt9kkO0iH7Qt
s9AVKVMDfgnytvRweH746Xq0SQPfN3C2leDxPhinLHyVLmLZtJ2jVb0j0uB+rG6Y5/2dcKCec1rn
YuAi1RUhQbXje2ts4u+b3wwB1xqgXS8E/HyGWFHk4fJgrUjKJ+TlOPEGi7wFZfBd8b5HU3qDBYLW
Um5HXe24fTf6bL0oauYhndllz9Q8XKzQ+aKSX9ZPIqO62bBEeN6PdZByGIMTCkgaW9s2gsYGn2+c
JODJkZYHbEGOM9RLyrHWRI90MadjoF1IvbskRkb22WPub2nsu0zUYQ/V9IN7Lp7HvY2kh2qbDQko
UIS1YVbe+F6DdnHEbtQ82VDTcF2EUviOp90JxZJ0/u6CVS40lpJDMM8SAjCuEbLYF5tAuEhNL+FB
9VX02TfolrURyzqPu1aC3Rq76gNDYR/+one+M/EA6thbBB36fL3FflsncVDh6aDwokw9tjubUmEL
nv0sCMDt3sj2E+x33MABJl/kyxB7+p3gx1/8z5u3ne6u727nagpSYB33KBbItLjXSkezegFd7hRq
af2G7J3Plt9/TqAHT3tpEZHn2UxDqriEHULKEbmAmIojXNh52V0UvvjQBCYlrgX37s0rxznhv1/B
OSUbnberPCja00LU+RGXOTQyQq1zh3otLHlb9i3n6gffZEWc7J0DH2mBsdxKyefeVMMY5QRNZwkt
vV3i35/OZI77p5fSYHNa+zi5Lc1jkqRzJgQ7vglfIRCBb0e+m9iXBa7bg1X85+sOX5f2LhmCsOtF
m9L6F8rAvrfed/R4aalIAjtoUKj7pjOPACLwbkYqsCuCl4NGpAOQZB6qQC64V4LphO7oPskR4UyS
2WdemgvNw3e1vsMsVwY6rxbXegj3IsAhkuAUj/iTifVfPeG7+9Xb/tVjlCMGpuaGYrd0It+NRtY0
tpnEv48yXMD7ON0WKvrNIwzmm9Sl4/vYuKhd2M8AZdmeY3Xx9aVpUWONwqB1zs5xgjevPVsr6Ndg
BdMali4O6TA5Zjt/4jodn8q0dh02g7fTXSmztWUkw7ItqMaDlgyFrxPw2G5rkVbstS6cwXjMSOGH
cTJr11rKzoUt6oNGgXTUL79AStK/L7lvI/rMQoQ834SLQMnu4E0mm8hV578xleMz+56TRXgVx4kB
6UQ+dxxcyAB0bX9n2ZhHrr4JXwE1bRSSey1U8PIuqfT7gx2BO/MDk5+pbBpswG+wuObGqR1M/z09
ZCy4VquqXptp/uiUu3/tG7GOj67GEn5epu7agi9UzQBt7xO9wQVIfQ0tu7rb5rAjbZlkUHtPIV9d
b+X73LNy+a9V16foAOk2xkdoXzshWjc8HULCnEBpo79cThpEo38/OwcBo54IxVlWu8999/kUJm1q
nS0pLKakP6PjNhBkRwAvuKVPaOzW96DIiy9pDy+vK/KBDeWGZVzsHJAemxIbMsMYd0pkm4/YlJ7o
ELqIENnVpVxehi/3GamM6ew7fONsXRoB890+3mFp0+CzjntOlzV9g11CKHm4Tf89OB2PfghPiluK
In9lCwDEBnRGXc8vxSDsL5csq1FHwL+h4nZl/xSTuPpFyRKegiS3GbVhv0Zj0dYSG0Gmc4b49x5t
N2Tjn2VyIvbOg3hh37vXD8PGeZ+bEn8XpD4xcAhMkhajLot/BvG+dtwRm2JoYzMrNgW5ISSXwt7v
OgQdkcfEsyZiqPRiuzSdhjGtRDN6Hg4M9g4iG9BP0/3je5PYpphNMZIHwoEVv0HQ97rhHtxZba3L
i6wQtqvmM9p56fKBe/5rDTxAWcTmToOfGgR0pXlmGa6/SeEfpYpDDDgvWDQAS9W0zhchmN4/upIW
MPSZT0bU+NFiFxCeCgRw+wIwLOCvo/kWI8PX5LCzAN3ZZi3yL75W3xbcTnM1PN3eprc2nH09acsu
U2sLQLupPdZLr9lG8aLB9gztj+zoeRSRQoTf2LgPen0masluAiAbXDGGP3JuEEgu5CfNjhnr65bP
IQZsR8+oW5pPiJ5/LJje7NHna+Ofuv+Zyg8JSeWfB8OQafyWEoWwmzGuptbtYbxJjxx+oP/urceD
26T1BqRaWIKGxfHrt1S9Z3oM+SMTkqG/2GIlDY4u61xmzhLCDXxtKJS1ha5uie4OfK49MUYSFx5u
OzJ2rn+Ln2js16N1bP012raI/Tdsm2axjULXCvNL+W9ntqkNSaYCvCKC/UrXCj7FAO7PQwhYgg4X
x72pEuM+PGtrc51qJ2AVF2AugmFH/YlIYl9f7MF9SvMjF11uJi3hNlLWoReRhNIPIpGXLDyur1ix
QaBHx23Isq3vwELphmdu0gvqgnhBsUAwrzIxgQhkZopOItHLIIg+7v9kvF/tBxNip57riLbeGEei
49W7wRZEsWmlAYB2SpSRNQP5ucnGmkoh40KlFYsswhN+b/xrf/IsBPKTloJNb8/1diEpuX/lAIKl
g5Apu/4Hcql1W3wzbU4oS8s9TXDpB7+FVGEKsOa25B4hrzhsGYeLXQL5ghCIn3cjJ1mNLu5DoMWu
G+/KhN6xPxnFe70NdDGHf23wwnYFk0p0ZrlhIC7u8YzkBsX9Z0vrjgi1vOsDGDy9LeCDZRCZQqp+
5MFwnU/PPqDEdsrnrkyLWOjDreIr1AcrAGKegsZ8ODHi6O9TtXK++sQ6A4wkk/S8w+sWrbKHzmxf
jAcyIwk4fb+wiCfMu/r2ww4p9nkXq52TX++GG0kqDEucnoqixEFZpRimg5NyCOL8dHGRrTVxbAeS
uNIiVMSIceYOQfF45hvBL7osPD640ljc1yV2StyjbNDZv0bcLrrVZ/7EHAJRFWrT+aKsEcBkTbfI
Jt1o0e9mVzO+tFxJYLMJQ2GYug8whpf6ZqSzTpEkHgjSrhEYhLtHwYucIokWh6RkqRe8VheJzrFp
iqQrT2YdP1RE9QEAadRS8a8FrtFm7y+QAzZyyS+MBDp21yhkSTvtG1OklM4OLJ3CwLgFYG6qzyxi
RPYfhxEPdK9f+Oja5MZY4KkSE6j+Xe5coRI0ZlTqht3Ne1s16thpJHq1AYMRGEUQ23UKbxO1j5sw
y7K/KsOe9zTZzEHdIq2IjW7+LxifIhcfUVO92RZMWzXRFAS37sl9rWmLvVXyZ/bQ9rPbTvXoklkA
F2qPP8IFbLZL7nLcdpuNKaV1QTy04D6/PsXKGqjIT5/hTsyogGueuqDsylN1+1q6Oq/AslaBpi4I
rPrQhoKBe0YkRJYu1wtaacvhi8ODqKJ4K2p1x7SMeMp5O6zCbfHQpl+h1UOdSWV7ntJYzdk5bD3g
7RY0A7dAEmA6N4c/UqvLUbOpoOG3R0blB/JvwXMWPGthVEEEzbaqyipgrzIZ4hk+N+L01f8DZay3
aIlmlKr69md3uiK9aTw5X99FP22XMI+HQGzR1dtENZxz4CO0iOLoblbFKMSIoXSw6KrEB9Av5/3n
CiBTylhH/uJEVKK8UU4Vt1wccZLBW8k4GmDTtKvRqZk7w70hQnbAYMrE3Oy0sdCWM9DtsWveMloO
ZzcO6PgmGmft0cIMVS6v0SnE472lnZlOhKDDCKGJHmcFBwkxPUIoNrFG+7Z2KaGbY6/HbQ4iMPsO
pbKFxsf8yH3MJ53iaH8d6AXTS9uS5hTZCWyx+x0APEWz8sC6CPXkVxBYIs540beCeMOKszXoOapl
89xXbzLEvK92AFrBCcjYzETXHK/8oIN4EERYUGKRX0HhxKXmEW/T2sXBs8QA5ozLzlX02m1iFVq5
sTwOXq6UDnIRornA0R7s2NkgRpl5s7t/te86z2XSFruN6qBXsG80AaNqXLP9OM3k0ZGhE1Z1OrtQ
XxbWiGeB2xgKKOJTVLpngOk5YUaJXf98Mi6FHMDdXuo/tQfjr2d4qlxUAApNFMDBMOzyAU7O5Rhq
cYdFCLXdr0ncnYC/6PUJtZ9GzqYHTtcYJNIqH4iSFBVmhFX1DNDcaBy7R380WZNt0Au96INii/iz
LG5mSbmU4/DrdbfeehrZXGUA5KFMMoQf/cxvHdEajGq8REPXfMzXxcXj1aCOuf2aU0Zv+rYAn1Er
JJI8CChDi1c70zTjPTEWJasCk0U7okvlSIDzxonPTlDz/1FjEQuLkDq8KYW/Ly8IAQthz7xe2pcW
s2xhHBDfNMSBHRyr22aKKfIXl41u1X95WwU+U0IrjH/VVYPOcUVz7Zo7ifiwlAkMs7a1p7rPoHFp
TvTcZTjJyBjta52ozCS+k4lnEZKT/26Sx21nobM086nxPAGAlGVi3YsOe5AlfeYR6qd+aOXiu8Mf
I0t3iv4hwyzSwrBj+cAW8x2QKKGfO7pWVK31Zi0qv+sGffIhazN3/6fS8XCoBATuqSWg0UidY0hK
zXrBpb0UZGZpF/v/XQxDNpMV6Vz49gzHgUXElUz2OPC5WXDJf2QIz8GdnIOo5ltc8XbqfMd4kq/R
tobNFY+omm5vziVjCYwjomIFaZ8NQS5xx+oVdvsTDb4v30HserYhHbeyA4GJmY19slVVUIP5dhmH
rpSQyEjZsNdm91nIgnkFVc/ACDtONFaYyk1UAQ7SgTpgvCo0+hM+aBJM4ZpFCQ91Unwz8f7P9+dE
sK8w9h/540UVJxJ08v1gyvfmvnn5yUOld/Z4d7BLHctyrF7KGSFTxlwWjHSinSfk/upbecOS8/LC
ORuYhL1zWXVIi0HP0ITxJlYmbRcZDI4b8ZAq5pfiypQ2dsEwDC/M0a1iRF95TCAE+vYMEeOSOj63
KqT5F6cKwDt5AxUryjPl0wre11T7JC0tHI1c29Qmsp2840ILIjyoLSKs6/aNsmTpNJXC6sCP7p6q
IyB1jNcVNF0T3qArRxzSl8PXByAc+SqrzLNbE+T43mnm2ro6yaVzuxmc1CJ3O5KUv1JvvHGoAWc1
xxHxILi4g6CEShbbsm1ZAWX/Mhjd2t8YMhqqIpdM3JCW1+2uNTibTjp6DipxE+PeoJbUScnU9RXg
frSLBhbdVHUfskAT4mHr4wy+ZGO/uRezF10sQDJwmGSyzhF4G2uzoIMHyOArbZiUJHx6vthVtBcq
nELGjJ4nimrxXav8VAhZxXKCVR9et34V6wQRC2xduD9BfyIdwCAM+4chfhkLutbc4uBTdr9R33fH
BXEdVIQ02fI/DPObnaCZfE6fNhvPcsXn+7YWOJh9sGLOl5tVoCo9MPvG0/1pItaAL695WiDVG9zc
YlvlvmOMC8nwc+2e4fuB/E3AUl0TUhYz/I3WzL2FXftpZlV4/uFo/nASxN+6XqBDKIJ5qyHYg2j8
gqTvp+XmULUMsmNk5HzIu4g18OgnQsHPBXvhOIhbTI15Bd0wAK9759wbVw1QO4HQQHQxY3KR92BE
uTf5FiZ7DHJ2WW1hcs6XfW5EZkN1++Synt0Y/tHKzuhPyNf3/6vf2LgLVlDAldmxtjQJXakIeqoc
9jQ/M8NxCLBrlk9m1+yKd7iWejV1XAUu9GFYm7NVkaFdUP8e1N27Skx13BEF8EvSZ6k1+dcXNo7Q
ynVKW3Vl5sjOyANWHZBjQfc102vRYXAaAnrRGKFxXacxjhi0xo6SG+MEjSjPlF5O/lNRhDuJa8cH
BAd3h4XO23fZKSGWiE3rRHgDMjm5c30gIexzyoxALqfTMqLlLmSjtNOS+uIQHTNPi9sxfKoYoVM7
hfQSgQ7w8MOTpL187TxqhGuQjJba4HbAEDSQPe+JyovucuMP85R5GQTkbBGIaKGk4Ojm/OyL3+lP
Ai5ayz74SHp3c1Ayt2FkgNFq1i7Sv3S26ft0MWrLdVIXTAIlxsMeBuIRAMTP+ytAObJy/yBcV22R
VK/93N38d8O1JEh7Wb0iaIbwfXnLkHCaTCv0kAmf1mA0jAsEURe5xYgjTYOJGNpuQ29d11DWPZW7
DK/0vLFdT000qBZP3oKd0G0+0BMHkbjY8BLbmFLww9N1dkqJAjXPwgw/r2aF7BJEWWbB4nOz/dwI
Hr84O4NYV74V7x/1DT3iTVdGordRqbWv2M8eamrUUjQIiZ77AOlVup0z7bQBgmuhlckrrLxBNazV
z8rEh3uhf4t1dPaSyYzDCI9pWK1WcqKcV8LCE3GPl6oP0/+u+ZHqL9sbAQEfxiS3L7LyzkWajDNF
xX1Jd6mx0jUvfxoqXPIwJJBF/iHW4GKMcmoJERXKRJvzdHNNfRHhmJC5zBifdgJKS8WzNw2lsExy
gDj+XRj00K5uMMoEeHsiF5951Mr/05gX61JlnV3mcfyl5Xrr4Okafg1dBj+iGWuG8od8NA2U2rfP
r7I6/L+G/U0ZV5aH7Dkd7dZKs/RpvqSx+wv3Ulij9UfICVc0LBbE5dq8zl7iAzixaaeO7R0dlLkm
8VkVjWyOiJYorjNQf8fziw9KSo2BLdEwu1KoBMIbW0igBwOvudm04E0qrVi1rnOenIXwGxOAtJ5o
K9YcGsbf6NeQfQ4i1DBkgteqy70XNFJm/7WjGde7Dwd1MFfRaNxVwjBr9ib7MAirzUsR8iKNrR63
DpQ5U1DhSGD5E7oBz5yTxOxQTajS5J2yR5geamlvJ2htC3YHep+InNDjAIzzHGRwqxdNbcpZ//Qm
tv0Vn3157092nTfwKScCdMB0dG6A5qBEnj54hhPrIYk62DOAFf6KrQoqIK7dBMnyOzo39nohh8tl
KQy4CcN4E/+3cbCHaOq9dd0XeeX1FQ7fhpQTVbfFNkiPbkDu95nSYQelHecd/K6bJZ4rO/5dhpOQ
pB/95dMhS5t4l6gP0Kw/vAIA2OiCbKkTYSXOlbTIGLey+PVmgqIhZo/awjvt/Uc7qCeROHimrCqI
+tOiIZc6Z01JyfsbvAAAf4m2HNT2Jyi5zPmRw7hnCWuQ6gjLNS+A/SEvq3uAn2Mg8JJ5wB++OcZ3
M04IJ1LF544nAfRwPi3wX6EwCJJmQEX8dQMGQyZjt9ePXIVrwB8O6X7adGvXI6cTuTMwXvCCswDY
Sx2MQJinhBafP94UMy/HEPWSTTpzDnAX8FApgwyPPfE0FUqhtyeE+bEZFQUhR0rlGKdB/JC0oJGO
mav2yK61KFkt0xsK6ZBQTL41UtH7HH++s+9Yit98MXTPrDVK/uL6ljjLNZ90gBHt14nCtM65MrTj
URFUBwGOTfQ/WFNkTHHw9ZdG7PXk4joK3OgCBZvyd6p5V7jM+DoRvfVsXPrtECJJ/roLGlzcYP3p
Zpp+9Vo8Twt4varqSpdKgfRfHQdggNAHWN91AO//MTqSneKkc7AOBfZwj3P+0JOh3cKKqjndZ27d
gNai/JCMFIKWzL5f0gPraTX5rCYo0bveDmcUUb4kQe0gP/DJWv6D3zKd09k09f8RPoaozNbmp/57
aVN/fHADYr/8A7s/U9wtyN7nZdlLC0e6ompn/1tyhEauRQJzS59LRDQzPT7gk3lhJkPCuMJnNX5C
54UUgrm9FaCYtzjSthyFr3A1rIZQdy/ao4EQb9niGFv7SxJYh6ZRKEfcnsntEnSZZyeFQCzACnDg
R4dO040bf9qh7iGYQX2KxG9rXZ36UFvXspEqKD0qLn6jUoEnwHldKix0H0aikvPoj6O6xNWDy2rV
D/PQ/Lnj+TcLxi7S/VSpltAfTQx285UyVK73tafsM+amBGnMR3kSXdNq4vdbuCroN5KIl43Qf7sH
z+e2/gBBgSN8L7RsCMQoxWqtH5mzEWuSYO+u/ePrrPupkVRraKMmfGnUVbsv7tKLmZLyNd31T5Pk
HewYoG4bTyzo5xkqcH5hZoUMW17NsXpuUngS0o+EYB/QCjX6fOR1rdESk9swZsFqsSs14MWqHmbx
xUDfvalHwXPxea2TZVAfB0jM/pGNofBBqfj0UkwWYiyt2b802V4Q/zz5xUrIlvNlOJElRH7kLfbj
yHL/VKsMXBCg3krdo54VtxKrFe5FH3qyNwwDRGrQloIGQaZk+/xpG/kPv4wIRdvFrbA0kiRMlqLr
H0igdPdDWIawbqPUgO1yw3NfZhk8vCUzBuVORZidL2unolFo0QFtZRpl1LRvSD8Z2kFwVVze+IBQ
Vt7XUjtvZoQ1daE8MrnCAGyg8P24yf4HK8ifoMwkXA8jkSLpF/xRaUlz0K4wEy6zRH49AvP5n/cF
HIrQqC2mQmVFh2E7WhpG7c6CEzSZ4k9kD3z4kgVLEUxzqYV1H3r3TIeniEBK7faM5VchhHfJc6lr
+FQlBlkuDXyyX8Oamm7T6ohFaeWA1cO2UeOCaAhowkz+2ngwZ3ptXLkZVXVxNsJMKi1CC5e/AVZF
7NgID0SAaVJHDxgrnvKZzN7SFCTy7IWmoWqMz8FTQCY+YCmTWzI53S7NrWc/GjWrtXfDOX74qdQk
mShqbuVo4Kg29F6RPS5OXypuGIUqNiJZ43Im73EMWmVTt+70+YtoEv4AdQiCD9f5r5Jku6SiVEwf
uUPny94b1zd4/VoTpUiXONeNawTFBKmAxvISncwKbGnA3Efhz2wH0iJuVn2saLG7edUVhB4FThnC
nR8k4VbWszhkbWKKhObcsoPzMOK4utDiDNXyKTRI1d5rjhg45yIGIPnhfmNM1v53hOLmdo83NTOO
OoRQ/rHiebjnR+6FD+gzkrMhBGLpy3DHNQ5cme4F7CKzkl1tGtL+rdSCHQo65/YZJy6lwbDl/Zh2
HbZ8dGtsKJrTAU2TvJUUH4muLnJ/EhNqqy2wM+BmvNP2SGuxzzP1Af/lhSSqG8rs4sPwbNq831yt
c7LJVM4cw8HNHgMX6yU/ktuKDe3c0+5umI7ubbFEAZDIg/OvdBx99a9dI8b6jXjkOGDXWwYaN70A
fh1VvwW8qYMlfoLDvnLURCWj+A7RiRE5BJVTIMNI70j5vIEE0wZ078jgbToZwPALzA5rXY76hahp
KB//mxAFlkC84cMfKR0tVRfDfqMvG0ElYYqQkLyxIWkhW6ECz/f5aAGQzy4J4EDm9OuRSPVDACjQ
N9zAFYR2elTF43xNGEduXX5TkqVGb3So0VUZm1DAe6mEYuCUUVSdDtnin8YHmQicH5KvDmAlOD6T
X9ji4SqfwD7bwBJ5WxFOYJQZoMGbS2SKAERhUKa7/XwVSeO8ZQzClkbcbfnshe94pMzbpzrNJrh6
zVvmLjE1577bHJlwize6bLV5N1Dvx94rHKSgoP0ZoxyAVsPK2fsJCZIrKv7/sRjpACUH6qnRn1ws
8fA7KWN8e4F109fp+aF0e5TTHqzBbZcElFbSQ+yxZRs1IW8inPma2tJfxzETOEV2sIfPixLJDaF7
FBOesERsMkqZBw70/Rlm1HOy4x7WnLiPBW0ZI8VTDnZzeH2tlkLcohNLLlboZwf9yn5WZ0taL7a4
x86liiITzI0K/Bh1swpxigTjdfQ5XmuGWS2Crpk4vMPd/GQFH00OXUVGn6mashnhBwXGdkv8r9df
zeJCS4CdVebgPRfvbiZS1NWbf9KZD0znL1qQSQoXl4S+Uc/jqvMhBXVGFP3CAzNLYvGmwqCEfwqU
e3cyWuxOcFuTFNuV1utbEpW1Q1V5+tLSHLpnrhRa8rnXk5Ws/8Q52j+JrU1wNlECWIEpnCe0XYJD
R0WqQ+f61sGrM0Z8CMwTlDo+I0DB3APpKy2lPzBJj6N7M3TixLioObazgv0/QrdrXTrCz01FD+gd
/v+u4Gc0CVOy06gpNasB8faIMSgy071BQc4jGhQq3IH8QaGYuvkUM2Knu2JVg20m0K0UevH2WZ62
k2evEQc//KRt21VAhxCWvcjAm/qOFDXHLuNcqNKW1y+EvJFYFJ+mFO59U/HWOBPRvEIxb5grTB6O
Q+18oibyiX/cMnJFhu8ns910rYLtzSvBzP4aOCVESli3KPmfb1F3eHnSydQfMzGhTBfvTENUNu1x
3beja9P5KbSGIbWXkJzEl2+/ntEFFhL/LAMDCam/+R+lITgZMT1PEziUt6y1e4XrWHLl35SY/YVX
4Aqxod0Ku4PuRO9/dz1dx/WLycxLQ3y1BkZShFeKKpArNKDPUAWWCTt//y+aoae2R4g2glNtr4vb
Qz0b+7Y8W9BhoIZXyeF+AGKiS5azkZbBe3TonLMYejYLCJtTVJQksIauPBtyE3ekjP6wq0iPSlLR
ocvw3X6NUvqrfum42ppKIWLemsaHBzw3Oan5JOr2Sh7yAbV+mySD4BdLR9yGH49x+TsnJEd+Qerc
EiBcq3cUlpMoYh/O71th5lbzPjWFsd34P/tX2DWt/Pm8hbfC1NqiG8HGij0AqxsaH3GH9sfGOHLd
BcndVuh3K1bzlaXaEETJcOFq9Wa4YBiqP5jsrz+A/6HKUctBzIvM7ifH1Xj/CQysA9u/1qQ/T9nI
B2B5t/C1fDMBIdxi9wMu0PFDjtPcc0/jF56IObAV8Ra5OkWYAVNwl1eCCgM6q11OFM40sEn/45eq
lVJxFu1Dbzr91wDzUntjpbt/3VuFCWfXZ6o5A13tisr2hQJk21Kj/i9xB8gNy2rhdM+FziVCBTej
RY42KrQWBeAPR13r6/vR8f/Qg7DpyjLAyILqnwuBoPZqJYGjCJHBFmV2mXj24WVT3fiH66mWavbc
jNFhScjdq6SYn1TU0XoaSxsGbE+FYPVtDCaQl+jinpXsD3jN4hB92EYjuMEadkoR2GxeETNrNQGa
OfiiXdXOYV75XNBhBV7wLc7KfWAh9Hvt2jTWurZek/j4d040b5fbMUKMoxRBGA6oNCJ3G+AKUDk5
MgXBwc2CKCopp15OUbScy3lTLFAiVmGpeusoV7s6VGsv+uU+Ou7WI9TWlf4DMgmtOoYJq7UyMed6
KgXuft8K76+g9DLv4fgk3nFjGj9mGqQCB635+hTf0cIDF8LctmUaiDWtA//xGNI9hvBFd9wWxlyX
rVKDW4FzDLkWf32sPKYpQRwGb7drxDHSoDXhU71dKLjEp5c8S5Ebfldyd4ilsaagn/1XJaAvn4+R
EKZIKFnuvdHttiCHC4jX8nOkYef4+eOf85jthpvF6Mm8C3Uza25kthW2gXqUt5P7xYv475chAyLa
A9064IDclwWrrP7Kp7Ku0X/01y8bWxVCgsDxUIa4eb+mGxsc3U4XiAK8VkE1L5sVs/BCI0zx6EIs
IpOUw4Mb9DJRgqI3sxrYAgpi6owr3s/Aq20WwtPXfLhx1YK1pNpKrNNCsu7B6zS35jaTutzPuaPv
EP/cMBRkX4Fwg05udQuMVrmslz6HFLYcpeH7UVPH0gCKzMTg4YbCpKZB2+1xrAT73HkKDCXJ5QQl
jiOli2+l0hwYk4j5Fgonu0CR23Q3tTCeVFTGKa3nvShVD5vAgLgcDddgNSJshByF5dWhlhmwHjoe
zq90/o5akF/t13oMTFyWv8nzsgKzqHXp1ZhqG5a1+r+yVPYM5/VTUYS2L8Cvz3CaaklVrrGP8MOb
rzlXOjetI25lJgsd/9eVupqh9yFn/9a3zBt4yTiyeOyvRzNnkHZv3HhPCOnwe9mkyW2y9i2ffwW/
2kffWEwBFFy3cEew7Vi1s/BCi2ql3fQB5pTSkr4HaUzz5t09Vym9Hg0ayAp0TC8dtumlGY0MmEnW
zgmhtcuiKEYrP3R2I43jfMOBZGCu4H/he7JCQ+srahEJPBZEuwV5K0sWftlNxiIHLV8hktzg0s9S
BcoNjydobH7b2PV7WYrU0OuCZVVF5aF2aiQCCq9R6TFg06fTHj6VLpfvKFms/NxYrM/s3z3K24sm
LOSD5rYRvWHvxuYpe1sKIyau3bIci1ypYlBunqqUc0jMAwhNbbLu3RDnckizOwlg82BaXks7E7WQ
UDRzL2vhvQqAz1U9X/PAsKRG56NQiVB6YBMsXzz/3L47A2kQYxq5/JkfJyHn4xI1ub3Re8O5QQkx
1csQ9j80Xbj1kyJTY4vGnaEVY/hQUjpBcSN7sKIhAO/radTRdfZwJNY9N2PhsH25V2pANRAlqLPY
nfqj1xEBjvsIJzPFfGa8HQHyqrGzi6PycdFF61WNG1N6c9wX9KQeI3y+vCTqej8yIy0VksFYkDDV
c1MKHagXjKM0riA6INydm0RHdKoWFgAZfCKCW6/PjsJXmyXEAge2M252NiaiX29ni/tl0VvzP6UG
45+4/+QvBeGCXhp75N1KAggbGd1QX5H7vRb9A/VnlNVHp6PxosolnrHqUdatawbGnk9WUGvH47v+
Vs6q2TpFWDkpN6rQOtfWhnv5LEhfG0gQY/qYBsZcYA++ZUYzKcFQS1cOYMbavIXa8KPnx6FJf9/I
ti84mbEtRdOnOA631BMBUbe/M+MYC4ffXwwqqHPio7SKmFEmanM8U5RVRMct0ou7HqiRmwHadane
Jlgl0A82uBepVgIDMKwpJR2sE8Vx7hPiI7yRT7QVGk3QYlLHabASr35+IM7WFU59n0ZjLE0blP38
aWRwSpFZ11tqzkfnaIBniJ+PQxIe1h9Is337yFQskAMe9AlbktqcpRx9GxSrt9aNmxzK9BJq5r0R
moBSdYsmBGOeHnypp8aFeuYHxNOStSe3dBPsUQdhR6Ir+Me25U5bRpUxn2yIU4E6feAspZPRxK5X
IW4YoUv+SWLhhiWx5P6WJqW5Gh6IV1Ac/mdLme5ctHxZR06wrKIaQnN2N/Wo1XWPty34vzrdysBk
gbRKUPGGA8lyfTAkto24DJUvUFU7zFRkz9GakLSeMCqpJ7q8WQ4moilnapGsvfcN2hFAkiX9eWQp
8v05DhjO2h6GVBBE/Bywi3EUK3df8/TQivEop+c06Pmhn+7dRjB86cHR7THtMa4bxDDSmxOk2SHW
Iep4I9gD/mMpFgdeIXoHcv55zjb/XjVdJuvVsclNgR/lkgwl8kGsq1Jgr3PT/WXUWdg8prMhUSWD
7J/Xq55yxma9WK7IdxJT5bWrzCGbA84WTDBzUim+ueATMPIbjA4i28O/4lBhhokCWJdFxVt6ubpU
DNRQqw6twADlMBjGjZObOZm+OI8BlyMYmidfmbb+EUvk8lsRpgZUWYubdZuGJxXjJEBPJZ8c6HIh
j8kHR4KItqQ7ecetTykTv8ZkCpnMQR2cWA1YwrzfACoAv0f63Ost1owoqcDLDiG8GqHwu6ZQLSLC
ByPL1HS/lrO2mW3gSPS1bCBDOzootIGFHoPNNEFO9nHsfvtilSH1gtICFoUIUzMFJbXPHiW+Wx+1
AETX5NCui7kL/HErGawSN4YTbE35goVs9jpVl8ViObvWZRU+/7Plk6F3058NZBJkGZy8GxyNF50E
GdbP5kHQPmCIrRbhl2n9Q/H8rA4GhqDoOMDc2p5SSOKqaKz3toNn1VZR76LQYPAI5hxVGFfStBdf
KgLvDGvh5bk49vE5/dIKcJ7PDxIDWFY0cPxmGgM+HVeRDGwRW9rdTV/ld6+W5VA4OZ91hM000Lj/
3tZlpWXGLbTdaVccv2vtp6CQ1/XhrZKw9VMEudsWirTeD10bjGFyjBbiwEL+gupnQcDVpRugmEW6
0vHCIlIxDXdZU5qIbzcpQAwGe6ybDu8fCTQwKt7rhxd6sC0v7qNWHCSNkKn4kcbGn/ZeIIRXVe7M
jn0aFWIcLjcele3/5rfr5SdUsG8N6SPFCm5afcgqusJjkqk5zcwTyK877r45cJT/2SopCsY9GOD4
+ta7/udDLPdshMZWfuXD97PA7veDcwceRaqQPVKY2VLXN9fjl1QsyKVNsoMm9paNQMSAZz2xVrjO
v0fXZLFt8RRGfeFdsIsqSM4Es1ZcqeW7ZWzjfrBpuQZwWhNF1EuXVgxgHPC53cSBnvuEoTiPQY3m
4VTniCSsulHFD+UwOUnWXOI8aBc2XsGWA+lX0DGj0po3AjDI0rnAn+LECuOesPJMvTj5qtxtV8Xh
V18LysqOzufzvogyj4oOmBejKLxoSnNrP34ShNtfu20WNlUwa9ZJJWFrHkSnjj6po9fpHoBi1BE0
nV6VQ4fNLI7lY6GPT1nraLoStFyJD4p4RdostYm/CC15dV/+0F++n588V9S1J/Igr4m+DS+U8reW
x0hrt4UjD81Cncg9AO8s3yd0zGMsFn3wurJFZQfdGeFanu/MreF7WEJuR5dKmiV0fEfnBKKKtihk
GqWJVw3tO9bTYNm/5aiDwTPnl9ViA70Xowq0DogkIGxEwZuDdIwP+F4UnG6ctEqn/D9ZOpRMoeC4
+ieUpF4eCWf9odu6pWeA4kQMrP3pL6Hw9OnT6GBUzwUaKtYKWiBmdx6yG5OY2h150c2dMYSozn49
hfGbZ0N37QukNLECQ6oCtnsJ8+I4qqZhnhh/3deg1RwlAZ0Qu/97ih5DSxRsS6H4uHyDAuq9flfj
bvMGU3OYvHAi0CIG1c7sePFtSnTuw1MAMoDCu0KNY1xqRw4/QvihHFzva6Siw54wqP3S2RhfHHQ5
IHCRp+lEhBXuL29oIsAeoswqDO5Y6y5/F5jafRvXnOiBXCPv1ugXcfENd4DeIv1hLCZI5HU7K9Ap
RmuoYNMaNDuusrcNMhaGbZAQUnBAKTEEveEm0dySZiXMuDkE35xsEzcoWpVbqYHGKEluXjdg0WXi
BfXyiYT9emC9CZks+yoBklCtMznYvYmgyP4kzXNa+5ToCop9ZZMVbplDNHeEL0HboxJGOiIoCkB/
BQw0YswUsSUzbl4uuD2/lzd5JFM7xnuF1Ss+8hkMBxjjFPnAKyO62qvUfT9TsjGZj4pbFDFxndJm
I228tZOCengUox+Gk1nWmzjz0sbgTb/ba4u8XJo+LdBBRC5goO6PaNsKf6IHiMxbbqjQDuEa6adv
b0GBwKe3T33z0N+BprnN78yllNi9bwPa9joztKdsos15L8jdBFpDmKTiewrS/KZSKcEOMtKTvsxd
ZzXWLjJZDd7qxcd7giunRxsMKTAT9u26QU1OllUwK9EiB00sApMmd++6sT5vwKkm2JzzrP9W32lk
e/+f6BW9FhffxSr0gsUs8idEUGM7vP53EhV9tUlyHkVBH/GeCC0RN1qtQG+8XnR+E0jjtLaEvKVF
aN8+bNT4dBPS2KX+HyJo/G8xubtrwWaD0lLpypzPbct2Sp5Kgudmv7gNKaaTHQuBySkdHHmWk5+b
zkWOvJBr9S/mYeoTBL5mCsu3ygnk22auq4QjZ9PqfPPw3rIwjYg4IjHh+SySLnQE9YxNmJRIusMz
29H+gb1wgi0ddrGm2NXJkVb/dB2+rBh754xHmy8F36M7icGP21A1Ah/ESuDfp5v1MDfao6Qm6BPC
jlrx8XK2D4+HGBJWajwRQuZ+gQWix1npsEypJltbk6Z7zT3KeNbkoGimyc2YwUx19l9tSj/zJxfZ
0IvdObhoy8VjSoJ3BocVYYY4JZWGpA+RFR+XI+mrHvhYxh3iJSQ0npsYjECh0nd7UAZy9dYv8RU6
gpavEgZ22MUrbpvJVHveqC6CBXVkCi9ojUTRR20R3lHPWqXvJd8c1WUEHTcYbY0ZkI/tGFVyrh4b
JtKSZ7Psv5RjZbiLQZGexS/j7tO3fTkhZtb+s/PScgcuXI3ewwJVu62fqsqOXS6xSaS8Qcqfp1/z
08AJOwVNR2bDcqR6DAWWc30aPu2ninB7tbgOm4wSPPtvNSmjETAiLIY68NW5Owu41Z5cz97UCpMG
SfPe/sdrcMQIMnW2R61XHQYapyhLrQ/qFLPPQIVFlE6cEbpKWsTbnlDzoIFF6EPHjUcF7rcjWvBh
gXV1N4v1+YDUC10TSC+IAWNCVv/9yYmO82mdRo5Ub29sZGPS+aTXeB+mGULYTd6NkI37yFyjmk34
+eYVFwkfngyESPQB6py3PFo3Tf9+OSUCCDg9GYkRRWZFFNqEFi6l6sW5+/5yOxBGJkGXKqXg7Qwx
umsfAGXIx4uv4M8xLyiL6BsvBM7CvPpcJ8BEXhIuhJ1w418y5AyQTl77W4a2WqHH1vcVC/bhzhhG
ZEwd7xveEbA0hgptmOgx6sPbvHylQXBVqOOKw7Z52oJ0rD9AyiM/QufwM79zUV1I3oNArMabxaIl
rq+Z6XwwVN80FIDpeD1Q6oaSuvxBHRxS3bgBjFCnj858yV5Xf7gsZA1vfVN7pYLBoHyfb1ZvWW7u
IO6/M+6YMgJO7Fw2Hllg8EhZtaiihmwtd5ntx5AqTg9pE4sI1Nr1jdT0ByX43TJA9LAFCSHIm/gJ
GsPEX7vOX7lGC9aTrJ+HmRVAGEoZR1+rPF2BCXseliIahtfF+Ser/IDekb6DvicebHf7SyqEf18S
iF1zPMlK52dogp5D9X/7uGFTD64dEyMFD5jSATE9qwGH2+oSJy3LHl9aRNrsev4hOq6jKus3NL69
cWRYuUlgJZoM6J0tXJEt1tcmtOMwdw4ZHveiSpg9FksL0j3H+lHatdTfRDhLZ/p54SYkisiCLNKW
JmCgnDo8viP0zYCBd/I+3JmJLEMjHaHLNWPAyKnCFKfN2ByO9S1M3Ej/SqLFu+GldAb53lT1konM
T5yXxPI3L9IxASG7wqdL5b5t7Vs/H7t+u+Pb12s4xxxMLiCs5hQsqTYEZ9QxXwEF0uKfj0s2qlYG
IRjj9DmT5sqkAegEN6Ff+FRsGRHmA0F4O9tVS62ANIBevjr+Fq7S8Q9qGVGDSx/JJiOfX+zfseYq
uAxLE/bpfWMiOKiCTn25j2V22qJWnbaI8GgwcxfXAZoAa+a0jeIQoo7ThYLTH7+mJXH4nq3zcjpa
fK3FUp8A9yD9xx2g1EC/XLZbBjpbtwBf+DVOaOJzaLQpV4SBhGfdG20QVUi6PkiUteKpCjh8y2Ye
NXuoOL5RJ44sgSTrYbS/CP1J4Jmoh+3ctU8W0nJQduq5gq+aVttVwTjPiQVAM4qkD2Wsjq0z5S5E
LsdhL9nFwjtmpRUwl+zzCy6hLC/k5QQahCPrZK7LazGTJijP+J2qZ1Tqeiv3zszvKfyzNzIXSOba
ia0BAHT1YUtf8DqhhueXKdRknOw1i/HQMs16cv7i+z8VMqI17KH8CU58lBep4YYohyA0eWKwLG88
IIfQ6xssXE1iE1J/0w9dMNvHHfWmUEfeD2CUWzbZpMtszo/LnYFfwLCD/OVIeW/hniKY+daRly+/
T1sEhmemQDnkjKEheGtz7+tRX5mve3wdA+A9kRy4w9jIuy+6bdiL08s+m1UkIyco+/tvno+b47DA
rZrY4vdA0a+OAmKz9wqerp8ZWLAmYgqMLZDByT8qNJbbBo92lHVPxorb5DJYAGiaknB+rkpQcMP1
j9cNzt1GupvNeIll0MwEqzUk/sOjRgoYBi+eFlS1Hrb9Dog32Gj7m7UjXWhPvMbK1F0tbktlTiZf
T/5n2Ndp3RT3EHQ4ZCncQDQoA4b66kiAP15+wm0P94fj0KWWnVNRN4LaO+Adrxi5WXxMUkulFWX0
WSj5iRSJ0nEge528zIPlt6a5+K+d23/obR59UBn3ENSynx3JIyvhBHB41tp+tW77dFGCs4VelsWq
7yCzwMZ04TlUBDvHPfVJYcOARSUMc0KJHEeZTE3b5dgTshQatzN53Wa1MJFUTMO9SthgEIkmnbsW
6XA4Qoi5ZPV/nftE5Uhyz16EKiHJrkUGXmfaHZnumzfsmoLtwmYmMc2UY+oRqePsVkqkW5UhRD/y
U7khPwx8Qmx0MFC7iz045YchgyKe5g22TL6LbSUBPEVuGvkfV5Kj9DroHz9HV8zzEq5kc488lHmB
5YIvfHj+cUkztMHRHOwFAR/X6aXN3FS8HPaefsF1WMpqOHC8xtPSm1z4Q1Cw4ZVEAq8b7J0zjGa8
o0oZx6xi3V8wSMbmI/+XZtXM60lvmRc2yyV65f0F3XZRiAVtkiWTBqXiK5XrmhbmYYgfEhHUXobj
PlRVOUHQhyhCkyAQETZV7lC/UlpllaMVXbt04usj8jxuLc4K15mTudnEEE06vhVAm8nQo2AlNReE
6lN8LHNrodery/QFOh2BkiwBmDKOGly1yNpIK0qVUEcYMN7WGib7DILDYX0KJVF6/rcPVgO7bFpz
ZhrwdwKCBBVeq7N9nYCPOvG73YdeycBABj4kUVlZQF3kaB1xu+GwNy4AKqc6epHp1BTMTm2bEjqv
IUouyJGS09HKQ5Kp403F+vRJK+z3St8YjBUhy9std8Ny8Wggkf27t2NW+Roczyj60lKSCg4wedv6
zH27WK5Bq76hrBSS5QOr8oeihIFemr9EvaNSMFXT5HR3HVbEsZUKJ5JDom4SMCOK8y/GCqulTWR3
rA/S37SMXSXFNqIYWwlIBJCZDB3eOfmyzkcXWxwbDVdr7B/hOyH8MAPym5T9cRONA/3LkdxLJP30
/2mfKaWDm6f3avk2F36VPBCeqqngmhXkblB7d86C1PL4O5xWFi5Tg+mrfMcfrqML8km0mCHcpBFa
/oj4jipFjfHVDFaG6pRpbE2ZtC4TaGme1HOeHPOxTUsiGa3PTN28Lu0kSwEtLNW9hrqHQ79DmDAy
Ie59LAMdNRpqgbvW5wwOhAtVdBM0RF57hSMehFbVHk0MAIL27Dml9pfOXy3uDiRJ/K5AOeX+Wpz9
kl4SxjVAk0jhvGXk2eNGTW4PuwW2BfuBd1SrGbXwtP5T7Fyl692F3Rv72Z4YuGsYghWBajN9ZcTK
2rzpKizKZb5rTiJqkL3a1Et8F8pchIuQ5lFrYFdmc3xYz6dHFpsHNo5VsGg8Uz9sn0m4HvmvjdTB
BisOdQVaOwD2PO1u2rHqCo8gDbpdfG38MFwxTYPQ0SgxNCmn5z0vzwmM66lcy0rAiwUkc1dOBwp+
nA0tsU23Nkj11tO+jCNf1t6HbFvzQrA9DnO08TakfMht7nF42sT9kLMQPU1CzYoZxDnyA9HyDJCJ
mNe/6WiQLjzM06OYhox2iAIcYAJ4xcvDYDVtHV54gSbRtpw3gTNyAJj6ijqX5irze+MOUXIEeL/J
/6g1KA1e3BjTlz1mhv1LYTcAma/CsNU/KIfkxkH5hSBWyFNzQrFLhiZATWvmOIEM6r0z+QcR4AT3
b1zpUABTXo7YNPKNckQ6Jz+D05RYldXUQPrh3Pvftwdb7hFPpVO8AdUs6vrEUkqDzGCI6GFnPYlU
pSoZDhYm6wJP2pQIgd1O09+U/TXYAuoODvdSsAR4JdCl60sqfPJLtXCgSbNRl4ugrN78p4OqrLSr
aZiiNRDHzTiRhFtLRLjev58EsZdIbVv1eJQ/7QMfQZS/uHfZ0MjqxcleBJCFpJvHyWR9ZoT5Oyls
bPoZ8v2FWWGZzpWnV/lyDZbZpRwbR/A4QUk5U1wPa8JMUM0/Tbp+TuU9MgVQZHHnsRDizLTiW7M9
hpwgAFWkUdaLUoO9lx+VQGLzcKeUaDIh9EoS2iqADqsrTKyhF4/IHD/wKRI4ylpPHgld+VeDvBJy
+7o7GjudfkUQFO5chMvj21gpO5XR2DPyW0XspXJvc5RgmP55NQ4zgnpkrGxFwQ2ouO108vOo3ln7
wjVkIpwBUlGYGCTUpcqD9nfR62e6b/MRTN2sLLa24Weo5zO59p4x0NvGo6MeqKwMsOQk+o5zCMQG
D5M6x4iSiJsWzdK9GBiYW/Wnufr1RqFtKO1PSR4lm75bKDtqvKtblBBaIosGpbreZ1jJlHxat6Ze
sYB+enTFw54ZcTGUXrFen0yJ6mFP7pX3yvXv0cCvEdr02zcO00IkiOaNFhccPfaBhwI6xQOs8R7+
1ZAcivXsEL06x+hgUpOT/MS8/rAiRbKBlj5HuPC8juKFGs9gVcPTvYoe8wiRHH2QEHGOxC5UnttZ
4qdKJ6oXeZrVzzK5SzR0Ea74KGFmLTfQ03fLDhlq4WHe8ertaaLRYKCmUauHesp2qU6ZPPWYNIHD
u73X0MaGlsu6zARjwJqUCPIE9O7y547RA9S9V+ng1mQqTXUqOf7ftJmryfm++Kbfx6vGHR8mfwuO
XxPyIFj+qpvEsBa6V0G6Qz18NAtwNScx28nZwxT3JBuFnhuYOkZ/cbOYcY4NKhJMr/xF2EVf38LG
Ej9yeLnNv4N6hNuJUVDl+NIJnBMZVV8aHFSTkhsSS73LvefOe5VEbFD3S+7zptKSPEji3PA8+dDu
oAE0MLL3anU8zHRA/yUNO91Bw5Cswov6rAPuRpzqmWzVyYJpB0wNHFZR6O1FsrLqaVi+sGNMkyKy
wj/uHzzP/8RNX7sg2cPOGvppGyps/yN4vIXDHdIy1AUNZHp+NK+domWhyR0822lR+kRWDAFvGND8
VDRNWJwV2I0POb8Cu/vylDOLrQBprfsJsrv2tc0wD3NJLs5/XehI6X0Ft2JyKYkrAdDrjvb9vpLm
9rM3IDN5PZp1QDO2d3dBc73DCdJA444f0si0KOUiCjwi2LW9hJzD/1gkPbGqCyi//oYLBCVLcQoR
MMmSHTTzYx7GrtlSeeNwQbhwNgfO9ptRFb7hRnxlC68sh4JY5SxcBOylN0EMCMvG1fNtZsSkBUgZ
+sXCPSHucug/igk8ulfB35Vm90mLsL9XrSXgy5ZDvpW8A/vP26f8qvLwoRUoxQfg3ZZlNqq42RJy
jgCrzvIJpdThrr80XWh9gAM+9Z1ab1JhN6ESbHSu4IMVzLyBLua3H/1E3o4V0a5kO4qyA0/zRIYy
T56V7/TLz7dyTjxDK5HuySl4tV7Vsp9ExuZj1KqGu/eqMziq3ctjj6ejWvcviYPK6SPWjXrEDBkW
Yz4OqFUvmlUzd8Fvc/HtJV3XajjB2JGGVcQ2Xvl2/Bhm4IKhLtRv9PBzbJXOXhrreZcpdo1p+Z9D
yDW5eyEDx7BZ5iwluqXIHaOvREVfkFMCafEFwCU8nYpFuhT334IHk2GGNUyD/cZPRT8EkJ6zzT0t
Ua0mOMRI67t5eKsQvfIRe4khGIl8I17PHkHdtnjycmxgqcSgZPeFFZeaVTqJHXoqLR5LNvWTIL/J
Db9HAYDWIvVxjwxhmV/aYXIk7Qcuf3Goqmz952XJVdXtNk5ZtHziIYTBCa57dYhwCX82iY5MWlRK
nOuQ3SqYce99eMp1uVfkNQCMeW1BIJasv55mwYEGPuWZUlJgkw6RGI+0Gra/CuA7OPZu78L+VaQd
c4oiyTXbGdR+8enRgsyVAR9iNx6+yt3tWpoy7kKKtAc4Sdkb+BjJ86ZwrqaAiLy5uSIOxaTsItBT
Kagqo9YJxoofZx1s1jQij3WC2oKOKeb+too63a4t804Cl/yFXUwgiB6PgXyNv7DFo1kEXOrNvZ4X
1BsdRt27TicotKNwjNfGd5LJQxBA14FAlpGwWUAsr+vbIEZxmC/vdGsf/KbN3ltAAQw1di8GxcBf
7GKSqma7QNGVOA7o743rrmWVrM95kBcnNilUxOxbSjfqvf/hpqqUGX5XV9S2GcENkzO03hGcZDVZ
xBTRj6JDpiXz/VsdtraIP6wLCQ7I2B3ORx9VDJ2nFds+cTDypuKEu/kJ53cwxjxhm6k7P/2/4N7W
XUPymp5QpsQ0J//yLRIY0H7b1jQ4U9sgReAF+iW2ZrrqI1orzV59t9i/+zqKQx6SUfu4cvN3IXOB
g0sR+gduQd/ynTtRXiGGc/ZOHguhNYLxr3I1cuSaq2EcPVenGL5O42x093e5pLMTFKyGeQ0JTTEI
T3Rd2DWeyUA+bRYN1/Cy17TFbTaPZf08pWNZtGv9eFa0d8I4vhZmII8TugAYENyzmJyg/OpWdUaQ
qSbMG0kQU+69GNrhngCTe02Au0vWdqMMZ8olR9KIAp46V+E00UHG3lPTzJc2/cnjFGt55JrNzHXS
DcprEg8bgs/POjpUx/xBs0NPu4tp4B5PYeoVtHkIhg/caWVwTVZhQUL30uzNAt2hC0SI2s+86v2b
mIzQVb1U3ko9AiYo2c1bn8Z+HoNQo5iARIzdULvlpSlEkqONGs69HzL0fZ1S/d6qPt5jw+zAdwxb
s45VhayOTYZLp2NGV3Tepe+uW4V9ZrasKvkmgWQbgNxPZCykAE/8p9D9r4wTbv3MBN0LSTvdYiSk
dX5ZkSiNdiN5zF3HVubRPa5+pGb5CapnoqzXnHeF5vYVyYtLP0RSxAMJqxfYnIosWpT2hTs+l64J
AwJ8OXqpsbWPrmn5fuTWsHdswx7cqyGae1GikboB6waan/xY27Rci4EbNOpuA4WjWiLVgX+ZDmea
k0PDarQXks7xVZHBY7YjKbSr9x69Dql5gwyJn1Oq5aHNVIlgYqzaQTW5JnBhHWtHmQo4LdRfPqN2
C3OEQ2X0wCeCpPagXZiwMqE20UlYpCcw+46FN7Y1uXAu5IR4qWV3XUXDYLQ8PJb8YEoamyHqygWq
F7JPnt5E8ewM0hxHLKw0s1TBkohL0/IenevyFCuaQI2I8JR80+L9ymldK/ak4iJo2lxevbgBx3We
HgKVtLJZprmqe161xYIbeMv1nQAVgWSKwsAWCNFLH/mjJrnR4S4k5lRBqVb3qYsR/43svjzRFg9b
9JbVxmW0KKbpR+et37o3VVaAY9SjINIujyLB7OG8fpxV0LwaNd6t4qcfBVZULqX8WIxiHK+UAx3s
dDXsQBZOPMtjOQGyPAZqO61N7vViYl9MQ9f+6BKSffNju+gMA3lNnsgeiFUnGmTsCYzNYIfAkWW5
oT5XHJqdU9OwQwzUBRyj4oAVMYkAArJZ7DO1HLFF8Y4K/Hr0JYZmmB057zc8zPtQwC5ztyI5MKqr
7EMH6+n9B3fdR7fvhsdnR3vM/PvgYYFJj0BHs1pDDLGdBDwkNEgnoAKC1B0USIfpQyr4MCP8vkST
X9QdIf9u7HD4yIRS6+PqN5QDgojtkCN3rbbcexglDGVxVRI8HQIsZVVRNdzc6W5fczGVuVFaF1oX
sdVdRbOzaxZDa31q+iuKj10E6xYuiwrvMvH3pCO8xEuAKLbT+pWVjjBVWQyzYelePcKMLx9lY8qJ
aGiLq2Xxp8DZLUZz/eFskY7Wlj6187oqyjyocSQfoW4EAzLSRcfQ8TinsGHH10t0PF4L0GsJLLSl
Vpp1FlT/rmbu5X6w/MNnw6XTmt+ZHWLMCsKAuJYHhyhRboaYnT2mOR0Gd5Viioq6A0zqYOwWALii
emHPaIaeU0oHCVNDpZqXkL204CrQFatfITJnohPhbQc56HBA3oaIquYhOOZt3DYj4gPImtwiAVKO
8W5n3dNqJrZapIeEWdnAuBZ4Vsd1S7eU04mRO40qfnPny2EwaodJY/vs6GE4NtyFXx82FRm2K38k
5ZzPQn/A+9ugGfaRz9LBK6rIQPreOrxCZwiD5TN9e8BSRzXATeAd3SmK8v0hAIqRbWfY77Nm0mbq
HctJiND1MLOURkokK5QULdjfDT2H7acmabnSIdNPBkXwEle6hapaT8r9kVI+euShAV2+EJFwSatl
qTVo8QGmv4ZwJ21icAqziici77JqLCe2bADNKxF4zdXCRfGu/3r/IDeYwZUUqG0SuBn6SMZYP6Fs
B57p+CVd5UF4jjt0tTPZ4oP/V6qBupj/BhJF7OxN/v3fe7hOIYLRoxuQzUQ6E0p6C36egBYHRAQt
mIo5BGL0No5w4eoHQPStvZQ/XNcFUwls9fj3ED/pE9lOrMAney23B3idgG/WDsUYoB7L45pdDgcR
Z0rSlIkzPilCC79D8eKLTAlqEe24ZgJKmPyijuMqvXBf2d7kzuBqalmgWB0iVN16iGaj2USHRyoy
Vnx6b5Q6d7IUPLpskrDGsNEZqSD7j3LbQRsFLcVnqP/pH8c7B/Nokd6wCZPJ+B3wRkH0o1mt4ibP
9wmob2BKN4x0AkqHxS4+9WeGRtmR3qimfMhJrtVCVV95JAxw0i8A6Iq+SDGawSeYXRc0rFU51ZNt
2bNJdVgYRGnfW/Ze+d7Gr6R/H+fM7THFoAKDQhNpqjxFMrsVeSjLjgVYKVtLGGA2HM4OcrvePOI5
uPaYqY++zHCpeTl+hgDaC0rempE6vUgauBvf1fH8dLYujvbG8JPCP3hQauOerP/9gxjhdqBlpCaF
lzGHmQlGvr0Pk+PMoWP+1u97rMN4pt2n+2WExCZY0RikqsPx3lTZgkpLxHli/qDmdSPfkjRMEio0
ZXHKRlVzy784D+5wnPWJtGPfxs/rQomIOWn4xl/tmz3st0rM7jEXCRUkLPeM2bm1eXZXt5LYpt/d
8ipMZO6XA2RhyzglPL4xD3EJbQeQTF5w6GAAVHlxqs76HYUvSvIZB09feUezUWhdMY1JU2bbvaDa
k4GDG2rFW3mdtZaRoxp+nCdm3TMU9+/XU2ufxxKng0SrCGNjK5TxUetNkhOPZTF3wi6K6Xx6CM6l
tAFQg0lDd0z/etnz3Qpu2nOp9WiLIc9RYXjk3SVevs0loZbU/lrg/p9D1Iqw3U5HmWwoq1nADdSD
Ze3jD7snBMNPWB6qkUW/S2UbMACBmUD3yPQNIDwh1dI1xzV3za2cPuBy18k23rlvVHgaak/EKdDt
JnTj6Gkm1p40AvPrfv2TX1VWkJ8CE0Gm6Cw+gcSDJhQTPsEikUpO3xUWmGGz1fuJjYO/y9Tqgw0q
/kJqXZJt3xG5A3IcfoBfJ+DN638J6Tw7JK31+CQ0Hvj9fc6GiLu/9H46MF5vHYRoop38QptGrM9A
15FkrGZKX49uLavaj4XDsghPUbBLJjiL5r6BxvncNfN3DX5viKrk7hq61t3AgkUb0h3LE8+j4jH/
ZYom9+g1mj/H2CmyiAC0MjKfn7mifj5QO4BSTfLivYBgGYGGxYHV8eYSAnEP6CvZ4ZTLGor/zidZ
g7ANuGjv7RGZSXujPK60XOQbARIVv/rGSfAnSpjCtYXM7pVgu0U2MBhUEWc3r2aE032uFAsaQbxN
Dd/dSt1XwkbuW9IznR5xgz+59yqNOF0WQ3LiM7AXrKCElahnfOHBFY7qx8PMsUmDpQAb4ZuYwFCJ
ncG0BtKrP8u9jv6gXLyqvGVC5AaywNJ5snUX8yBpZWW9jsAu/R+csTayhFlUQJmFHj0rm8WZBeP7
s2FrDfv90OHF2v0bCkaM4xaWfVaS3ok8EAJBBObu4iI5FjbCpgs7Fs+C+HT5LgkFl/KYKqFe+3zN
erJXHiADgsgvU2TN5pnwuS0Xg2TOCmSP0C5J9WAxh76k1U9Vt7rNAPh7EYcVsqX0GWcHVCzoaCG5
NBuVAd2A2fe8oP8xg2mGQ4SqxhQwWtOGmafyHTUfDlXP2LPlRnTQQSnjmHq/kzMfh/M92UZQITyl
Np5lAwI4pVE4fjrlkXqZdT0PclesJmiZ7kWlfKo0q0NschQEhv9tRfjoIjzBxUJUtv8AWx54N5EC
KR6LvA7tiQOMOJabYZI4SeuJK1aoEpSVC+SvPP2S59avBJi7couNO0KH5GySv39D6stJ+0G5/HCZ
lQg5kp8vy7l8viCMUo/VlSjcsZXHRjGFKWsNHab72xmcnI60afyQr/H15MMoBiXgyQTbzob/RwD/
jW0z+xXGmYB7AzcOG5+HJMiXH5OYSW61dAj+NpYdA2g2e8sw00Dkm2iBDEhA16VkMJsFw5kq2pdB
myC3GGdd80pxiowcTmr1c5pZQ1vMFnIyKUFgZ8a7ueZSYxFwc7aEr5n5Qnh7j5EcgkTVNVulx3Es
y0h+muOImSK7P76OeyfyPESGCTW78pTd4TjhyL66un6WuQW0PjIWciS2x4m25vup8v1+Bq/cLdsd
XcViQRZ6AUyZrrf2LW7pduh7Uh/tkWnZkiRSYCy73vuRApQFqYUJbNmt3UJL0G5Okp9zQiEzzsgq
Wp8mLrTM1oUrl6vq5SNCHYV+0YV1R26HmE3hxAp92CsWTjeJOMWKoKa/yH9SUgG3ls7bAdv4S/Pr
HMU4Xf/4cPN9W1LxDGpAtcb83CLPzB8OkkanZjd4m17OAmU9Jx1V3zmeBzhGLEb1xLk+lA5cRhGM
CEgcL78LS0OnW+tI0N4Dx5doRmezNl6FI9QnFhPGNqqlwe4cK7+sYmns2JbCDLp7L0sf/EMaWIPL
LJQ+GysLb5LVgEA2myavN/a3UryI92V0neReD3092Zh9LkEJOIsib+ZhT6qSoDfJFqw2WGRPD2LY
bkl5MFZZIUkdtVmGpUk5/vFsqlZgp3xMEA+7DYcPudPUscQ2WIR7orUNRcJtai5810SukXItFRxK
jSksYnBVxSEm6611J7gLGB6U7wGR76rb6jhd7Pc21S94mEvBChfq6dZtxIOL8zRI3ufe+hqPNwXB
Naqz+wn8iLQmcLD9sKQrXikE/6iTCC+ou8nUe0nNF2um04+RUUFEIST9tgDH/+osI+z2SXNGEfWB
k52GIoc9fYo5Wwze7vXaEr+klFBxHpmkJE0vB8b7IGKzkgDJs0+oBFrR4cjme0c+Wze3oOjC8fBi
tkTn42LhAuav8LfEjV5a5H5+eqi84KO3qvTVP6cUT9gsIxhwuUCVw3ehzgSBTfIs7inGmlLj6Q39
g4QBC3k5MENkhno8k8m6JGl5UgaX0OgTyoSVAKYonFonCFUvnJVEoblK/uL9mjelciV+GkQqp/xS
xM/p6xL7NkCOMn0d58XwccAnaHfdRFCFgY9mWkyccei3wPhaYHxHMITLi0JOdOLeN1nIjMZbXx8x
vTmtsFWSvyReL1MdAVIRq4OGlwzEl7cc2v/0SEr9qtSCf0OQyHaeKVrGIF6D5n7lcVROBiE/JZi7
+1cGspsqAW/gD0W6LGQevdeQQuvULmxuYbDYHnSXK6PO035l8/65FOT/DqMhawminp/gluVNwlxm
uoaenPyt6msUYhTf2Ldm9MxeGVvlrqgfBGckt+wak8hNKJM+mvFM9Th9LxIdAyCNo32CGypnxIA2
kQLXE/Nkwy+Kfe+Khptnw4WQrLg2xB7L4RSFPXmRe7P/hQ1N3JSJ0AiUozyusmpp8PkfMdN94B7y
f0JDAHFrHLGWwGLub9EhJSJ+1+0nK0ig2oWcMJHbWsaBhtvpqwzul6VDZ2hZu06MqD8chKQ2V0Dz
Wyedh9JaqdF+IDLHRapQLyqUOOaLAoSazLeC4DBOrfwsf2WmOb9pAOFUWN1lx4arpnuBJhJQ1DpH
GluhQ6NCW0GTOKbXB70HrkE5tkWRI5HSuziEBqV5Oxmpds+lUcSYzrJ4cW5bfoP0zdFX0zaQEI2D
/70BT6h5N8r6f2rLErKND80QWA9g+pi78aAvaBd1sJNMnIdjPajHFIusAOHrS/dHHwTXH9jy2dM1
SIUeSlmKZrYFmtfjR1GxCnf6DubFd5MlWrMzTL57jp4COwg1Jt7FBP4+trhJ0lLSWcusHV1cEna5
1NdgGc9sO4PKJUgDoDA6GS0xFYRYfyK2mx7E3081+lqGd05dwrhApmrCZRdmEpEfP/GirBDs9eex
tOTfayD1Rl11HtxJ5BGDxW4AWVtmsmrHo3z65/hzouFFWMPOLEzrWMwnTiukLbb6QvBSbyUc2Y9y
ash2ykATRMij+zhDY8TL9EbcsA+G/kIbpNi7K/uq7wOLtu8/X1mFZ/63WHePOV6DSt+wyH/RmMej
8d3rFFx8dkfzWTfq0t3BrL6xdCQ7fcpi+zj04CS8//jLhzFmypIhXzvIfA3qBSrQ5UmoxD6WTyWo
6LgyMxLsOW9uLQnGXBKsZ6H0/Hnv55nB2/LqmBR4zWtUG9XYE+1qcjyc4eFBvyElcZ4W9w974eqT
09OZuiGN0o15N3dgZ1gasqE1HRcW1QMYStNN+F/b/iBsfqF41R/juSIiUWrMs34Sj+I8pFKxcjlw
NNAn61wuzsCxU8OlI/4SDt+bnhA4jFjyvqE6NKmb2GyIANJm+E+5Jgt3THndBRqxYWmQHBRnOjGG
Cbiq7NBfDRUbHQdcGLmi3P53tUNkvzV30ru5rUTx8PyJexyOYOuycx0791nUfurHC6bYWkN5RftO
xGMu9bkKtTk4S9RzAGb4iqfBvjikTX3F0ME6M8BJKGaOciFci7NZiJvzO5cznUVqkLR4PApxqWBc
MeIk32cSwlj2LOb50u5YD+5i6SlpP4VxyggdlGZ/iJs8Ce/K8K0DSfmq0nt3fpNr8IMb0wScQJTV
c8SEUwX/Gd8Ct7TnC6HfvZL/HCaBSMdE8wuqy+PxcH8V2cjb+f0IQBUi2Ux0svs39fot28VfGkOW
n35gLozq+ZGA0pZ2f2a9CptoUDJnEWyiZUIvQ3OsmFfX8Uk5EHqb61mArU9xM08BpjkZRtyyfqLH
8DMF+VHKogrevHA6uPIC+rAluYMD+va++T/4P5eoqu+kXpOEiCa7nDurYJDboCi+MpahJc0pH+Re
+hFEiscFDQjEiqgKQDIqvH6UMVYHey7ojtUkjhF4zMz/6giBzrFL4NUMjNwGTpXpZ0H2bCJef9lT
f+KTi0YaisnadSVOTDJW9NiS9gqVYQseIuVQF1wGcobuHymonCJnShtzc+R9WL25H37g6aZ8EBjJ
qjP3DTIYg4288DoADV67ehj4XxOOwLmK65gvORF5PhFGLSIramKCG3MWFYXziHjTkrsH23UZFGXW
FDtWsYTDQo3xtyDxl7sHgx53GObGzFFCW9hOZeodPUjTasQ2e4hvO+lsjNn+Stftr/HA9bm3w6Gu
bewre/kqG5x1y309eSoBjDXLb/jcFGoNUIuPo0uHl20qF2Z9qu1+McjU+zt82m6tI2U7ExCkwLi2
PrqtrrC/6lP9iOUlvGUtrov4uYJuGw9RFkUyHmbV7A01aajhM3kWrVWB748a2oSoqQNptk0NyZPd
xsfzXd+bfoaI1bJM7KrK6jHsKh9aoSTjc3Hv2lrRxgSSbnCPi+Qd6stPqioxps965aRU/HFHNDkw
ZnNJx0odxEurAf0oIIRnCLkm86xxErBVYRmeU+OwxFskfk9sborJTJa2/XfiKw+NLtdiC42l46eb
cHB9vs2WKBcPur2JhAxPYZddV+GXNzksBisDxFbcXD4z16jnZHaRWSBTBJEfhsAH/0JwC4F3T7nC
5kTJ3i0Q+aSFIWH0gGc6HRAamvq3IPkVotr8Q7lYMK7DEfFu/2MY7f+LsAsjQURqkF8M8amp0TzY
JGd1AfzOS6EzhcDBTKcrH34Yq3Suy+p6Wy46nAAuSuvhWSyRJ7MYZIEbY2s4usoygZ09sdgkhHNJ
7xvNQm41FOP5piVb3tFCJiqqW21otY+IeSHbyRmRmLs61CtWMm2iUuCkHgI1011VZoMCjdsadG4J
6prASjX9oU0HSjpaxM3RhjyMx7JBlrt87eSir2cappWoeE4P6ZmhfUzP04LY18eGB+udxrsGJqtd
303WGmvV/QDS480KSQNqEe5gy+OB+gYS/D7VSi5G/QIRwOxN2OBTv3di02GKNiPTSj6L5INGNfvG
MvtxZqbN5EQ8ZesBxNilRvNnNXblqp91EmgECDc7jorIpg6K5bSeWF+GEZviMT+ae2a2JRZWW20z
Eh4VsYmUsTcu8hi2AAcAPTCJPlqq73QGREaM+Vf2dmDtLmnF9cHZ/Ck8rCs5qtz88qbOjc83OPe/
KbMar5XF70Nr2XzumjD4clyKXFrWXsmHnO4cha9Cqyt81K/ag3vifdcoOwpNyb4Usk9bqq67ytNt
tkMFph+yTUWsr/gwOKgJExzeHYW5yFSp0Lr9ByB0odZiwAlLuR+iW1/ItPn7eM4ndfdCzG150Wmd
KVgk409oChYOMuT8iubGnjQ9wFhqS5aqf2ynBgL/XVByr7KlH6uC4qmzTrXtGU2kCwUo+Igs0J35
F2GrG5yAYoVB8G8sGmFNKpWD4RlpuMmV4BSvQKChCo+zPwY/ngfPEGCyO78FQbXo1e4FptX22kzU
4L0bOyPbnoXqaB76NNBUtO2VPvfzcUX77BapLTVIi4v45zTLlx02qC64WspKjqn0u7MOlJ8ynh3K
G5QqEMVsEoyEdBjv50TxASGwD6FGHXHjmFlPDjBz/ALlZA8N7pmF5K9oFJbTFPyc/i1JEDKfLdXV
m/7McWpG+plVNrvt95y18ycdUkfb+fIpiA+AbM5ymJWUCFZoQkkrRyXm+dipYkufRy97zYb8R1qt
LI9taL6sm13Rhxcc+sUox8+5vR1gF1o29iKU0rtSospLhCV8ZLmmy0m9aJvroml8XRwgR4AijDDq
NJh97Y9Dbz08AOF1vb2SH35RMxBlD5VxnEoMKnauHAEQBWn7gqvvOpLXq/0KwTapF6r3pKWHJrpg
6cxPB/p/rKRq4KZfDxIa7v8P7XLvkMoLy+tsQ6fKPTmvWp6DSxcDhqCPzlkiODWMY7AUvYOIqcne
OrlhdSV44ue+YCuBwXTd/CCh3DaVLo1JbDUVX1khNVWW6LBIhjG6QLJt6TuQ9Mujv5v7k31GQ+jm
qAJECVeKKB5IkQ3GXXV48BwDc+G9Hm/sHZkPhGafomwnvEXnI5ztZx0L6M9BfbJMsjinOQ/Qmsbl
KWRH/lUmBi7PaWGa9FhJ20ALLxr4rId56jMoCJMcrR7OkIWfHFZMQ/jzKOTxq1OtGOhs8eIme8f1
SHgIRyNv87gef+NZ4ULeLQk9RGNwE6BA0JTdOCnQa4z55morjE7mJajEHb3aLUjA5NzpHO7+vkkx
miKhrE92QAiZct/dnkHsLMNAjw5aZcGtDSrMABx3OP4ZnTJqEmBF49WNeyZCVG5EGWbLrG+dMy4e
1eYWDLzmO3KZ455zylrJnhqMzq4HDdCbdYQ3dJGbSZlny3bVD48fM1Jd1lsT3ONQ/ogND1DH8spL
rKD9ZYVj8/SdxsIVpGOp9rpnkYTegAOOw/uBbS7wsvMNOnEt2ENX11OBT4V+kFuUqZpsFu0IimJo
Q5FxZVir6VLoNKjwLgXdO1o8cCl/hnVwnq4oTBD/lotwqmytb8xiADRKRcUAY3WUAuSme//7ftU0
FVUxJwXlSNwLRvCxaBiP9LawofYhntyugdSad3zQrfeD0j2WaXlley/Y75ileHtZ4ux+SAbhL8qL
q0kPAtJe1FpOJOYRRpqwPlIkMZXYpog491mJLPBIfjFXK9qk7muGPFV2V11GIZN6edEeFScbrMG0
nr5bxLd1Qqf3feX1+Bn/qDOw0JsY5WYeE2ih9orPDXvqywHnbgWAZNOKXuYxz6vkjvo7PlXsL2mh
Z8M4oeoktC95b+tFyyBrfjwR+X9lrD42392dq/jx2Qw0r0YCjfQ0ckP4ONSbng91yC9hiFmLGc4a
JEwwhySCup2nlyB1teocKJu0XqHJhg07bcc+pCcDVp1wiQw6ZUn/82VAOEr3USD3mRk1WH+wV0Ev
OCHnsn32mcZOmJyBVbiwPP7nmImRR2Y0A1F79hPI/s65WuAQRY0Dq4Da+grnnhvANeFv8SjdnF12
UZcPT2Mq5oB47+vb3GAYq9K/C7uUigVvy952r6zeCf1C1/PtZVPZz+yIZXIZq9mTw4JzFWWDi64a
QkxOXrgbs2SlGVml1MH/x8tddOtcDYxS/x1p6l4FCEwzPsexgdCCVu3vniCqQ4MGaoyv/k6s6OLq
PKW1IwWNUBBMpwD6Qp+JPM4YIpbXXbM5cDcCd+ONLHrCoWyQLazvXdrb1J6mU6Sajq57L135GLvz
PIGbPirR3Qz6EJ1QtI4S0QcpiG3idMqWKh2c3lhrDhboLx3wZWRYr1TWEad7Ty2MRm53h1YXtwKv
g9/47wGSncDJziJAMYa4QLDKScXGKGERzvukpHEtV6dV8lUhJnhm6/sAvl3S8rP2ERFsh3/XthC/
FrJHPi+DN4CSjhw/Z4NE3DLbCRCvpTZO9RWgEw/niUForFW2PNvQeMiR8RLw2W0HhWamZlTZYERk
vdnNvQoY+kkhYSfiW4YWPDjNl6indlqEQADB4fLymdFSGfJoKv2VWFfdMeF9t/KwoNPNkBtHl2ht
2CUxBaryPaXXygFLZuXA28xigBZuNYScembT8etnO1C3IJTp5DsR80a3tEShMSPtp/5RHbRVR98q
Kw16SOqluYzvTxPZDiPQnPJT8bzbZ3HuvF8zf6Sdy7Vdjlv38zzcQpMJUNpFyss0eVPmZZEMZlmn
MSfIZ9D4m0S3alheBaIKMEAhTaZ2jM2PqIGexGjJuhlMNEK6yphkZIpSeV4XuWF7bIRzQ9NDp0Ob
/4wrJWGWIzKv9ZgFnzW73cgCFMrZMyE4m4C8JdJaHnx3YQbiv+v7ezlvAYUowhwLT22F5fOIcFMX
ReRflrJfOVdA9xm86SM6DDj+S4a6svrJZUJh9t5Id0VUrp7At8iE+eAHboLG4PpNTGDmJmv6OOwu
Y7dXo924TEP0Y4Po7RttYi7gWR98MCLHRZOGrHSDy8QTUzXXpzYRp3x8kC+ZNYEhQi4VsmxJIQoj
2LWQYzzDiE7HL76xqkOEX9vgxLiOof0J+ryreVCHNXVULzeq4I6axMw5LNr9U9xeWUkxWQpj8b7I
NKCtNFo3dI5Eg+jhQplatnbjtu5VVXsCOs4VSqslrbJY/ntVAdmZsiX13RDlkVsXd/Ww/c5CSfZn
vTppAkhukOSBxhbdhRLAqJAftYtJkhWVrzKOlNzqbiJNOMOudc8rZZdQP15pn9FZkAgXfWVQdkY9
JfpR9OZxbAN24VHKKxgh7zCp38Ww929WT/YTdLYNgb7WjB5rGWqeul3tBEEFOh3q8J/+lP5AB3oS
+uhQ3RH+PjX9rTs1iVqS4RtB4/R9jqJLXGRSic1vQmfrnKDG2TkxKL/mx49wny+4wlm/KQg3E9zr
OE1e3xwQNR1VFQIYq7eTS5o3r16Vm8brYPwJbBZo9Puasa84dzvlFLdfSP0tmwBwcnOQwrgAvlS3
0YXtkbrsXzXiRRVCo8C0of8y8KTIHpNWx0aST6zHjtSHrge/bVzFat6pXivRGyijzHGwpdhcUYZv
mrJ747UEMyLJapt17lYNuvtXT16rqUNc6ECb263XTNhfu7RieJWboWbcFEoBdDp9g+2PkoxDxeKw
OVU5nj3fgLICkIBMDhPvYwlW0LlEFkzHmMiC6y9evsdcaftIjGC1JSosEWjHamoI+TPo4HFJeWmM
mPiMXRyMez0Vfi/bbqjDvDx44UwtmN4QQkUtTVxXWdJ0OXLu1ZmDPTubmfMHkArsUwcTIHd8w/iL
KlgGBDTb3GtQ3upzaeQPsmiIsNV2WwqxcKl4l5CLdwxmJP3awIURLduD1sWsAQWwEv5FjbyW06nz
30SjOP9Q6mzJWJAehOMH6x9f0+4x6PjU+9xVdjKZrxzRvrvannZIT+n1mnHeW4hrXAwBSyQ3crve
CzTRTDdZUCgDV/hAyYGWbLm3WYxZkmc0pT5OL2Q15XwzS0KLDxbRVv0q8kWvGalbShiNwaEiQq1p
e5GWh/7IMgPwk2GJNZSz7/NYpdIskTbO7ajIFIL53IReAVoMz2Zg2OGzf6Nx9KCWf4kSizFNPVf7
jmXo3LeCJOjLx56vQ3VRIX2YVeGqiSVwIStFcYmU+maz7sCd/6pmFdcTUOPMxzLl8RAAptr0Rt3a
wi+WMpBC08fxGPw+TJcXr+P/PFnfkt5GxrCC6SrH5SByCslI1wZ3X0teXqEK49j4ekdPoesiSQae
rC5xOxOaN/zloOmxtPvZ4GoxBAY4L1b3tdiBEr2l9gLXb9KTKMcKZ8kCFPTJpwqyOrmB9WBCnZcs
KOa/k8A0zt1ljH9SRifFqBDvJpoO45uWZbme0fgd3YlgAEhZy12JFEy1fUsB0uPKQCNjNgxQvWDO
ABK75X2ibRE/UX9Y6S09p0GMbUfl7699FuU6nT9slizyLtBRol5rDFl7r8uZF4WkAYl2GR5h/yuM
sef6nvVSy5tZbp+0xY+zPWxJkYBtvfd5RBF+lHnvK6OeGiVcaeCqIYIB6HCHg6V4PjLOHNVO1xav
RoDsgie85WwxL4ZPQ8QCEie5miF0tH0TVBX31wrmlHw+v3W9YfJ5xsYIOkbu1lTS5Z9MGI2EX3P0
nCLtcor7AEx/vsyReu+XS2F1i7IocQXEd9cdvgpDORLfa1PcbzYXnthypKaHHwKAZUx0sjXfTGnW
i36C2RWideiutTwmQue+mS0b7PYxKTJRiSzhYWE7qVgSiLDXMPd13DHU2MBQWn5eFl0QeWEnmAvG
18W9vXsBUEjTvmRPRSKoXA5fj1btPhXny1YL55IqlNCkknOYDS66jymY3ToDxs6iSh1rrFrwlJui
/0oPv+q8kyWzdWHUpNtuacKN8nUHtknse16EgoB8Q7ou23QachfBrvJ5+FwuAE7aSVhhkEKdQQAt
XJuDcz1t1+BZivH5/gii2Zsw6Tenpazx5TW9pES7KPxmHhZ+4LO7KSlmlq9a5r4keOgCAWpQfV9L
h01WqTnNYhXTmRf+OAcywu8ci678u7xOp+4+VYPMzMUBLfsLP+Z6duyeAmj8z24xp9MgiyEtopts
MMUwzqmAaPcv539EnBbOYAql9eR74w3HpJDjoVdaBdVUR6t/sCp8ZfObdvZLL7zjUAL7KknTNqdW
kPNhb5jMjeJaDff3I91H2anFNrRW+dM9FbcXeO7vtGZYKUNJJu5TCyPNfg7tf/YZTxizfxLBMNHp
qE67CAGs3o/fvKJdvAmFEFPyYoU//ZfYrxEEChh9pavBCpkhol4TG2deaVt23AV3oP/fJTHoIFHJ
M80x/mRK8YJdCScCjVNzUKisXoskRCKg5RvQrYmsMogMuMx8K02AVhYJKKCSCKRUCpE9QNEDidrS
ouE1cX2rJW+lct1WfohdtXu2pNPsWyeLe5a0mFE17bBt9BWLzfQs0TwAS18Y7GOW+MgwA1+0TVL+
rBHp8HWjRWFBFg0MQ/cBIFmI9WR2Xmi6P/vtQIwvPbOnIR/sJRE8A6F0g9TMXYTc9vaSjXnrvtKq
3C0z2DjlRKiwB+i2pBRpd+Oor98zWUjteXoyOjkk+PK3AZlaLXNJ/2SxWWbIj6wSu5vox4P65tlF
DRGeK+uUpDRMvJ6oLmcHHtDOjX13bZZfqnIP7OJsfEj+ny/JpwRC4QV1ijDqhOgawEE7NI2ds2N+
YYvDjbpq0PbMtsUKiMfbHIegz3pP+dR5/7nLkDQDGwoQwk5nrimi2YSWpLdADFmrCbItyPqvDJTM
lN7gXO2SFhmaRR8uo5zwPBsakPS13vTziTRiyCPxI7YWsf4Qq0ksN3psgYX5Ui3b3OHWaFgV5bz3
6rbi0IfnAxzNJxNOgWHzehmdDoDYJ80ianBkJ+3Gd+8DZKkSu1NbWAqoqmtkA6HatYNQ4+gmOxAN
FWBqWmlzV7wToxzlpi4U+P+EOra3fYjYPEmAIcnynqUugPqZ/64fGJ9I3JV4DFeB8EHNGfDRaHQk
cM/ihkwMLC9BtgC+0DLMaGjGoE0o2PbdwVOKCkuymZEl9egXZLR5zdU2lYnf5U6gj+OF2B1cP/Gn
OFxBmLynkc0/dRdt0B9Gs7iZlZhiVdsguL9uKXjxnUgdM5WPFRi6Ec4y4D1tz7sfI7B1Pzf0r7nm
yOol0XEEzvNNo9POufUEpQYjMEGUrAZBoxjx1QmmUxR5uS9o1PACRM5glvOxG331UezMYjST0SH+
5siWRp15XGcAN7gN7aROgRbIt+/f8N4vY01ilHXquo1XKchO39VG9YRgPR0p8MHThcRlpXkgxWi3
hb+4aWR9rG7pGf5QL0MR++zCrZJTVukhXAv/xzubbY8BKadeLD/tItWnFPF3vlk1wIyiqgPy1hqQ
dkSu+gfjkqHIrHvGAS3p1gJycf1YL4J4oCL5zEgoO7hgbbAotxzm6+xWD0e0uKqH3Viai1H8IL91
DLyOjWIVzInaLs262BapOpGpYBXMVAVsIArrERju1v7JA8T5G0cAdLIm5ZXJWa7FvzJwpv0duQKH
NJZMPGtNfbln1uzblzIVrEcnLPjI9zwRqQkWG8GOgvRcaAXstx/52hkJFgqF+N7CQwiSwj+1ujbm
sGhZ8R2PoVNs2LiMXTkCTlaW4JsIv7yWC1vQRmdy0a6ViqbcebvRXvLbAReQclcDRycvfExPtFBs
HHEXgktx9GvfWiYm2uMJFvymD2evfwEZYEyQyqGAT4pR89jcSiGJg5p1n0VFTrHuy2SGACeU+1tY
AZz2kcZaYCK4RSDmfUXcDL6Z1vDIvQE8NH9NIae6L8jFx1AMNjx1d4Z662Lpdj8S0W+31V86N6y7
TZZ/fQzv5KBA7pGKI/0HCq9Kw86FUN5e0Te9j/IDazMHMWhaW3Yilq4agcF5Qnier7ONKHLZh/TX
p74XkN6qQ4NsUUhqnC3rR/Tp3JG2HW7kdFQuD4OJcPXUMRUZnC7ebt41IBBvNKHrSiyj1SKbyIFP
/xPa8LlFriUmeUEl6JT5/dml+4ucTOe1L2aMQx+o0MhT6LRnGVD7bV8hbrCHfetRc1hUPt/ohbEY
YFWj+35BAy+k4KEOSVWwEhn55B/JOvCife/U9e+/Qc5bMO5YQWMfhP0utPqSbOsDrsMWSLW0HBa1
SDDBjr++Lg2GNZCBdsvPV2GMp5FhXz0QZqLgEmpaBUsJf7ebv/+IulAtuq9aB9WNgRhr1jw77I+R
xNNXTJi9RLK3zxyOfTlHb1tQ0XRVcUQlOWFWfDbu5f2CObDrnqN9923i3E0oKCS4AFtM9ACpPfPM
KemBqfMRWds/9W6PHZXCDlJFr5TCDkYL8drAyfqEHUZg6LEsfWYOVUpULwZIxR+p1CDXHjdl0mSZ
3Q+hvGlRK9WKDjbo2WqWQYuT7lEzhe5DzXe85Q/9ZirkMm7d11QXmUk9nEDVs6YuXLA08x/9O5Mo
Oflctl16a5yB1bdi2vA8C9QKxoOYeIsjnDGB8emUzhO1etrqQBugdVQftG+LG0SxDNUCd69bESoG
FsIkRSxC4XPI/LsYi7LRDUw0t+Bwfpp6RgChj+Ys6YOmOKj7JNsOqj4UEqlM5xs6KLo/OitfZQ5M
heCdl98Lvxx1N7C9V/l/aDlXlYRvdBCmuxzs1SW73QikW+Ft10lzm50Er0wYPBS0SjZWhxgL+cgJ
Isq2UOoQDDPOHWBQLL39UIKCopxM2vH7w9smUfecVPZn+7XFywF06Tiq+d4tb5nrtiC4LAQ5Rdjw
TBwXycd3M6OYVAU1i13wXE6MW3lxPsDRxOHid24oj6S89j/nfuP1ZcBrF8SAszUhqaq3uKqd5Kpm
vY/ZvYyvLB2N+rAA2HY/IA/anbSGrECT/6mjTy5ZVE4uNt0Wmrbgt1dcyBPVEkT7+vqpH67kQzvg
IX/99bv0IQo5n620QDnCdYSjHO74R5SAvHG1zZDrGgkF7HdndjyXQ0zzdwyO3Rcx+KhyLlc9SOif
RnxQ3AKD+QNQORgq7kEtKKQX0Qutx818BCt63TjZCtWaWVvzNqoWc6iP8QVaYAsRsaf3n0ySjBw4
1m+T8CFfPrjj871OsoEvtEGa9QrrjRN1MeFI0p/Qpy5IukvDkywiip0z9RGbsDVBQFidd2HMK0J6
UXaoVXh63Pwx+dhVSoke0KkBky+hI6FgWgdGUsCaaRMOwPbU25Q8PWVhZGAhatwLHq7GrQdPfX9z
TiZvFQCFEq1eL4iVfucjgC9CskMgkx7t7RmpkGgsBITLYGTfwxyz5C48WBwJCBqX5G3Pu0XjBNvs
gZG7LZ9hdvsjVROJAVGMryrOSNiXJ6/G3Vp5B7lCSWq1XqGAKV3RX/Fdt6DZyrU07HFOIAuiT+Wc
VxCx1tCN85j34RttXfuroe3DFzCxiIf2iy69Ht09Dnr1MeJOmhLJXZCYcS0jhxuEhxAPFd/aNqUQ
/AD/LlVaVSJhSKJapRKm7IcF5TFBMrotc67up+UnavkDPcQLAVdE+q4zmD2hh3m9pgDMubWOsTp1
P/vfsubCjquESCofjW1QoC8HnZuEE776p9ARGIdUQHJSbn7+5SubdWRDC6sVFHLbPyakPxGza78O
RLkwWE9ppO8nXdItfvApbXZ0j1RcGsZOhUp+QuZxTvbXtAKy06E+e5VypVRjJA4Ebo5SDnIa9k0V
WYaCNb6AYpQ/w+q0OOstcpQhQphVxWCAlOozgxU0AhvvfU2UWoJuJW4UTyPrLldgPdcMz1/Tdr3t
Z2mOcpA7P2924U28Pikaki6YsePOM6xpuq0UP4GOAKT/GHztXHjHgUX8uxhib6KSCILiPW9rA2UD
zDb60ENBXbDobdewvgVN9ct6GDF034CA6UFSONd/qpDP4H4XfADWCTyiHdUkSy+dBzzjSjjLXGbD
Oeko78DRFSY/5ewtCVQT8L6YX+hYcQznb2nPtdd8OWpvCLs6chnY6XEsfOMPbnHEMUjz5lLv6R3U
f2LsqNN+cg2X6jG736pmMhIhYWVL4ScTdUa4k3xbB+g+Af12RX+DOGAxDxpPB0usddKdzOPCBf7B
RCNO8Jpcy6Kwo0ZKwu10OTif67Gvp8N0lSIREFkXWufhtcw0jnvW4YPNdgXoycZOuq7llqdvRH+/
YI0iruREbo3Sz599mP0hIFpbLd8CFWoA+xRyRL6Ik6+gDQYEUAVWWijEwSzBC0+h1a5kO7VGGe3e
5RYuqAuqr6Yrfub0K/eyz6ZFcGAZ261cLuI9AKkLfrbclt9QgcILlbGpNUJKdU9ZrcAT1IFcYcD+
MNNpo7hQ371DuxtALL2hQq2AlUmTxPycuwt4WQoK4zSTsfslvCeDITzDtTLknOLfJ74/zuVxf5vR
EmDD/RSVFxx2CWA2aiOohbWvJkq/LFqPAdTpnpiBCaLD+PFMOusBqB3N0ypIA9RGwz3zYJXy01xf
95HnjAjBM6Qju24v0wF9+Nbnwnep978AbFLeG1gBY+6X4gdf+Qyb1lVUQoTAnyvz9onKNphUjq8f
HafSF2ZrRTiZjEw5yBef9St05gsOJZeI0UU1ssvEiHQxhxJil2Cjbn3EH9VmR6xf8BvDqaK6VjjR
NgThrG3y4wSjdokvkKBN6hIh829l6hkyNTktqySD1/7OSiGb4eV6X6fYRGIyCuEyvMbagOMGzYcX
8oSfPi5jlxfEHG57g7mVJBgCsiHk4NIyLipf610+8wq0TD4tc13SxFlFh1J7pFEPFzDIObTFBilF
goIQChjUf3Yn6IGuDevokHiCOo+nM7R1g0kAGyYvaQvQITtrkkv0gKB31ScfdPsGW0nwSsIXW4kO
8E6DyxcZFOMhsqGMpqXOcWa/44SiBJj4ruF0P1U8WsGBWrsW2FgOmoe8a1pONujnpKDDSs0/WCuG
oAX6ltx7vk3ZP5/mXJ7aivfx14/CF9crDBXumClH/ykXDoMLBUM8LbMH94BtLJVJaLSMLpj2XGt1
EC3AMlBkrk2QszKoH9BpvYMScv3MzQAQpmZNNj7ZDKnfZibN6BV9MRcQR/FCVcz/Gd2uNIJsRk3U
SzmL+Sxe+PPhW8pZwQFqUjdkgfjYkbXUtWW29uOoZJJ5KY1t8/3ek1BsPMSbdQxOPO6XYOYPO9EL
3nmRcSpTuw+A1XwRu53xAIrDza0snL0cotCRc2r8jO42hHpIFOHQgG/V5ejNGWSKBxgJPQ/hD3Nk
OHJ67AA19gOPi3bML5Ei1rxxYVMfUHrBDbzDi24AfsZSR9fE5JRxVgWSCweDEP8RHcNSz30hKvJ6
gbguJb15ZEmivs05Y66S3HAWCnSWF9/76lN5aG5SQzh+Wf5tz6Obi8BDhEHU6K2z1zeg/kGvjuvO
me0+/Bd+73RjFtT/sDvXIG8TyaBleKYQTA9n8uOgrxmbuGNTx4detwJXh14iJdOJxooGf5+2sg4G
/70jFLfG/Kbkvs1JLCY2PTtYIyiQw6VtoLq9hXMlif6LPEqCE0vwRi+Nvm0xfB0j+GlN/wPQa/nk
+vQBRpdTiMr1Whgdug1O9PVq680Wn/LggEqOlayU4p6hsHA3NQGUVUthkTDTD3Lo7n1XACK3BdbQ
5YUpdIipiYFgq+m1bO4zmRCM2Rl8vV8PJSk4K5qjqLe5rsyA/RbrKVzucetMz5Ho5lG5yXa5fpuA
9G1NNPcCY1LyDk0tTqYptX1QNPiTJkaSPq9kGVTNZI9fNn9xWI8TmsgXev4eElMv3fyuYUPQMgtg
ZVsSUs4pGs9PqQOBWq6WOgNG8rKf4ZTeN4L/zXwgc3yM9ROPYwDjMalzzym4AjZFeaJbftXKr5wl
rCXD3X6p+RNIIgx97mJeDaWUEem4N5xlUR3lBsN13o6cvBD8XS07l8FgdAscWywviPwVbJdxJiBo
y2n4X2e3nqY8s8nKewRhA9y0uJAew+wk54Ql0jZOqJSS2jC9hH2p2I4CANCXt3pihZP9MdaID6JI
FBfZoJj3ee7CfFywNbk6gmysD0q9vxZr/Czs+GDoUFyDoau7YfcRIEcsPa+xDuPk83Ha73seUye0
xnGqgQ8JWcxyhG4xf7w/JqbYxOvAMDSqzyq7TeNnBNuF8iou/IKwpuQUTkUp2asVvqjWm59/tBK9
PLWhepsn/dJgO/eB2rHC4537+rzrFfVjpwBLoW+yDZjTBWhK5Mt09YybcjH+2j40vLD5+SymaEi5
JbQluvVE9otqqOAG8+rw3axaFkpvf6k81ghlD2MXVTVWeLliaovQJv9qzJeg4frj50IBhBnS7jJs
kLzk9+N/Lk2lnKYARjGQjvHNoyu3RkFdkY/MnWi3g5w9uYyPGuV0z739/LDNL5ZkaLvtAU+oUSVh
FXeNdvN2b1QUR+WuR6WB6PgIcmCDgwn1lPo7GdYUlV/LN4mkjYVALN+z+NnQGOapZpPsTiKBwLgd
/y2YBTPr180pIMtJ3emVnqyUIvvYoMyCVtaB55CzrguhyOD99ClxJEOdmz/l+u5FShlzED2EeGkP
03DilBznWJPq9hhwXdtae2+IKPQe5wqaL9PikSe88H8Y7RIjKg1Q5Q0gdsAXWACFL0ULfro1dTT9
XeBVr6rvhZ1JMSzxeZYa/niZizjaf3RT7gYW9oKP1m6ok+qpLiVi5KztiRCwJvEURB28EjCvx/Jl
y0x9kWy3aBzayOdGzeZjZeh2QwahZH2AzKizv/LkLDp5iixfPqWk2Co96sl8QOV+lIU1qUBJ9xnn
mFbO1ImVF8PpLawPBDORL53feFPOeDOdCsOLtcSMiCM/1jFhLxF4zQ31enyv47HHUNuRvA42eiBQ
Kk4Mo3tdBEi9pFC+U7M2zF97L9uh3P4e/mH8tMGMnGG10zo1efOBhZm9EJKfMxc+tWLtJqleMJbj
8MxU5ccYjqyJWJ1sG5/HdaHdQwkxUWssvxxbuQ07UX7odLnEM5DB9VfvuEtqhnRZZXeT+2Jrz2na
zgF7hnW4dJ+t3jS25Ou3cwlA1o3soRXI3iWqej9GmYCKVnmqBASMq896VPNWwQvu2zgouZ+3dsFl
j+Q91YWoyMuA8k+fg/PPVxITnsgwG9gD5nIyeqdBpttvf5/+jgyTUA+QqV5Opb4jdgyBXely75l2
gNerG015tu8pIo4Vwe2vWP34SHD8OzRQBGiG7liFPuzOQOaSawPsphz6xAam/dBfHx7gkqhQQjqo
sJpBc4pOKhzPy1dtWT/PN4yJMdqMdcyhiv5tJ3lsVH7XkQ80BoBt6Gn2UzhK0Oozd+9a+rTR2Gva
L2H3wxY5TPDBGF9gPz6tUv+42BnxmGgO1yGDxAybsStX6rCLwCZzO7bldQsLxT3xFLSodD2e4Dhr
hYc/CzfQMyUX5RUxxP+Pm/DwxQk6Q8+C9jEbG4zfd75ZnpQ2grK+w6wi8JhvzVzxsQW44Q1HDSAI
UhYFkiKqQY3RKlFJaNxRINSYfNBSo0wp9M/QxKJeOaLCLQHIGvTWocBR7cuLYaQORSdq85T/Yqqn
5TtL9sOtFuvYPuCzo+GiAl9fUOjJ3D7RuL3KK0pfPRSECjo+xAs8FLrPBupHKnzzoLBnRvC/Bako
o32osAFJaNlIZk6IcK6yGcgR6ZlZLMEPVPKnRc2svr1Dd90F/nHhkqmR9m3HbGhOGwF7oLSJT9w1
SxT5Pu6H+AJXu4Kz+Hy3IZS2MpVQKq7urvrctnpDS3+Zqsdx6ScutHT2QBmXo8v3foN0UvQ3Ng50
M4SPNHfDSO4FRU7g4dFwsQtRu4PM5uLoQ4+uskwL6YG78ABVgUpVTFxzlKKC5vLXBXy8HrO20q2T
JIqzK834ZWMwg2r5BUY4X1Ge+JOC8B1EnQLHmjwq1NsKR8myG9xYkOLXXJTp1kHbNUCjSLIPBzMM
ngsFr2He4mQd9m0HpVFjsa40ARODIEMUlzHyYdb/HY26lY0dir/YA2Fpsw6nLhNZcvQLtb0x3Lel
Cf35spPz8Px6gcMXHt6jsP/yOO73VltJVyFw6rTq5Fwp4OKvU4hWvOH3R3u19sZnnEsEJxCm6z/e
RIbYES9Jn84/+jm2zwFYG/V6e5Gc0RysvkqqQ3xBQJoT3wiXANsrB4bn6VYxdcE5YiBSBZsd2hCD
xoJWYNXIUaNvp9Klcd1BuwvNPl2TYVzqglF9LMYTpUX4Q2JtCsDIRrxzbbQPBQot6lfrjhSDNzGf
4qfD/4DJJYPoll1oe4+CSEXHMS2zSirnOSx1L1GvswXWCJgt6Ko2W853j5Y2KmDJrP8TBHZrJyh7
akiFdOglD70CYRmK6gnu47Sy2m5kERKoqOaGjGlINKHgjcCYrGce0DhJ+Va9OHh3vFLNN6KmLoib
d7paoZKn59sUQADWUt8AIYhV8clKt4k/ARHwCQVQd6F3hg8e7W1RJtvOFgH0FPSt41JXzws0qWF1
84ikRhz+KGXUSuGvb0YZSsbw5xxc/yiqx4et6rwnTlrB9SdsF7HQfokzvhRCwLwmiPGub0TTD2hw
oiIaYrgWqMxFtjgy8ScMxhhIzhSw86vV+s3IGfcgWFMAzB3H8UoAdmkm6A/tXPJ4vbVkJkhBpwbk
HcvT0GPPM1Vg8gyXzsi62vmoAXKaEMSrNzg3dr0Kc+I1r6SJk8mEy1lNtV3N4d9dGnkC5AqQjvVb
rZwgmfj5+mKvDfkG19T5+wne7TXq2ECKMj5AW65MU4/U3JtZjAquobdifCf1lgytPbbFs9cngdzS
X7hz0pXf1zcfyZV/YnN6FvdaOZ4PkhZamcMYQodKRSmvL7fQT1pPnV+6CJgZPto/eAKOv+qZrh/h
3o4o/Yp6JUM/Zz1p6U+lyRC9Udx+skIZcl0MKYqzP2ebARS9I3+0QyhyPLAZ7VYvaC1XMACvdyzC
VfpCxlz+z6V6cRGDfhjIBg6zVhIALwMEX84PFf7lo62cBTgDGBJ0RL9l1W7r+WofyMLbZA2CQcar
eIhuMyDSybtxmZVmhIt13BKPjgjwtjZz2/0YmSWE4bk5W8kXcw6q2JWLFDQ7xxpcczVynKM7spGw
VWYwoCTT/VfPBDnUzgjFLRj2zih26FtDamWcUSZeIjbfjrom8DyIGhHZUoe+QPuiRIT56jwtrfQl
ukOX+WiGH0t9FcmYxKha2hLj0EpSg4JV+unPoE3Q3ZtLzmsze3VzEWdOyQGCzzyUKt3684dtXrrV
sgmFzrliRexmDM4zhXQCeGz8HheD1DnwOgpQXMik+RO8OWRP+CsYIxvDGoG/LxOb7HJ7SmheyyJ0
lGw267Ks7UXzr0VpVa392277hdyOaXg6iC068aRRKmM7CdxTSWjM2eHBoK65Qsp4F0cuQ5OVkCHY
zI2aprBpphAqXh8z/CAbhFOFPLdtIHK3h8ixR1mJQslvP61WcUlFrZNJsGNVY36uQcXCs8iXhBBy
kGWFXbVJdwJqUFaZYlDI2qPu6//ZdBvztU11cfYU/tn30fGeeETkGCO11MkzkoiPh1E6idtUBK2s
DAFVqGqaLKqp3W1v45LEAM/SMjDxIRB5Woke3r4Q8HGemWZWakwkpDYYQ4wcBJjICIlUo4UkdC3X
1xzmCAkYlajkF1aOUoBnuhDUR0sNi+3NWFt/nMICaBnvlPQe4MOI1M/DLNXXIRQj7aOJDbeHlGAy
ABmdsKcZpla3HNiWO8ZaHeP/zZYUYmhBZUKn3ebAM0oYgoPwMb6fUkz34v55v9DLiDgD9waVb5W0
HYZBGnnhebYFUcou7BBbF0Q2CaSA1LS9UAaEv2rmzsbPEGcGba2z+8mvhKYXSMj0pJNy4fcu8hdE
/EyKK72U8q83+9FPZNI3N5wcAvzQ/xiNStcwerTItiUTmIhCassaklIDL2q5/MVlCqDsbM7UyQ+d
CO3GKUyBiqJzD9OKsNFqqRuFQs0ngwq8zPTO0ZDPtQZYtI5vw45Meqaa0DLehJI1aozaTmE4aSj4
/g7Usa+tZ7WXbkgwlnt8Z9ITOdLUgLyBLx4lXbvSmqlJz4hk+yW4dNwTCjEzgYFnG/X/6Gn3bQ82
EK07zptz8FMNLd+fETQffVQrue8DrCeW10u8NKtg0MWaqbo7JDRyXg3igvQQrwCbH/Y4MjKFJfV+
vKZNDZ6sGIK0lSQtsWr0kznLJMxOIq/KiOsh4nYrYb2o1cbb30j7Av3U/147UT6Dqw5O6UApy1Vw
jCep6pSH8RVbOAy3p8xKypAI7SOi8F26osKY9tPjDCdM0ZfdNW+Ih4oHK5o6zDQOLAlvytkmG/Bh
MnFVF1DfBDfuHAKAKY627k2BxWQ9j7vFXA07uYkvs2DikdQAZTQG4Zd0JWmbwpw9RIBX+XV7uXeK
VULywi55VCFYDRQyStR8b0RKiZpvIO+vIfAjzeOc52C4G/TKiC3ka9lBGg8Z+i4lqGLAQbTQfXQD
VRqvwN9+VRZ73QFW1Ar7EEYlBWa24M5KBV/gYrWp04kZAN267c98hafAFipL9ZOjHWBzsUmzainE
NbbOIsN0jPpgi46hwHQ00TX+ohSwXAQ1fDsvV9RlqJyZqBHgBxeQT2E4PRz08Pj1lyfQAOQ0kliA
q8bpjXJziN904aQNefoPPVknSGnNzSrKfjyMDHnorPgOMQHCl0rg3KpUselP1F4IzD8mhvXzjnHu
MuQ46sKKhkw+QeH0Ui1kv3lEmQaf74Obq5F9dPe1osBK7H29hu2PtVWzcq8diCQUxKDogyaXaZVg
9N80PR4p1Wrcpq+L+xarYaE7d1WAsfazF1q7/hCyMDgfOaACOkNP1uifiwaeLuA64pmNLSPovyQ8
QDH8Q6Ghezi22iV4/YZrlm+7ODBhjp6Prf19yA8FlNSYw67bolx/QEruPTETlWGwA3MTCRGReQDz
EYL0L+plsMsyt23HRznGmcncSX1A3DyiDD/7u2LbD77ZAJK37U7tXK58fG09qLXXxl26iQ2RtAHF
uaUe0UrBrbMvij2Ij0LDVQApPVH4kFNfy78LlM9EcThSOfn2CzQutwB9U6RpFQ1Q13+2yOwvrulO
WxxqBfPLTyxw3QgL+Ztut9WHpI8bMnGtQ5xa1fkYNcpmJv3wJuEuDdiW/WO1hl18UHoNXrSXwf47
gsOM9CjueWb6AI9Ct936RPfERLpjKUakZkjiipS8SITjliidzkFCt5XgvBjyBOYDefYVYojAEqNV
LXWcxcd7KtkWqoFb4OuBZToiKih5eiZ2vbp58ZQMIOKPUn+4L/sIIjyKr7JilMjznjZQUSd1ncsx
dLjkWwMAh6VgIPPepuroOhcb6TiCD+bx+AlDnkkPHVCabuGiNv1FdW32aqfGgwASDJ9hRvJwOXqL
w1zj5uu7GRj1nTvRZML9x4ERVTxBH/z/zjSEHE4G/Ww3mCdsduRAV5iVJWtnLav/VIv0l7n9Jqom
cvHHyMDC1kmVIXGLWHAGwIr0a6WoLqFy0mgeV6sDFuQmGngUDQviwp5ogUED/Pa+/CpgeujXjmZT
iW/a/EdMQHrUPOnd4xn/IDp9/oY9zmN4Paca0e5iPe7xqUC+R2Ca4nCaVlb8RFZ0pZqPULwwQOMK
k4BNdZhaaOMk4wRPzaHsTRamu5jGHMXfzP6y6wiPhHnjcY2zEuD8KeZBXyMocEKV25fkbfo6QxSA
+FrZSoBMkWdTV8tN9wOqCXQrvIhrvQqCpkk5jUWW80S6HQ7yFiZyMHtR/NvPD6ZqldrSTLZ7Tp/9
utijjb1gCtf75Xw5TJh7vlfRSENRipcyyOunpSVt932NkV16S71fYv9hZkjl3Uk3NKSZMqNbQXea
Yhiq5F7GY5K3f0bPuY3aYED/kparqb61NebMCi/h0/zMk1v1bifmfa7jZaPGOoXfUdH3S8inq6QD
ooyf24Xqy+cqBvTc6aRd1mGuDXnGa5OkAvot2ueFCwhgICljSbY/M2sYHIKIrRjhznEeKA8Wj0H+
PkI2Ek1Byg49hS2zho4fqDfrqIXCqgDyv9xesxLVebjEojNwF+QMoR9Q72cqi7Wh6Cx+tviwhH9Z
xtkOSfQfEjy+hyTQMW9YWysFEEx7gr7nYNwSpm3wop5TBtrRG+dPXcDV6EvOWuNusbSwf5A2XoZO
xVhKQxjDD0pOdun2sOBnG54SVmkyO05chXudjxbFm1qahDRqDkPMfmktYf/MzYXsUH5HKrcWnirH
4i+dc4vD69iv63w1C6VMgsUKEuJfhp3zIU1fh+wVUDdi4V6NLu6LK/7KopYbWC/mIoJfq84CNOaq
mCZXQSblZVGiuYco5I4pJUWdvhINc2FCE3UDAmi4xleEIMm8WwdJ5V9hrDX/+0O1t/E2AYKw8/ap
Vd/L5r31tj4E0Yn1GpMVL/hGDKvwYADrnoKaPTFawO99FpqtVrzv5oL2z/JOPSizIUVW/A4t6KTl
GU0QJB+/p/TeZoSzybZQ1eHX7GPP+UC2tJUSajLYeFEKU/aN17vfvzRNr+Qc1l0Tba6E0B6ccxxh
YcFI6HQKCjfiYIWeMDutgSqMVpcDCYBqo7Dp1YAhqBr9NLQXT4Dik9aYIwuUHTcJk/DB3v9kFcPM
yOOVfpF9PUyMQDNMIvZZB4HSAxbA+LOkqBdzU2S/Worb/alJbOJztatL3TvY/pkaveSncXCteCOm
aIoZLRR1pMrQBjigjKyAYfnfEr0wVUg34zC6jCiVHG5U7O1SiPZLujbbXo5LPCBRjTrEucI4EV6G
+lU+NWxqfTJ4ebbrYbFQ57j5klyDB6fO0zGT1zARmb583dkCZ4vcnrxQhsELNEveWQH4JHMlKDLV
cy0hLwjb9Hemldz+TgoYCPUcqyGwb2d+72cwHm69RhSx4dWidy66mHwXmqMdBJCRowFWwshxRTsJ
2eUDoBDfRilWZ5z3UXXp/CQGq3qweNHpwZG9QPPwV2XS9AORWxIqqXJHZfYIw2lyRcUULvMhEgnw
Ehy6o4UnNcG1yLAaeeyqPBaeYlDpDXpu6y3sWItYJE9vjn5ZsuHOLhivBJbZa68UKp/f0fKIVw8b
3GiTYzgpHhMXAZFQEpMFd5GQd2vH98Qu7CnDIezVzbY6x0bXM7K99950yqtfO17QNyfoDF520b0N
MQ3DQzDmPLQe16MFkXDOq/4jjSyacH9KvlxkEBib54/sTVuYVvDtP8XQl+7GmsVWTDJxdR8Y/3cP
mP6Hwb+g7f6OEtUXwwqzTqZh0C57aXl0ac5T3UJ9PdtrsvZajKwWUwftPnxUUTWJdS5xixTEq0VT
wpnliEYc1ii6mXf1qkOcsMp436fXCdNQk3fMGqQWF+coMGXm8O7iHXgUAwXNpK6rn3hOZZcqn111
4i9ELbhIeoLwEcfoIjiFYAosWIfgYNXFpLl7RDR9P4vxQhLvw8Mc5xgE2N1Y9QZ1WM69Q62PdWjk
NEuOhWIIUQPB4qyEieCBpHcWLwD3OxUATmueK1l+zlo8o2KDq0WDFMIkD24i2VWqV1S4LBRwgD9x
NyDBd+sgSoKgL+8qM/2sxRSD0e6mTVLRzdK9GEx0n2SK3fXqA+nmVWxYAMEz9RHrU8RLFZqw5pKf
taVq4lKRY64MYShTzfxy2gRlO4OboCK1R4AcjRxJ48Jybj8vcOp2I1JLG1WHKSW+7RT1efH5peSH
Gz66oAi1F8BRd+AYZMO4lwfKbSPmooH9HQlv5yJUgBsrXXKg8LmnM+SR514Ep7onGuXdRwBFslvA
giCU5qftgLqPu6VBJNr0ccIhl8dIVacj9OQloK+AdP7k4CtcGFSPOW0SNrcWU6Dir6xtTECd2e6x
jR6dIbti4tiq04v/18ZtfemB8chUfVP5dPZJzYr5zGEp6vmbdbThttt6G9SjRiceG7qB7OaMknAk
iGNwHI1sKah7v64MlzITX2iAwlqR+3aRJYrEboufLRlib8D6sLHP5t61KwZxFs+nKf9Q7fB2NMhD
L0amfIaMflrbQ5SYyC9jqebYOBRXy0VUeJpS7mXUrOIiJE8GkF5qZGSOVn1X1nh3hzbSoBAzVaqc
L/VXxqrU/qMSW0es7UXgI8YpOsAiNeyhHfCFXOmUbgVLPC2tylkLIVgQgAKCwRdfi3BMS6bjymDO
xGAjUnZQdm60nm5z3vLUb+t6YodclbP3fIPToM3+U079dbu/8uYWIWPCZfupIjOxClFdk0WbP1rj
1eEy34sIrCKZKXd1w8EppLK5r7UXqMZd2z+ACY6aNxbKw8wMffzxBX7bMj8MAXTIb3PFSuf9nR3K
3hddzRrH9VyQFJ0XKNxI3j+Nsm6CXvSWtJhZRvm9jXyyFz3GoLdHrPA2YKVTJnKXLb32qL6W1+Fc
KyjHcUZY0SwaEwbQ4tARit7TGxNsVHcMI1xB3+c/UDsHcyeuHbOchWwDhLtSUZfGlkGWZobtqwMF
Agh1ZE4X1qgRgftSMXZzVUcffOfP1TvWuG96d3Xr4JUAcsjSvLND+UbZmMaruRwHuQzoA79fzdpc
gb9kNIsChNFpFft5R10eN7w1qWVmBi7dxXZb00i/ewDN6ZB+WLmE0emjnMj51BtIrW4Q+jXNBca7
Vod3hLLk/YNGoGtXwIlirNkm7ocnU1d/BA6KKaWWq8ctWNS+OdSwycBYAa/dM4RnvAg5K1DWcKcF
TgoEyeg7
`protect end_protected

