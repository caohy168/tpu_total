

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
grYpUA5jzoYp1LlWmdZ2ALEfyb0iZaBlbu2Jn5TWbislv0ePefGNtLrxAsy9+neVRtGKqzd/weQY
1GDOlCD3sw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jJRJFGl+freuRUOkHi4uiJXF1ZSDXCZnSp7sify5hay8gI8WQ5QHE0Kl1tU1VRdOD+ovbKr3K+cS
UqWpgUyeIHMS2fFsOi6SAu6Aoshxr0Vl9PE57JGCyWYxhIS/bFj42inspCVQCybe04fBzJMNWaUp
2qePZYRz32xbymT2jPo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu6th/stm+M5ynB/TKpquW8ZkolQD8eNSgYHhWrx1S0Oj+qDq3ifkyYP979H5aZBSsmi9nhkBeP5
00SMQNL9WZH3DTym/hO1AOEB/vZQ4iH5QuRFIKccEqDq2JtY6+UDXXKzO/1rIfmarsHX8ltlRTV/
zcfaeOmCAj7ywQc9UqYmky4qV8fErTo0+Sdz/lesSXUkxz2bi3RdkWlaTaVx6gglEIQd+UT3ZYt3
+UGswd7jIOxS6vlCnneyc3neS690RMPIIoNUnxysnaeZZUGvdfZpjktfag6rjQ59uaAGWliO4MMi
6ToA8bqievgo9dlWIHZ7qHH63+ZPGm4+ACmZLw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
anxX3tP+OSA4f+Zz3xRPWpNr0NFYOEkjWa+yDywi9ewNNEKmVmuybI2vuUNyxHHqdZuNWtw1fzH+
LvHMudDHSvrqUXO0i+yPr/b1uULww82dKZJhMTouZXfSBUYYR2R6eOUHlkc2mpuJW1b0Yfgqe/lL
U2cURbnRhzUDfX4a8/KZsget317eHUxMWntDUJjMnFKpxAe6rTs57ljr+47CKoyVApxpFRtXyva0
iIrl61ypfwevW1NM+dbuq0A2ep4qpKF3QXqu+5quZRKiS9wqmBIWbGIwWUFzi9jVuDlWbiy7K2/8
HWrhgAyLQfd3aizqZge9Kid8TFg/tOAzl3/Dig==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hfg0jhNUSwZoyKs+dkGwZfuOuLOYxt8dUSYFBsXNe53zJQUTW2+PTKtB4x0Xb2iLN7gmIGI0MkTa
VnwntAtFN20kw1KSsvMMJ5tmSswwrxvHJwEQEUQ97ZGqSWO2GHL6Y1M+TGniM4GhJ4MqrJ9nz3bJ
lDbNWHgjFGsf/h3qT5IiPslEewuncdt89+9yjAvcmXEyKAI2nU9sb2+Z/dYcbWohVAJhqZIShNET
j4MueDXbjuGAb3rviJH30Ms0ITe492AtvNh8bbtTcCumEGRwdxdBrBtudooM4fhp1QOulK1MlV70
8clOJrGF2872zCxai4LigCCBOk0uSW3ObDKbXg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SbPUQ56CmxNuuFeULNmdtP4VI25yIuTqRpQZv4fdI4ab2e9QChHgoTeL8pKVO9WcuhlNTx166GsZ
+J7LQgSi3dQSR++PcS3u1e//zfZcwXePmh5ndXtuNKSeOT1YlsZMy0NFnCR74oDcXIAWozlvfa3H
+Ha8zpAYNJlEcIxIlN8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iBM86j8TSZyV5DU0rYA8Io0mzpNhxgzW55YqzBpIYOLzQUiY8G8WAdKhnnqwoz2tPjopVirg1TR5
tvZKebOq9UC6KFo7vKxpOX57N0cp4fFPLdWGp3bfCI0YVxBdZnmmB4Oc+YtxYdI6e+BC82GkMG6d
gVuqFuf9L0mulL+yXuTTt2uiDajwZIcjyq11UByNJFKgZWndCJNV+FkUL21qP0t0BgzJPx1vq9GI
Xcdhwmaqi5DH7ZSxtXWYHzXgMDV5w1iNgDI3RX7uYUR/uvXUFc8tvCukL4SxyVDekPuhO3EOq7lP
gm4n/MB66m+/WkJd04R1OsrCyFsGEkoFVCl47w==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TDm/CaHzF2sRlkHDDHosS/V53FzLYAEPesCrg1+oRNDDuRD9Xb5WpyqcNNNidE9joaps4c7lrYCD
3nRf5x+Z12x0YPF7kaiPnyDbXkFRv6Qy+JTaRUXeoTs54W+jPqxDrL1x6Wv9yIyFxShptBbnNkVI
e+UMuxDyxwcdq81KmTCZc+NgWtBB1VzY7ity43L6Zk/6njjEpAsUd275HuhcP4JW4NFW1TZDaNnF
Cww6OTyrgEG5hWZR86AzBS7yjfi5vJjN94IDbGHICM+1BbHZNAAylzDKaXvbNdWIsQbt3lRVnU+z
u9i9+X1Drqb7MWsOo8jYLXDlib7Gpm56+SqMOg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133696)
`protect data_block
S99ty30j7ef9ZYqPlMy9sjqAxM2ne3URVH/Gb36B/jp/WJVcbn6bKNCaClWCoxF7YcTY7mF0TyDi
7QcYMBd3kUjs9lYJdKOS1Yz32ps0UyVi5nipC6LDI3PlDfBDp7r8SfooZo5I2y8U0t9eixCVSVsx
hzTyO94kT7Ruy+li1sCSvFvffhirNGt2pEQQx7gsZ1zvLv91+lDxNHllkPUGn9sfiuCR16I8IM7t
CU+bXKOYiQIcchNwjwLSvhCXHAwp347H3FAXE8POJn6iC/RZZXzFpy5dbEe1r6ambqoQ2Dwi7IeA
+zRAXNJkHVilfaOrJMtw1jGfOLH2UhBarBgru+qB5CDrOh0xWnmbG7klXpZT7IpsDpftLtT/Gh6Y
+9u/4iX7fAwXA4XwzNPuFiyfPx+Rck2NTy+67XGCsKPMljxDv192svNGv16aXZNpNxdx/gfdSvOo
O50lMIQ2KE5YKR6w4Lr8kxTu4JyBcps3vNvAEqesYFvYmk/WTWWjCI1EQA3SKxSvTEuF3BFkNmFb
wyDgoOcq7UEAxw5v34/eGJNqo4sHi0jpFgHp8eBBxGv0e+4RaPrXjF7w6+pbWRUkMBzR4ZTLv3bI
XrCM4De+MUw4WxwFgTiOFPvvSmGi0rhx44wrDWkHaWIr2mcXEk3gn8ZfMh95LFctP/+SdFRx7isR
X2OW34BrshUwafZn6I1FLxmEgF3kYdJHdhRGe0B81lorSG1fVAHBmUdmpBMmuGdAIKl6JGCWbhLI
2qbNQtZQwPAlQx/oCe/ZHq2e6J9/6mHJvbdAdc/PrXqu6Xu/7VWAISvcZtI8tan79onud5tgMs8a
hhgBV7TGaSfrCn+JCpqWCHyv3476wkkSdJkbdXpWfgHG/aqszogSzBCp1dxCRGnQTUoVVfDx2Ism
13oV7D+pQLfFDqiJJwYFeD7xE1Ru6h86CY4C7t533dKNckJkZPUg5k9Xwm4Zr9iTVrbdYzEyJNnV
SI2k/LBBSKqtXoE+qbE9schteLDvGwU8Ikplw71b98H6VudgQQNOvwAsCIHy2CuTMtHiiWjbYbpO
Ce/R+EI+Kix7gqeaNSzIjBvmjIkvL+1YRIDxK6gRGlBnl+qVH8i2LbCKaGk9zufNFvpaWYbJ/hCV
246U2awQXo4qx7UomszfFCT18t7JaGeRxeji73cVjF3l8AXGaqnEV0dhPuTBunp2SfBsXRYSvL66
eHRe8dxeOaWZpbAYOMX6QURIeEE+rpiA+P+D7drYXXWckprod1MXDonnqgatv81nnDrQWCPYAjzG
+wd4YMw7xCKjHTknZC30VUA0bTJpz89rPllx++sk4okPoDH/6CzzQplTVQsphk0/7yatlSF5YS+c
sol/U00bgqwss853kGhMLII4nJP6uR9wu10t/wdVTGJ/UmqNOQibjXb5IvCcgKtm338sAf1bs8y6
oSLb2O10bqfkOg+Y9QTMx35uHRbtyop8IQoJ0LU5g4d+Wk1igqacf1fJbL7d6XsnanNeggkCIX8k
uRtBKur3TcjYbAtSy4T5/MWmX/H2FBZuWlirIpdKmnnbZF5Ahq571Nw+c9fmKDdRTwAgIjNRjkHh
Gf3JfPFoj7eaxI6/J+65TxcOjGcjzHnKHWfd2HGCNZwqyM/8K7dWnOCBLCImDxuGg0qKwxO9BWQ2
5RZEOyt4jg6FM/BZvr3hP1mWhbXgIIfFyxdGUndJxaSBy/rMzytvF3xdbNAR2XQDEcR3vCISbTcv
q62TsI/8m5R8DBAcyvaUROG5zizZASonUmMOaF5P1g9054GIIFeusYYl/yHumrHuBd31GsFIIaHX
+BCmq15snVJlqMlPtgtTrEA++d+FJVEoFbk0Tp4KQA7wkXFkA53KRSWeaKlYWYyzrr27ZXNfv1cm
CivgNIOM0xNM3lis8VdvELEBkQS6fA+xUs5DJ3sMjzn7R/gaI7JaehIAO8fnEH8SRJ8fAUQcQQZ5
93j81FRFOfH/jEKs9eLQ34fhfpY2dw1NE77cf3eFsAY8i0gyYW0+M4n7b/OTvhN3ES/2VKlqezTg
jNALswjdmJ/vdymvh21M9DiXcpkIDTQDF0FqVDfegEUheTZPdqZHPSuJQA+psGgKsXt61qs/JsIj
C+qUQk1hkLjdi+mPZ3DvSJkW56wUfF9I1K4DLftYCzB6tkeNwcrZZu14/HNNMzLXnGrvTgR9qYKb
itgkeFrJLBwD6nZdLHUuM6vL+RlelerJhfDDJdFYLIasHnvLgNvHjsanBZUt8OWWQE2JeAThKTmG
KFqXqpcPMuI8gmvdYJPkdHQDR5oqwyrYG6Iuyf28XALb11W8IueEvV4gQb96ofcgEO7e0lYFww+G
Ma2h7x1VD1TJSrcZDQ8pL3Nd90d1gepf6ZAdpGt2sA9xHxCzFr2kGwkWKXHR7J2lNCftBpZYp13T
3pd7+s9Xf1R6K3HeZz6Crf3zuPx+yNr16FN5AQb4LYbRMjtsYa636a1Q1IyfPNOKJTPkgtvLuk4E
EhXngOpVRXycAz+FP2RFdK7rPhJDECZsesSB6gL9Oj4lwIGhWxPGyK7qbdTvZIgqB7S1oLY6XBwE
+YkUGj2DvtCHdeKI1N6/BijnzZrryxPbjKxFNB10KA2+vF8QttUJYkvQfZFEx09+j0CHwEkjkEuv
KhfCgf08g8gpzjXadXHElU84RD/QbV1zdDVTFjD/s7VHre154OmPkfQHstUiinXPUGfzRCtp3LTk
H/D9MePmjG7S/sPachTGtu4cUsy+awW++paNFgsuJtsgpLOTHceI1SxF2ZFfOj0Wty2L548iiX7D
2zpJmzBcKOc0eoKtYdc/8UwGbINCE7qxAX222UamL+cCOwlSJZwpgF+n3lB5ss82i1s4bcaiplmz
tulQF0/MZ20/thKBmCODim92D9t+nebxXnNw2ZtQa8nv4WQuZO/uiv3aCKEoOdBQajwCRGLTZ65e
IOdKK8PvzQ6gwPpSTHQCIGrrilHxsVNiNbRDgaEeij21soBKOhdtLGXBmpbciWuYxCz2BMoJggbY
2EPxNSa7Q9k029xzqIjjjzakYhKbQjZrhtg79kTybdFnescLKQ5QCz84lvZ0G4EgMflbfrOR5VE0
NrEWGOrEvp9jMuxxT5FClc+40Cx+egyWryMAufiXnX8z9rhtAn1lw1eHqFSs6K/jHCuVuFfVgdi8
4hrDHScwd0OjwKeAkeDRnP/XDcMDntB5ZsdY4+XT9EW7extzwMQTA//+fjwc2wtdYOfl/CbUdcAj
LsEQFXdn7OJfkfON4RhOHbBTVt2UGE4H+22J8dFCe12xBgdzgjiUf1Svs1yrmIn3Xgq2gENcKiAt
0nkgcdEedts9YP3/uo6J/pIQjjzMFvELUmTmTi4EAX5pGW2g/NSRONzKWV/kJoaX6MlZMfliXvNx
/6kKeye2eaV3X/4kud0awJAAFeZ6kPqaXMeaXFcOs6pJUvFQvu+dglcRoPe+Jtn6V8tm3Nqd5NeS
9IcUBK5fkEiv/vyghw07VF9d/zqyc+6XAaN+hawp+dl0AeX8BpQmdUxLJgAGK2h0jo5YIWSszEjv
BbF92/2B9kZzZQ/T1bwRj8fFyOa1hfKb3JUiZJorRtLBsw+JtDzhTJnEDKxc8RJDyfbreWwNy/eG
k7CFj553TQdq68J+b163yy2Qbcq87BtiV6R8TXHJFncXTuyGAVGnUzef217kzjPNwQnF0aIrQPSZ
WEUVG/gjKRBEQaBDpJI/TUBiNsZVJwEYF0ZwWj1NITzg/OlDVVvmeiOYPRrL6uTnqXBA+qriG3lH
oCKgLo93Pw80et7nk512hKS23Nr5hSTNgC5zwrU+dkXyuah0BKFmoSTCIf7QnswT6uNp6Q93snwd
dEGP7kcX8V9dcLgjWntRzGBGe1caMHkh12/Q394Huhjv/oHP4NN/OY4vYFaUEpDHt1T0O8BEGAy9
W2TiFUsqp0m0l1zv0S3ZXFry6Bfwjv7pAUE5adDhH9ViAcT6KzVpPYDM1ITocX7scAlpBF57qogG
TpjTXsSi2o4OEz5uZle69R/F3zRlJlA3HKE+BvMjiVME/sgM3ldUiGqzWetZ7dt1ko9mRbSqR6Hx
qVFSlWJipMWCdjCDbqzvp+gQfBBijD/Z7LH71BfP6EiMzhu2KUkuSTclGCfd2Z3he0ECWvzJYxDT
jBecLLhHiKqMxguL85LNlxIlKmQiDyiNsKEWgXtFzkRHBF/V7HZi3sYUD5yAIauHOwpaI6/DY3Zf
rq1DqWvuKVHQifAogCIBT7ruz6M7n+Fa9l369lCKjkSPbVDIE3+OBilGGyYZOELqBVNMkpPDSWgp
T4GPDrEo6Bwm2ERrvgHdTusx8dBEzuVaNuPgMDmIa5L59GfrS/j0JvzYUjG9wkKu3HnLsl643gN8
qAw+1QdL8vP0Aet8k5d+6FtNRAuKMhf8cviLCrAUEL5Mfnfn11scZJWZFrsB76FtLsXH0eWUBz5D
YsGkKg7k1aDuJJ455GRqdxdL+aZHKfNy90sfJypHUdynP3Nym/WGmXxQA5m91UwzT9+qQOuGlh2d
dy5Tn4h02WH327Q49E5nmZs8foN4zThZd/F4IlegftpgIEaWHTe18c1qw5hdhv0IstYImDZoIPHm
VMDnhdX0p0F1pZKgXDofqQxR/ZgkAgWp6KKFNtAdI200p0ES0M2VIPuiwDkMv2BlaIe7EQDvq/oa
DlGCwz/7TUwfKfvo6NdDHuav153GPJICK057ClCr6YEv2C/s95ce5F0FWpi4DdLHzmBjCdbf1BQr
lS83+CLOWPKp8qSLUH1+o2UlkRUcDmo8F/MOHZYmWJiJVZYaJSLhoQScxciq6OY58iZcjldnrqLW
8QbFki8bjRjIOqv8HmTHSaX5tktlkmkWbgisU8s/8rukrTXT6Ut7kc1/S7qvzwYzxx2Nk1CtUpaN
ZEah01zRtqUqDtm1x17sYsQ5x4SXJbfNeWVglKwNaLAQd0XjZFj4bolPLLNuZVJgD8bD0dWVuBSx
kjghTe5pqlyhw735bH1rxJzdNIA7955DRQpXtGLnkSz4I3mnBjuQzwYdIiRTn790m+f47QpdxOKC
uQeuS0IkNn0qpQzm9aKM/mfN/N68PI3daStMbTdJmUCMO8Tc9TDUlW6j4UXLvrSn4Zg11yNSjcUO
m/mr+Vv2zmuFvpgsCodpv1q5BnkOiPUqwjM2RtuN8BkeTXhK8Ge7Ue2SAupk4xe7uah3sn+zaJzf
boxMfzq9JlmWjm4RwDYl9yfrhnoEz158+9Xwt7N+9HrBu0/HiQqn7EuyRjAnwu+rPyshcNrDS7Bq
S4ZIf5e9gXwSwgBmhSjsPwEWCQu5CZVMIgf8kYco2BPlRTZhh2KkaSNqeEGG7ZozFfJ8fJaif9q6
9tUlfbqkzreNtN1I9nfHEIguHcwkdAhonRLhDtt/djWNYTKvGxIvhxEhLv83sGcFewZsVyblHywM
rqhOGIXh3A8m7iUzC/9IYos4KtL2a+UMq5YqXucjTMTkFX3FRHQFKBVPTYnnHC5lnCeORXNST/fn
2BejtE59pTtFjEyiUFHiEVzqwNIHx5Tu2Y3YHQylsWYopt8KjFHK0qJDu6NjNyCrF9O2Y4k/il1W
xybbtovbxLIOqr6rcW56/ns5HzO/xg/lQNykJJSZoWa1+xoxCI+NOvrthoGNFItp30BmdkDKp82M
ZqP200pHGnhuI6XPfG0voC82ESXfpJHeUNkXe/h1ZxKGwHQ9yfQxV5PgaWpLagUQYKam9xkQ9/r3
4EGbT5VT+I2uGYDi9ZfVbPWdfFLYRKNnfuof0qVLOm/aI5CbFh0VR9NgZVxspjfavPDG2Q1w2YNw
33wqb439n5ExQU+89ry0AmSAh7EC/FJG+sbzngvT08ZuKTKbv2qjYyKsGpCPv08Cn0LSmBZB8EeB
SUU6Lc8caIylh76mbhbSPi8aZ9WHNxc6o2hkTIz3PkGE30qPLmTfjJGq2alMF3dL9IhHaM1xxMrY
GHUxF+fhSMgUGpAGhl+ukIoboU5gY6VYla2+6X/N6zvxYV6WhUSHe+oLwzY5e/nfNFOnHweq1Ty5
K/akzn+BvZ0gpG4FhZvQJt2yR8peVkj+gjWlJItCrOkKJgsJZhuYDY+wvUX00WO8fmezKn7BR83J
p/BUaRWSl2RapWLBdC+Jc8K1etDaky1zgaN43DxQea6lBQqKifEHHMWOaNJl76fcjgg4By45RyJW
xbcfvp3W/6g28DOs53YXsJ2XlQIqshX4MeNFznift+Hg3zw2TM+J9n0QMiPDFcsOJAyYV5R+Xwxy
COGMk/yOFoDB8CSZWRSkTXcemks1Oyx1gIRkK9IrfjsQP6xAaWWsFzqdIXyCE6I/a3OkyyCNqpG7
YbiT+ml8ZGwwwoNtrg8qIGkHsrfL2m27eNNG0KI0U29NfeWF7eyTxkY3ktp4VUOhFoCNoWuYZlR6
s87q52zw0n/WiBZ8V+OKCSGc9zLIUD07zESuwYNeUFq0zatH9LS7bMlUyR5hy2z8AMMuXX6Eafww
UcOa8M1+8ILGnEakS2rK3icjSuum5BCSmL7wa1NSQVjGBKrkIXagUxQws1Pnz4Vm/gX6wXLhm0wj
78y+N67wBjHAaqDmjDcU6fzQIHQxHMM+dnwJ7Oe7fVpEvZBZ6bzNX9XbVCckNseZT/9vNQW6bB16
Cr6KM6hBATsd8KxFt8wlqlndx33/Xkz1btB/Wc/RB3869Ut0x9AIQXbVHsHrnaMu7c2f+lQq3XPF
gQtSTh/iyNuwSZxeXl0rtfLU2YGFk1OCiZ46UWie+eaPBmAIhBS8NiUOc1E3pRzjeUk+/8EDygpZ
pwLcnVHZR0Q+Fv5Fb/UI74Cj52nm2mAiqZiYAIE/gxJYL/yD1yEPZd6amKNPVMSU6WWfeDpY/s8e
MbcKtNw+PlOOh4zA614+kCDXFqKS++yc/xOpoIJ1QFUKy+vGQaR1L8aBChbv2KwdJU8/JBxvwJEa
MlXRxQ3yHnW8BvzponY6kAOqCEQ1U6/ZVQSslWY6rcIUaBOFCOCR97WqVU9u8t/W3LtnXqN4QyO4
/56maxNxrJKGQ1b1HNZ9Ev+UhrI7mPrSWVcfHu135Fp2e2ypGHL9/5KjgOg99OotdGyaMyVqsMoX
YR9PSuMzW05pqvK9LHq2O7rDT7DHrG9CODhYuOrY61VgJyVE+sVLZ46czJk7AlfziQwIpCaNj9dC
5sOcKSpHfNCU7E7CCpfR5241kb90Q+6gNWPE5CEd8Z7NTv3rnXl7ODLevmbTMtBHNenLMY615muk
GjfwAl0FP8IMkgu8hxVcCS2Nlq2ebYtNt+uhbRlBdr6OsRgxwNZkA4odhXCHKccD0IPsSM0lUs7z
4btEHMXkw69FBiQiaNgF6QGZbcdKrNDLFnHUpTS6FZMa70ythJIiKBCLCDWmSRuwCsyMAqpSM0wQ
qNZAgydUkUAHGw8yhobk1uxD7j7EeERzbUOuQZVTfa16Uc21SLyUlQF/MmiYfZBxUamVWMpR1XOa
p6rm+Sqc6WSJz+t0xGlAzcporXL84wgo07CAtakoDT5DlfgwO3F2sWLlCtedtMc+ABRou14RkFQm
7QyYzHlYX7fxQdP5G+jDpkTExUElEd246Sp5gxD4yOMfVUM3keTRqcJhDF0Y4iejfDiqo9a9xPvx
dmZIF4uehrHnFkD+IQzmDj1v5mXGYi1YDdziCsJ5dphtAW93Pp8r0jOpxvxIjtuPhiweG513q49S
phbWyXH5oAY9Ns4cewNEHwLVxKyvpZ0LZxnMt32NjIXG+nZwkIxSQqHQS7ZZsT2WUpnNUnBhQGmW
2x8PJMUM0aealeWzQ8I/PXzQuKWpzIElkHTraj1D5G/whpXTTjBq4pS1U+xY4ZReCU4KLwGA7BdB
wDXG1/7xdXjL1fnL0fYehnZqzAZX7iwbLo9K+TMEeSWWw1IwL+ijs2yLytmwgVQEYZYtj3Q15anS
aTGcjYQuSvOP8Nt5A2hKTrG8ylP0T6ChxTJmckG8oWhDalN8vBW23GDVYMuica/0gsC26bnXpTxY
4HoazuaB+4rN6k+vVFQ23gB90TlNFNeyaWpqd9Wa2ew9HxFLvBhDxYrxRWR/QDIKM3VQLfw6wca/
0bVn6R5RbIYYfK/umezLpT8kGOQEHXGmKhFcauMu/ty49vQd46YoBmFPuuPl6SNW1x7i+0N6J6sk
yOO4dZZU7Nkf4V/Lf2ikTSldE0UngYKo2g+ifyG5T9C1SWlWqR+yI4PSd+OUDdmVNmK/TeVsYDTK
fAfS0wdf8Zl4IT3waBfDhCCNRn8OofkkoYjztI0haLqJd8dgr91X/vjoH+aAlmInROA/dEfLoC8c
Rdc67e8iBCwZxN0CJKsJFRu3NroZkRsbbF6j/JDWodYalOkv7/0Nc5FaUrMUhhDQieonFA8MOk40
A7LapLorDG2m0U/KsAp7+TWbhj7EgCqSVD99mq/R4mR8PQqtd/dSe7lih+Z2N25/Pshpqp5Jvj+1
g6GrJ3yvksfHVdQIDc3P6ORMl9FD9Mb81DSqDnQhoU48f5R85wPA/QdQvj0YvB0LExWtjd9Awm6j
QjQTJsP5l3uZ6B0gtcg/k2TkHqv94/Jl97Kc91zcRVdV5lkyke+FExsCbxpMSZ84cKZzuaRI00aj
USzbjm3bIxDqMnjoM+qKSyeBI9snRK7DG4O4MdLcRpISKPV8wp5aQBbdUiN/ZUSYxPCOlUTcrmwK
3yqy05Kigog6aC9Df+hrdGLOKDHEefG0iSEXnfEp4OwMHBIG5WBK1DoaJbUQvmF2K6PIEqJ5L/Wx
azuoRkOWhcxZyLmMmFZJlVxVh4B47ZHEA+ch9sCLHBwiCfTbItHAIu2R3s7ijnWNm5G2qU+kqgCZ
62T55ZuexjPBWZqbOBBlao/6J7yB5/8actqJx/ZSEQI1KIt/3QKDPMIkfhogMOX7FMjmWc2tC7aA
sGi55+3hogTdGA9xZ3fzazTfaetuMLsJgxiA8de/3eKCAZ7XRlyISyKzYMOnoCCUC8mNOj3TVdWz
iOAqew+ZZZV4k2Kcj8XilCfbLCVhImDC/TbOo7UVTn3Z+QXCTbLh2mKkh2iZowfsuwqhUEsQwmvN
QA+hiJtzK0yT0HUe7EEAgLyPd4rDCXVn/oQr8PriKrKdNY42iWv61R9Cbe5KiGQEeblM3/YAekBe
GybGLxFtWR2oLS8QQjDPCsbjFElDb+bHEZF4ykqITQrtwWsoaxScLG2YCTfpWFsSeY0vRpEW8MtN
b3Ou1ImoSnjXpX8I15oPwC9CfrfRQj6EmIZ5R23LSx10Q2E9gosuGgI7xuR0xYNG94vqDmktiVN7
YRMG3G44vRgg1PC9kgd1LjVK7ahlnb5lE92Nu3EvfaVehgICXdpE5lIlCTsVbcZ1Vywo9twLMwoQ
Hi7Qa8w7jPxHsqS7ZwOjx8NhBcrJbCkR3zQbslY+HhBgQlM2WlQmBQzVC3B7Vn/MWH+idEEyjK+6
j9phTJWrHNEYEVHqh6mgOWA8K+cOJo8UWX5dM+wztfVVayqgiR9LVubuEvC2L7pl7aXGuUTmiA5n
sJOUNf/IGRVPWdsmGbIU8yeWmy+BzS38TJc73oef1ZpERGCilmm0Ql/gTitbjMJQmDgbo/MGyqqx
2sXxGrrDAdEYBZq21n0LCRjE7btCEGq/3YqFTy34gQJ4CCzgZsQ1jZ80UzCz12qswGyAB01iPScB
cD954WcqlIN36A3KnKavIfIaSRECeMCctaD0vyHl+vBy0APXwvFX/Z11kiCw5/VM9T2jytz98xiK
ioWGOZInIpWbk+KFjCkHytw0MHatn+F4YNlzUEEhgpUaMGNykbvIJfTbJan8RQnEvqWeBPyI0XIW
53o+eB9rffacZpOQv8TOzLev5UiXVXJFwRSMENxsWfcF6quQR2uHlHRH7rkIFqDuu7GcyECSwwtm
DKNbI0OCeVZfCErd66uPna2jLoOMDokxRlYgBpKg3VvBt+kg7dfNyLFloUCsIGpkRr1lT05b28pL
fYxi+3IPTQUnIM5X+jvgwZIW4oJcTCMMxBP9LZB9Xwl8V0bFTU8ZbzQd5Z414jhaMX0fi9KWeV2C
p5Fv5z21uDuht9iwPXxGK8aOF+9dPyQ43XO7nBHb/BZ9Lf+czDC5e8EDtn781RUp5ExS9k/luznk
cUN9mHTAMXtD/ihDMtuXMYM68TBdIm2AFu13X/CvKIUKDv0lrHH1nMkKAi0Q9UTo8jpjQ2FT1y6P
K+Ajn4oOx4FaK1B1d7kaGooHyZipNOuOo/zG/qLlao/Vu25trlRy4KU/KluJG71uZyyaUdIHkQrO
BxLV5HLsQ1r+rcbLFNAG1MO7d1TxFmEYiWAvZssjpxFKJ+M12lBJgyZoqDUg4Lo0jjnFKsFBKSm0
1CZCvEZ/OOvs1/sjyTW2e8B7ZW5dismfyAWpWxtBQcCUnAxHukOQK3W4ALWxp8o48D/4qZ1/ttjA
gW+D+ZxdTLBccrR1Pvyo9DhT59/d6M12l+6G2ZJkBQg56PYex1NS7PJ/0xCxYSvmd859qnRwsnNh
uoPMRVdmcAgUTeYlMGjKf8lpRw5ebic9aUMbxwXQd9sBq5/m6q9Q8Q7YWArSHJ+Jnke+UzncX5An
+JiY4ySmOI2Q+GhDDKcWSscdDae7j73+aKvEbh2iuNB2+VcAQcVysM9mxcaDxmasJqAM1m6h6Gc9
H0zlU6FO3dwSzJVz1WervWbBNxkWvVH9/0PlHUbpgQNOka+W1364dz36kk771JroStQXPcGNWVSQ
xqg4G158N22+mltuKN+p+Ns/KK1CQssq0MxCFgEFOEB+rZiXDsnzg9NAcrkaw1hci3JopeXgi2bB
DWYOK5WUirpfXtIrGs5UoFeaSVwsPndE3FWX1I4fG6JaDrCONRZg5cNr2LL9rQYwfb+fVmPWP9ZY
4HlS9P+it79hh9B0qiOZxlslG/WlCWPsR2kgAHNw6jYIc1FmKCYIfZ1IwSqSOAax48twgFdd7gJI
8e1CbtHoGbwa8CS72oqkcLpCDCqHlMofUuIhaDprBUDUUFQN/7i+K9R63SHCekzGTCkA8lflKjS2
uhbyr2zCb5Zli8greMRkIC4qb8Q7mmGbvtZi2mck9c9sDfqEcHphXlGz4UhhYswpRupwoMx24p34
vIg0ALpcnUsJ4DZaIvHI3/dgYNBLnx2dKXVznDjnay5wBVwO3aPBknpzR7ILLyVFhpEWWkQCZyr2
Hq3u+33NeZNnyuPEn43jqEWM1WfBXjEBI3UoldzM3vxQz9PMqWMKWgFcThieIr870L64g39DB9FX
DUJPHb++pu4xz4/a6dWCqtM1pWllUeP+DoUTZeDBJT2oDISyCX1f2w2OSDWiTMBJrYFeUkH2oAxB
WsG3aISiN3ck3uxJAbv+T9h6p1wO+bWLNkWL+od/zQLUsZTMxdio3OOxkL7m/cViW9wvoVHRtJQs
5+SL79P9JcQgVXOIiMSWRM46CMPibKl9gGdNNmzI3vi8XqOzsFhYvv5Ufb89DLll5Ux6MePErl2O
WKZjQUzKWXRONtlxigvkv2fECSvTJaqdOTBEgQip1wVvg1oXn7axhYIQZFPju9QJAaT4MdjPBJgu
30ld7/9LlE/W+DbznaqK3s6sXnBkWublqB8zKitZQLaKGsxKc9cjLeHWARm9IelgP5xvOPzS79Ah
mVP1tjw5wq7fbqbmlqQpQ1IHDZ3YYfgNqLK17RXgzQMa6M6hf11ambt3mDoPG/WwtqtJzmu+Eqlb
nQmrO4PRikBX8rFynqvRfgdOGoELttiuQHKKqVzAB4pb5bHsi6l2ZpULPDI2l1dxq59Zdlky0fhY
XEJ8BKOjzxywU73AMkT/Q0Ryh7ZR7m3S0TzZEtdpR+D0f/nruAcLMQf/87vIEkPLrAs13mKgnx8Q
riEFR1obb4flWYnRTc0NSww+u0i0EiBAiS0T/uJAxh8y1s6gvML2lGcv0yu8sTrPqS6xlncQ9B04
13rozxM5ydtzH/HZdxOMEy3Z1w9NhkM5s9HQWdZtR9v4PqNrKG94Aa/ecFIP4O9w5pVhpTjCLueZ
tX+dkj1U3gp+YBJ/kg3qsIV6TJ4pg8LLzbwdb3zeGGH7GqcoB9Fa3eXDkwsccxYQ6MknBdIUwpJN
crwPgl1ndfd2Xbx1alH5azJWaD77RPNTwsWo3zbUbhQtO8vhddSZhILoqDdskIm7RYrRI77VSOfY
aSj1oBPXp3Oe+IUIolGuM982YL8hsF5qgC2hu3sm4QvpnX7yVdxevgaXbqf/mHrBFIkOmPfJC2nq
+fMkePKJGJ/Rz9L7aqlKPGFvL8rxP9zt43YvW+JL7vR219QBfq81qzq0GlvQ/Vc7OWJAo8jpUkCF
Bh2MB9u0AkYnHg0jGuHYh/iePUrykLgNZmftZRVF4nkxolAqgZ4hhbAaWFsvP/6vFTgwe+TO3f4q
udBGeP2NwOiGxr5O1paoR8pLy5fjQ9bm/YkUBsqguDmwDMk1a/YX7ZjdhPt5JWKYEICOhYmp6FAl
o7XVkSUAHYftfHbyKmgtU2b5FNk0FPxAq7uua869BZFEgoBwxmiis2IcARRn19A2KF3+BIPum/Gh
KzDVfVl0z4OdcC1IkQaN5LVg5Q606TXZp+VYdjuHo/87YbZ2s1YwXVunca6aSaAuUVCjpTuK0QxX
xAWDSfakJAEQCHB5dtrHsjhINJQBkGA+TOEnUyAejz8ZGT3c5klOZwA/zqP3eMWDfR9XL7ftt0uo
T1lZIg3Uxanys2yUvSbHb6cBZtaFOOCD97eGgqJ1c/N7R+uzatP5izED/xl/JfhGwIn9cgmkrlKM
2S7dW75uYM19SO0mOukKMdWS0+BKidxi78/GU+Dz76ZHrTo5RdR+zmzHp0w5vQEN7OPyutbOPgOa
g4lflruSX3WJTBFzqe+zrtjxq//uiqB9XodxFKOaK869/zwv+IWuMc/G2lQrADuxDIgsCZFN3YHX
cFCZZ6WNve2XQI/9w0PcNrMXoL1PF3WkkbRZk0BIXBe99TThQ17OQKewxn0YC/pimhIRlrSMd764
zm+l1tCXwUWKHtfrQ1hWGCfkdQmhgY+OiTJ4IWig28D4nDdxPz3/anCH4c3yITwIjQ8tj7a3YBdO
TDAtPuCUmd7/zLq337WPIFPwBSgMxoF48Wh4o9MDhCS8bKgg1mxLqhCYQfoXoLXrwk9MNwKYUpva
/SjlEfnMzuqI9YhBoaneaNNER1bQiEreC3BN3I49kOsbVUjbB4nJhjytgFbnAXKZlCav7gug3KEC
pHW5g6kOBdbFaDF6+kVuxBkJE8gyTXryVXYRuq2Q3azJLO6kEnq13i3ZcFGJqgE5Ke4Tyq9TKkZc
dlRjKS6ReRzPJi/cHPb62AligXWiJ6YZr0a3WfJW99b6OVyldZk0x/ZcSjNxmNp4Z4+3i0LEp7vL
oHM84V6PRDmNVW12GF5hScpbjIw2w7lmjVECBpvSNs+s0aztWIpws5egOWPVf+f9UsJ9mMz9+7FS
//3ZUz+Ue+2G+XJ/fiHIMySIoaBOn/exJpMaPAlNlRq/j+PTguGZyM3DptjWop/0dWWkcBCBAJQN
oD+uTsb0HjQevTyqhCYcXsNmNeIOW9QY3Dh501wmLEyRXP9VE6OOiSqYF/qhpUeQ9mHuSvlInTOP
6Gk31M6pFSaLe8kyU9/gulC045zY2X0ZwznFkb9+6fhGp9XGiztQMMQJMMZmKUIqrYFBTepm8Eco
Ue58uqeX0cHlNSZ/Sf0aqo+M2QhI+BZt6sj2w68EuOXvACChqpXYgU3eO63pswoJzhJWya6kaw/H
uEOuoemB6d6SvV1Vx/tLORUKSOjV1AcF1OZyelEtrMTEpRsJyFG9tNIKkrA7NYhsS/up5akiAFhd
/2Kyx1B9SL71Nk5orLVHV+vXs52D7zOpsNsWUL/oFpXJAEgq/RXT5jMnDnPJLXoR0o+qT4+NEGl8
v8Jg0mtQpYylJjowfX2gUQSkKHwnwxcIFuo2IU57I4E0jOlkIc2J31uUrQK8lYje1CsoyJsecw9P
BbnvkAoCYQWt3796sGvbLOFPajyaCOqcJocvA76+c6pX7wJ1WMsqrrUJ8/eiMzNONeuBUzV6Ooem
tacJ3G1WZyh1iL3zE9i8skdcrR/7fP1yKZGcq+/FTIEycyfG1T88yP/VY+60+81ygblIOIQt3A41
nVXtR4QBYL5f3JAKIOTvAyAGc99ncdsqW9RBLToOkaBjl8avSPcZpSPOmwLqoVCaAgZYkKCWv6WU
dOkpWl/ggCQC7Rx5YqxeQgX3Jc8gRAa1v52mlQ0DpvwJqcG7Yw40DlzdGqRZSOqQjI5IKj24fIxB
mft1VKzq6kzKQoRUXpxB8V1JjsprcBSLGhyFCgaItOAaV8GH2CARkxux1XF0rfmBERQRjjSxEWwe
sLdEl+GLCe9R4HcimxhJcDJD4Us7d/4FTfYyv4IGlLx0JMdjqaZihTpOIv+ZfK1Pm4npDPgbF3eA
QxkEHV+iBPC30J7GZCXzzz+dBiEEbErh9Z0BXPHnT19Ii80h9p9sxAfi552W0xsvqRVaa8CZRSrx
dEGWY5/y1lbCh3PyTwiGgU6+GNm0lf+xIxb+TkXR/i/NnSBeqWYy6dvJTx6Nnz7KWfiwzeUkxoYW
oPHKKH96sU7pmg4I++7NRWZ1dWoOIahPXQn5KyuMDoHWIOxgTDhnIjUEAHa3GxL69AztWA+yzUCx
T2hKpNajuFmcLNoxI9u/tcqaF+1NNqYnr6xsh9ev8jQWVrZGQBOc25uJozni3sBp5z37Zu9FSXvi
QKAueX6/Vu9wir/+pc4Ir3uWXqNoF5fa5Kcq3nBke0xoYND/EQujnfhG22QhQFp1aBdTpXESQ16D
wuaf+V05uP2hlw0Mf0otoMe16DvArLzfs8progZ0o+quTRYght/K1RwlRINo1s5ucUFOv2gY4IbA
Pskc4+ngysCZ/dzdZRnRS4avlDwDfx1d/ropMGwXEqzxDrSuxVnwG3YOXO8JAKkDf4e37AJnVP+P
avUMEU6Szsq1bqNrhdzmRjNtjsCoZi5G6GoI1OWWHhDb3oexXQYH6e1Tld4xuEKsiis1nC/FxiYt
UxgaExRIfbxs7qAJHZ/FJO/0OkMzYdD5Y4KUTlAuuLbMoZ3x42l27YuBrR3WEZxZPqlBk6uqavXj
iVjurBsZnvbeg4gJ0cGKHkbl/GezV/XJgh6rrlBU8xEfjnPNkxMsYvJ7lZSLnEwIHlkoKloeqHaR
6z+0oMJSoDPqLNZjQ/xxhPouQ/V5B0K8NG3UVhdMhhV6Ayy3GRGY4xXx1c9aDYBysCcZEJcAfM6w
avUSZozGA/jnRf4yPWcgqgQgPt5EVzotBXzZDX4O0QFqZ0YewBA+9gy6NI66VdimcoD9OPlbUhBv
GRSi0ElgdfBileoQaW1PEu/DSDFWcPkKtY9dNWS6fCZzyZ1bbT4F3nKOelWALRLPJ/6TxX3qlU6V
9r8BP7BIh+aY73P89wTz0pyJY8YWNCfqWY6esSTbhlRBr0P6Ihrw1m9s+8+l1Va8HOA5Aq901ZUL
AfLBlRFdasxXMMghk4aepx6I9gtrdj3+zat9OOre6uIGOiLm76Z2rMDNoiXExyGjRg7Q0EnTVsyQ
r6mYBS5xPFvJEyov6PJH612j60NmgQ3r8KZxnMssdndAPrx/WBtkQT1zkBxh0R2ntSAHNQM3fwYD
TxymFQbGdUMIvObtYottlGfIIMDgd8es+MIWOIRyHzQnuKngTNHiWvDmxBw5iE54E7DoDzTmhLA4
qN69yxJsfoFs3WEFKzqpmIFNEFWHh/JDLqdY1+FPk/tNWjXBhJEQg4pGMBufzGeTuqR6PRM5Pdoo
TKu01V3x+1Y2HqtLjQzAqVrUHYAIzBHX6U3c/2/0BuwpZfi/dL1T9fXVqKoIFRp6Jj2kd3L2emDY
9LLDKtjbe+u1C8OLPuCprEiEYLyzGCRCH8KPVMpI/2+lqit4EUwf07jCX2xOIkGskSovTXRoVMx1
LwyxsiZz4NW6XGz0sNgOsTG4iEl890eOFYPK+OguR3DSTO04nSoC1M2xOEMVHmRu+XwK/cVi0lfU
kMMISitETar/Ei1NiGRZC5W4zDVWQU66reewTkHUBoKjT64AGj63kNdTotHT05ccZLhnA+4O07WA
JJyUHjaOinBGtRzeHnGkKAxJYIBM51hNuDDTU6qRsB70pv9LuzbwvvHXG0MIxzhOAIVa+tLkIwwc
cde2PVyybRVpBx+jYD3TJ/vhQf3nBbCXZPopqC7ONeZCzjS5rOMFiKa3UsfNcq262yjXw21LK0BO
gFrYLNw0bENGTDFcpKt+uEM4fkP4Os1aYhNbmPtfhjPwEdwY1O9V3e68hvgUBrFGWi2gTSvMwDYV
NoiUrVmIdAfv0c+nSAOrd0I9JMRTlXzGjCOnSIfYM4S2uytY+1FgG5trlWl1/AYLRTQQ61yIRBfy
xNHmHjDwffuAUhglMekty3cd2gtaVNQnxZqXmXrmDPz8ZdTqVzUirwx6r29e89rj4D/j3JE3LZ25
HHn7fhTKTL66I7gQoDE+iPT1rY3+DS7/l9CLDBX8wrl3dcK63ILNDJKdv6IsVliAClo40M5UKkPU
uivEtA1aE2OxP/GsVaFSSURJBOhch6gZXYqF2LnVrW4o8FWe86yreYSAMlroUa29SErd60Fa7Q74
Shf6TXQ0EXo3cZMZWgRpOq/R05J/zPCTuj4JNpe3f3Ec3umRLsod/d0N7O77qwibNy/RyJJD21lp
WPd6S2wBLzyQh5ioM/y12fyCKQ7pSPen+DcnOKHh4b/UU8eh40WpcMjRulYzjQmizTxgs86NMSoq
WkKeCx7XsnXrqtRHcVzlOTzJWYO3HwHFq7KuSDVLqUHi8saaUoWD+8M/r2Q1PPKtzHZwVhiLPgju
1qBgpAkzelMi4i2bjACotMWcu4WaRi2vh/RPTZf0uw43zGrkNhhCCVDDJQ0A0AB4RUOn7r9ppSod
jz7ZzCdXMSelhC5ym9SqOOidM4c4lfcD9oIJ4YWQafg3uzKRydiNWvOwaFTTn6bLxv6Mq6uxHRho
A/34sjKv7JCrL35Z+Q8JixscJ+DF0rDp/mUlkWy3LsvCElHmKsYwHTGHuRNnbYrnFuJPtcAk2BZx
XFywrzfjg3+xj5osraA/xZJbVRBa1bwTXLLUeeJWrX6UjloEO/8MjWp2pCGbFw5TUtnTJsCOmIoX
eRBXAyOVRg6poGt/mmWiTKZgb1F5SrQED1IzSk6R1fO9Wdoxm21CVry3MUYbLXON3C/3efjE4ANL
nc3U29uB13m167NEqsmVHGruSW5Snkv31yr9Fykw9roq4jjLlop4brZoXYLpKKu1mk4axj7gUdki
CG77UXbPgfpSgZMLERIhCmRGGFPmpQ6l60178gowyeKa9j9aU7L1e50GAruCI57ISCHBHbsoDmJD
dad9MYJKlieF3cX2+nx6ZzUsWPuTqc9MwhrN+RZYS8We8SSmlBveosnPn1+EaPVXgKGqUlevA2U4
bdWPgplL7Zr3+ZmPFHkd2FNwWh8/ALoprM5EzPqlczEd3Zqwl98iupiinOtkFpCcoFph9Z7frt03
yN4zXCifsG9OCQrWKSUvHmca7jGnieWspGyKxvhji+TYseTCwS4e0Yd2dduRdCoK8PnfoY8/IA1K
6za+BKHXTAfG7seI4PylybUluCNy3QvMQi92ixpx1hs/tKgkstM5V+GOcWzFrVcPQ3HCt3wPvw3L
rid3tCz6KzK2quJRtzos6LF4e89MXuftD2MA0WDjDzY6w2PikWXey7HLra0TEqNaSCXpthoHlxIz
g3TGAFwqFmm73C58gOh9ut7+WnTPS6ORxYQlHzsvOYHe6n6jYhpeLu8qS5gW5eysiYzZCifuqn1h
vEvt5m+OBEtcjZq4cJvmNffzF+17+Smw4HZc03zoIW4NAkQWjeFcdRTF2525dD72gLeSnTX3vOl3
2Fo/UZv9FGfCe+m/9jZv1w37++zrllK1WHEnwvDN4g9dXSR+BwYOOewInxjeCsYAFaNCOAUbIDVR
ucOkbO64Y/c6vStSoMFg+S5QCs+VndEn1n2Eg3nFQY2IMZjqJCjwadCpvr1/1THGytPVS6GbV2jJ
o8hd9mD0JQm4sFlKm7xdgd2HkE448F7HeOpQYuKQjl1ReK5GSqlg2Pelh3viQ/NWPY5x7VOxzHEV
BYn6hUYHxjpN+ysGmgVfvskygVjRhzyykIpsmeEjCdHsj5997p++P3k9Nw5akQ8YcccCNO8o0aEi
yKvN/PdEuwM+SpdnGrk9rzknc26rGc6dtBnE6aXjr2kaNzjfewWE6Rj0NpnxxDb00ndoxSfRUL1R
GeNGmQTs3l01cWZs05kz4WM6MhcaZRQ+8SxOdnMG/7DNRZtrd2Af/0SpwEUnkHh7lB5V6E+4xfl9
7UQ0dO7QdiNj06UAvvCyupUUKKRFvZgOFkNbAMQh79/Mu5Eoqr2HaerphqaHB4iy62tcCG57ptSk
d3JDpGwzfAFYJdRT7VM3dENErVi8VrRkg1F+MQHXAPLbnsAkCPIrjKPv5c73LwaXog/1/IfaxgHH
x78GJqItHnckCivQQlpt2dZyxBWgmTKJCKjTO4I+08SgPlIDu1IIYhHbhNUBwfqFPwjp3EuUI/Fn
FYMRxLhF+UiZ789RniYdEJLBxnB021o7gHKB0gQzC9ObUY9Y3F9D8jNIpU3xySscwGKZSDByusAK
vhSPxbYRBC/LvsZ8c5vGRvluOAPMtFNxdsLYgMoeVgiD+5x23ZKFJwqtQkRV19N5a78MM3oqU2uE
gVbH4jHQhlK/uC5wjkleu5vO836LbSWnSubxLt+itL+vesj/8r4+acXH94OHwryiT5K9PWKR78Lq
m6HPed06df28tgObpWjjg9DBt0CyqZX6KZK6qHONZzJjmkrv2xwwu0C4iJ56pZOWxASqZ2zSc7RC
JZjHcbFYFbn8C7k3x83V5r8TYg6UJKnJ+gdPB1JbP37CIlsIpwc//8EQgueQ80VvaTwASI0W7/Pg
Bw/1kLqKo0Nt0curyY5pgVmp+ht6H3VSlTzaODhzvRZrGh9y+DNlkdiHtxt+G+giz3awezDtOKy7
LZXmmJ0vMbk6odQx3LjrAL07O+i4PtrANBnz5SD+ajTgOFk6Q8y/0/4pMI0hnxt/dF+YWysXiM49
RSX/O8i5YWiIsl7ToNx/i2EraU9R1ciobEqjnroAcSS0q5zfd5zd0U7DFarjLkpsjUW/ZulIdWvr
M33u1/MuUZ9Rc+w34RMDSfgRoXz70AoSt+BY2BkBArbrhxcrIUR0VsIIrcDGNKkFxIvj4p3kNPNV
zrK7MN7fJP24rD/E9O0+1Tn9TWf4bd8mvI4EIbMpkCM7VDHjlrD8WkY23Jlegok50UGBN2JtKKSV
NLjp6qLRvVofiAhbFEGbuiKlJSFHK9+ehddOpGdEh/d09WS0WwvpDy9echI3POurgcLDPZ/BPmvH
J0TuCnhU3HufrsCb8A7fF47Dr7wD4Z5X3Lz/BVQwr6PuCo8ZDn1iV9K/DOoOium8JZClAd9KqC+6
ePMwt0fvaA6YQJQtU5nduRp2RoAhOCwi1pyo+aHGSPkeGslkgXQa10ArXVlodTwYdTMu6mnopneF
Y9e7UaKzEzdAE3g7Im5Yh/oTxWXpjr3JmDW+jY7NDqvQvL8BHlQH4rrhXWL8s6iIAlaQDANu9gCw
leyWdGVqNG31oVB3aliLSyJ8XRcdvv0wQdaL44/ukXZMKGRph1eG6aY/99rgh4dntftBVNs/7W71
lZFESOtmnF0WEd20nCMFHbO0oD0ABl56PwjvLx0Ph/Ol60WMB2QvN9giM6lVsShFukbR+PF0mK/0
FaMt1uYvdw7bPKsyFTdsk0p/XGPRenPlyoO8/W6VcYOchKbi9dvmxnmmamGApGRJyeUbS5ckeVtG
hyJQBNte1FATcpinesj7zwuTVbBZUHpPW0yVV1ymyAS+FZibElWFuTtIvVhkDTekb6veAizTim+O
YBlXkGK3trx3k29digN9VKZggMX0DcdD8f1Rjh4E7Cl9m1Q/zV+Ye+oLHLN3CvlwULc2oA+WzNg8
CzvMkRlrcEsm/YfjUUxo5IkeSYv83fJnPUnChyu98mhdT1lUmQ16L7cNpSWghf5VCdkW66dpjQ3R
xHe/9/ce95IPR/Q7fyUm5O/eEFTV7QoLcdvy/mvvgFylBUK6kQr5coc9qP51DIhWEnoD7OMnYeEU
qIQ7j89FGnVeL9xzJv8aOeBpA0vw32G2s54y1dPHxiHXRp92SwMpAciRzN/6Cb9tpp40DSy8mN8E
Y2jYxUZuS98rE9/8TZSOuOEQCMSg8hwXH2SYlPCwLimVCC5lUO/L9orfGwHBsoGHBSbwnM9yRoqs
yoVFjO5p7I9FLSJxC3HH9Hq/5evLsTzS6MSWamMNz/0lOBDTTY+GTarf+1Np88M/+pQoL57fTwjy
zaYGG+EOUGpBrfQI2iM3W+ne56PpSwDgsVx8a8ikrw0QMKz9Yo/CoXwBgk13fLRhHBM4zG1QfLDW
ePcIflPOPI15OzDriCMkV6CTTtUygPHRhfzJXby/9jvmT7JqwMdDCNZaf9Dpp5Ct+cqcykBYj9L4
S99Ju/kt2PZBHSEaSBeZDor6hh8sdtDYnXIAi6n45WhHUUkdWTrMl6UVqktsF+Gk+joFm0pwspHq
UJIs02cFF7V2jTHyQ4gpNYHaKLWqFdUUaxKsg2fAMX//+5Sh0ffcNHwwxOQB8wyVDjeO1VvYYqTB
fWyp1JwZWI6o5d8RVZnZ5uNDpLn2Qdc4N9bc0lcAvIeMGh/ye1YGE90KQseJTfTY4ZozBwsyR5PL
PS0TZsq5JuqAu1FjumoeCYATQfVWTbbcPjqTCeGnj+ihk8leYkEFnuZapUOP0SRKM7oruaFLIIp+
kw+XdDaG9OFN3fg3G0+COK7H/xtggfKcoIhNz7vb1v3XpFFjm/7IaEIUnXDiHNwDfHFCyKLn6G4O
kxupW7mDCg4q67JMXupydFtVylicgyylKts/Bh+xbPB5JDVhzKkgUcvR7VH7SzAXZQBdn5siDzcs
b76kngXyVsG1th1+XdKzvBxnV3P3ltRsKq6WSUkLTYXeUAGDnrPdC3opUin0aXFzV1K2+QSlkUVY
Tb8MC3sdrXiM2uyH6yOaxNLXipSU6nzQOmpXWH2bO0GeW1W0rkivOcbvLD6vjmIPNUsxiZg2RAYD
3ZLevw6ifQZQOQL2mdraeq/ytPjlXrWU1/qicJpUznN/IarRxzFl5F4vyfQco96+Si7BAgjz5h65
ulebIv4D5GiIDI7lwzwoT5Je8IAh3eJbbuJtpQKS3FtHpQm7blfd173bNCZQ/ZjcBo1aqbmahlSU
tW4cIeWmwSEfIyFjehRs/UkrsSNwGkwCh7BaQ/FkJUbWH5kfR83uB193kHSBA/YfFt4eDCUs9HVZ
1SUidMDhdYebmsoZYZDOhGazi2wt84w17Zil8xHuz/6FY1/T93C9rjkV7uWic4kBscFt8+fcdql2
AIvpRBsbFivmGIFwYBGljQVn/UFqfCQpejZRHwKix0QMIix1kyzJnAQouGYMuPmjeiSLG5xrZN3a
1h973wBUOCDs4eOSkiH+VFRm29JOI8aQDWG/nVr5HBdwaQi1YH0cn+a+SG7IjM6ect20iFWlwvuW
E93mLcJj2ziJwnQUleJz6XQRL5dQI8snJ3efsQqAwCXzPbOFz4uiIuCs1iw+0i63wC9ymRwKkOW+
DlOuVo1nKFhSN1G0d7YCOhHoLv6ZB+eY4Yn0+3hNOWxHsOA9e0O7zO6G5kuqiMPIOmIbwQk3DOBD
amtQRnHxfhVwaagnSEY6hTYoRtwsxYmqgk8dG3mAfwmELGc/xckmJ7ma2DhXj9j6XcJYX+5ZRwTb
urNLHSWQNo5aB2fo7+SQcnIVHaW+buAC418pRba74DvB8EsF/4WDLdI8yb/O+L5gMUqlaPcUQ1NP
WEyNd/RCGAxIB+7DCj7DHEio+1cFKeX/uhQWZcQPy4MsYWrVaUSfOt8UHWVzgZt+OSuyKGov+rBN
jcCDtVyjAP3xEhURxwmGdxfUBj1HpkHedoohcXZm7AUOyFXABsnIqg5aQK0euG7E3T4W59n0KEFS
CSNinaeiyWaZ2I6tjUGWQnHl5llp6YFVJPiupIDsoHsG1AYcLs8idTUdgF4ClMY2yC/K/JWv8RqG
Jk2yoOzRvtbAH/rK8QT2JrHowfLKCdJ3Hiap+VThC1HHtOR06M0eIzqVvxBewvfffsJJUvSqjYkD
8yjevPmDs8OiblWn5UUIWXSUUF9kUHlYwXy8wHPrP/tjXFNbyYj96p/K2i5KXTvQlaGb9NGMNFmJ
W0wKhJynSlNfKS2RBjdDTT+a2lh1l3FGOLX0hvmjN6L52KQCqzRDw0frj8/tSPwMXhgOym6bdHHl
/o4vRgs37+f8jJ2d1plblWJLJKk65nEJnkq1/hJpK/NUzwfHWLRweleusXBgN2Bl8Zws59BJ3d7n
XpQ+qJoNZ3tW5JcFK3rJTMM63lyMIcmlqSRWjqw8+S9dAfWSkGPLcqBiXBNfD/eVygBSCEDpg8dF
uLEiRmMuzHs6LL5K9Xe4Hl+E/1WFp5ifBbfhuwxIL7z2PQklWtJR1+FDiOShZO2Da/WWI/fQWnSN
IHeB/JGWbYYU8Byw1vlXQngKY3CNahTv3JIZKdGBZH9ERqsXhP8mkv93SYQQFd6sOtKCGh0/6UFb
T/aW1z1S5NUSQShHVS/cUjasUFzz6CtlxIICJVqu9vSXB6qZ2wHY4d/aDD/+Itw2ZJC+VVd0Xacb
nclfCnnRAO1ExTnsCgnp88T2cI1dz78zWxvocz1a2V8KT7betQJyBr6xNryaQ+GUgKKJzRMyCw9R
yiCV5MFkFT4wecR2tg+ko21HNcfqJ1yG7IAcj1mgUxGSfqpnpis/OvpivKHsIrEOPZaWMVbSaeub
HYJ1t/jJGpo95sBTem8p+qkAbIyeMyzUSReLHDprU78HeEexdb7HJxqfQOCx2MAsdo1rR/utQqsn
/nMBX1uofz4FyQTUE4PzPQkMP3cTe3UVtgHq8xWL/3J87A04knMP8Ndl1sirRDyVdBekmSoEWV2i
V80S2XqQxGrtObpmXUT3hSLAjw9jFe0nLhvp5Q6kBJmFkCQFTaPfDZQjoUCphvmRmDcuyrKfKiwf
fhff8NhRYB3D1+bFR5B+uBA40JDLjTsoWgn6d6fibovcxlus5MCBSL6oUxcu8rWXau7DNbHfVuS5
1k+KDppAIkVEX8J9+hILNmWspeFv1+S0DkX947AmTokZTdzNDpFJC7G/bOD3z/bfsT+PTS2yDTAH
g9jlj0/dWbqqHEcVOK3IRnQRC3zMraSozXuWLAy5kjOtjGc/kLj9J6SEAhMfpJWKUCAfrUIeqzk2
Wb8MgcF62KU6q939mzpQf4ybeKOm+2fpoymBdG2fArGKgfV6DS8y8IKYQv/XGXEEFz11x1ZsVS6V
55hXAF0C2N/eYBwDNeCYeznUbiKvm1/Xgwd6RVAiHGg24X+nsDdsS9jHPEKSontVpmsFzP8OhZiN
pnUQFqvg2T5kjRdafqS0q5gSKIrLcZbXZ5sCwqyA9yfOZH0R4dL1oOPnohV5vCn9xgu4j6TDW/xV
8ErIZUOXx1apTL0O08EXQCVIgJbPEKEzpgWizUWnPct/T46Md/6dFp3V7UkEnHFQbEkBSa89ATP6
iyuIBrNhNo3pmF8uXIg8/gADLWcx1IINWk/TpUE04s4sl+cfZgFldOp88LZvd3J/YaHTJAK467cq
COp7bU9nNKvT+iYEVcJB4DFgC+3VJHlazR+dKSN97OO2qPo1UeW/lm4k39YKGeoL+pQ/BjPxf6eH
G6Daz0xo4fAFvZOW/MB729KScgeHr8GQ/fSI3iXq1jhK+5482/lsgLIkYFzIV6W6r2+jGqCUBR3S
GbiH4S/VdgHEgpx42WsEDVZMl4nRTHkGzfB965wxc6y7leG9wjpXIUFwqh8NMFFCydQDbMsZYYzb
VbUkSqpxy1ByNWcGGuuafqtXSJhrZNmIQG/Br6JZOuqM7956HC/EL+vqzl0NHEGgSrvHVA4Jefqk
MIpALQUy8a0ACnP5p+/dUDZUyKFOP8J540FPhCBRvq1otr1/VpajanH8/jsxizi/DT/Kh9ayUpVZ
F0lxlP+HBeUd6VzngEzgMY0cO9+MMLBce8cRzX+SnCBQ7in22WUPkq8hJPvedy1AAUm0f3DS70wh
/sxT8/d2rkOGeog+28HJuZHGxzKzv9QWKekJ9RLLMtuBDhcDVGiCtUIz305pPVBxXG3DhmYC9G4N
w8bQ7WwMCd8u0E2yD9d5v8Lpx0dPKm+QnFKmJjFrAcKkW+8ZIbOdU8XxitNn4CV1c6XMBBzCmbOB
R2U1nBR5Q56EwjzwozVFLOykPMUD9qAzWPvxGF6lnGB7DzklopC1uuRPRsNzs6rahNLD3W0cLFIc
qtlk6qDSaKJc4DHBeYCJTfYvfO4/k3UttPzjZu043n4kG781qpzW6LdNKJpD5zZeqfYsnc7W473B
4NxBWBcAkbQUXab0KwXf+prhyyVCh8c+FwlVPd9ZuwumEwobV9hvyDgqOfW0ycDbAjSa4LZ2WBW4
GySwJMmnPxpa34L8Il8knZGFc9uUWh2M/6eGJayoaR8v0I5C3Vj1GH1sfOKnHKF4zR1ccuMqwufy
GE0NZb5iVlLumCX0rEmXGphxAxe+QSbcvqEi4zA8bwvly1j6YTsLbp0SG5lE3yN11KcKmu9IUFI8
ihhMDl4p6/dYXZ0x5toPpchP219B3tt++vcz84CTKnaqptbFN0HU476Wm1uu0xkJOCKWXn9kBinK
lKq6CalhpONSHqRvFVCPJtw5b/VrEqnE6X/3i9ixlR5DS6fnf9sr5gFc3ETMKQVYQu6G/EagpfRu
6QdV7nOXYdyHdGr1wBJHSHThuPMD9IgObyqqeMt0J4C/2N2273vMZF0qMz1erBYQOEVHIP7SKtxS
+Xy+wIZXll7cbqx32J8h71nN5LEPRt7y9Gt2PU2RIhsZEOL43BtGiS95EJOE6TCJN7/y5FfQjeOP
aJjM0dP5wrIAXp1ScQ0B7n7Yw7jfTeerVzv2zv1rcz2c8J6V4D3tsrXXvhOi9OcxMuxxHX7YW/SP
bqOVo/YyHOgIJcQl5e0YtQyCbvjbc+cXkPhblFOtAT6r7fhwu0nDvRmoBK17Mcwtomhye9F5HGmL
ks/itjIjjVS9axXCdnbsiEkJFVyKBSKj2ZZ6LhQ1gf8nI1pWwhSsGTYKyCLnnPcBfzF8GY16v4gv
Qj59XToCw0RFZFY4dtFGfaFXKnQy2Mct/NfV4DHjLetMpTFeJ3+9aRb86zlaeFeQZo0NluzP7FC7
7UPMvsEqWhHjet/zbWu30+5fKFobo9+Inwqb4iU4vHOaa3tJpASgITVAhUALzt4qBIiDnQZ435XC
kVNkg9Q7Ny5xNt/Z5U8AopxcwMPq5hxwQx/FaktYH0HErHEUqUkvo1SdxHUJBMXkY2FXNeTDUGhg
WDIw2Gt3TDgXU7dO92+ecozcjT9YBN5EvZTWOsrTw/DmCUBb5e1mKc8z0TSmdlg8k/db8rLmaNPE
MS1INA6grEO7S602BJ1SLL0VnUsjN+BqLPtd8GksXuGofvPiLcUIbFvpFKGEfR258dJKrnvJ0pf4
n1iIek6hrhcRtSmkXZjfSwXz7Iaq4jQ/shScX5Tt6tZYsV9avbBDs9FLIHbMo5NxlEEv736lZkeb
dGZLghyLeEhnzQBWzQC8sMRIkjnq43Ro2jxocK+wPJeZsgruKW7hAYFrLnWOIH0wD+r1kU1Jxmi2
DqkSsRDtLPj3TFp5O6mYT+DHWIEy5U/aYZOg/SKbaTMe/Y6rIyy3KaFZjQeXV5DcxC/KhfwbeIGp
U20RZwvEb943ipoRmzK0lUzHAR+ZY89t6KUFdEnDiomBOERyVTzGf2OPlkinsbjY6ZRBn6QQVBX/
snKUL/EXV4H5Hj/W+pDqai98z9hqlwD2PV3QlyFfXnTmvKvN7TH0RQG882PllaCaRcPxJktYVSry
3DU5/Uy4ceGfgwKQh7RsDnDofP3zBhwH/MeCHEwaRZs70cc+/spPXxepkhLFPNfWcWJIK6KqmWRs
LkGuNDnk6D50qGjFgav6d3SF9kL05aBjTdV8eKkGlIO41azvMztrVzzeKjP2gDxAddgP0tZIilKY
Mkj2qLp9BkXc0Ub/Oe5O+brL5TnYMF3XGHqLwN7TWGFroOXiv5yogi98B+r8GR8tyPPXWAduZerC
UroBLiqm2FYeaghFNLVF4/vPXypM8CQNLiDPZwBBfocG0ndMk/SiSwx7yr0q3GG1nznAJgzGsa5G
s2m0ITtRX0yRhfc1SbISZvZYLyNjn+DYqJ0QCjKZX2yiM4It1W30Ui/d7jxeWVkzPBquDB22A1Oj
O2ox+Cc+vDc5kGZIr4sjNED0CBW0v4u69l8FAXxbnQKfbjcgCYxZ5BBLMhNoj03g/MsrDBiPPItK
HHgHU0FAdSmxaQtv7qW+kWZOVA8d/O5zpJ9rDf+AWG+hxysvfGK9q3KR0vhx3cOlnkM+snVC6UBV
+9WQMefBR4YAA6rZL7mgGbmPSK+2sGPRKcGxFgNL/8JMpkN2faXXv+/0qHaZ/Op+6KISolhdEOai
xJ+4Ul2Qcm1dd8JagNd5ttUSeGh+voWC2uUYm0/e/kSWpyRPzELOp2NdjYDs4cxtjuld6Ke8f5Vv
xSZRpkez4/OXF1Kt8vsDtQzBY06rKH3g1Wc0TXFNQ7MWeAmpMqSLmzi1f9EmXO0JQIMiokfEf8ZI
FbVFHtVqnggKgGge9r0yPgjRmPfNJk3u0k3IsNO/ZdRe2KtyXFKi3OuGUfIPejE9bjkWMFVTYUCO
MTWm3T+TbniRSXgAlgrYkot+WvTMLr364t1YD11fOtr7h+QlWEcaaSRGf+sYSZneqgKPICByGKUs
p5P2UdUuG85EX0qKIMcE5032Ze1Qii1ti4X8XHaLSCRC2ojHsnUSV6gqq20XAyUsPufy4LqBBqbh
jhjE8f/M/EiUIC6oYlbLov1prx9T5uzyaJ62pJb/7kBwiJTAiWzwdczkV3edNL21vaOu3fJzgD5+
30A2h/5tTiRF02+j9XbvDd9OAlihT3Sx0rE2ySZoDVp9i4IfRy6MnC9xVb2K+iGwfU3yWMDfofLd
+GmIkNGK8RUS9ytMU9EflVDUMVeUZB1LrTKXYMSJLH3AhZK6Vh3Q96+4P3kKFDt+8Msm1hbsnhn8
A06gIz3+qCFLq+PJN+Vfyw3MNp79f5LZSeJ3v1s/6eJtK2kuP9iU9PsY+kVbQjZV1BrZ6fRpvLgh
sYyQvGx9gyNuCSSOifhxdOiVS6zzMaIjD8/uKdpyGnxTGIXCgLAxdzDkkFmva3O7yB3piPbzmEbe
hVPu9icDpkgBI2dAVN6evpBYK95Mookqfr/ajdtGSmC2YeJ3lEew7SF1FbJPwSkNqQs5RNeQhyGI
Yu1+0+3Q+iPhAzNefTP/YYN2VKy9ClcBBqBvwcJJSt9RzmMa6Ly+3Cx8vS56abhWdknE1WiqKP2p
dUjBhv9/NyQZsW/A6QoORKQKDXsOAH3D8gAdyZiqsA18O5w2zeHHxX0OBy0+4kOus9AXdljLx5Vj
rN8mabUHP3GmEAutfksMHoYQwQCshUb3t40Wd10fpNjzM9aplalALJb0N4nDd0od4oNh7RfUdQmc
b/mHRUp1Hd7QzMSkYKaC9sFm2mfOR65nbJL0fnG95LR3mh+b+sdm0H2S/UnigKAyjH/zGEj0jpwL
iWA7zOp6uZB5RasgXYEyDSAu5Jl2p83YA6peSEZwfk//sOBkZVpAkoXWvAPzQW1Q5Ahh099IExLQ
uK9J/hICEJrzZ2fzClJAWaxr5VLTE2dydSGPtdFDheLzk9INVQ3dhWJ+erTdDZiui5iDHpQ15aTM
/B+BmW7lNuiJ/KqDkO4vGMk40U2JJEcsDaiFjyVKSxeCr5uBjoVnxNnMeuuCDV44oQlZz8V8UWtI
HnMEBlD8eRWMo6V3J1b80Icm+8fnLopkYqC0ye4gLjV7JrbnV+BLs/zgPodQUfNH0daBJG4YAX7f
kW+DtQ/pfMX7GTXaMq6U/zCG21dyb/6WDAA/aZ05Gw8CSdKRx7B1DAwTCZ4AJj/g0X4P4ll2O2tV
EcDE0Bijk9xZxrONXvjfJ83u7+y7iSmHqYFNF90Ifw59clStYcmaveyokW2HhqpXNxHSPg7B4/pK
G/f+32qUraM4ha5Tq1f9wgq5KGANXE4TIJYWIvQLb95Xc4Xt4wGra19Sicye4llQNiG9gZBVZQOA
jJfshj4zKotsyeQCzuVaNK8hJYE/Sid8mHeiNCqle2TIP+2bOvuIlGpjVdYMm3dl0M4EGexUPuR0
QscJnUNp2YP7wVGGKDs9u3n2FtaODXwyGy5+kbWcc4URUcl87y2gLpSIBPJWuMDYq9yS66M47j8N
lGJwxyl7gT6mevwQ6guXntk+xeol9knc8HRyhdYBi2DIJ37tIRR02bSeHPLE9161Nxhe/tngCHpl
wTUpt/zqQxK3C8rWKv+78Q6jgn7NOiUjF1n1hTKgFTPT5dh3zEx5dd5p3kLnvr8RDboyv9aX00/U
yIY/aV97lBkC8a+sA48roAorXg+q8cz+G8+S8ZtZQkad2iQ/+NkScknZxT7z28DDT+Mj4PzXSwqP
DrZ5hDdM6pRU3CwpyEvaRJChSym6SZHvKdB77LkbBLrbPRShNFqRW4nQ/++UT8sAx/JWOj1joLvU
DOpfnKDbB1oDYgxUWxmiJwrdolPEQdtt13qiV1nBnvKXWT9jYDZdYLaIHll8X+wmz+GThpC1IBe0
CsoBix5Iv0yBWWCUAHrBuxmhhWc60P/MYY6HD4fXieemSmqgQ9ryzZSfCc//iecmpEDatafV93Se
IuUw/BcrQbY2TXeauFLAAHv0IyHZlPhh/VfDux5gBLBKmDZCMstEEidstxNz7v3hAJprTLq7ZMo1
8+tVGGBuZGHwjg/1r7LVblvZPdlsM3QUcVV06LdbPshOlu+eQU36+nmIf8QBZz470GgCZ8s2Nnl1
7YEyDzSh64A+bXy/JV2tAXGaD/ncEZwHWRiphha6LLLipBmICciwpMlOl3VjjgiBkM8FexfUzOnt
lg156Zu8m2VBky2yjw33/ycsLIGHVaRr41mPno74lwVgMSEuiuF0LLmUKpt9FQzkuoyqKeyd+Q/t
vjv4Ij3HIL/y/FZ6zcMYzVYqV2LB78z22Tbiq2UQ3vtI7NouhGiPXvzkEMvhRepz8WSB5GFzuqVM
pYRh4twSLaD/WS8mMzNwCoxSg96lqaLa9+spKLP52rjPnnkwtwO9KF3QKqjLb1nNd4Gy8xZFj3Dx
kCRJxbk/uILI0cKvC00emZDNksyiQ2Mrz71kozFADqyd5HxU5qtsfcOPlkNZCILlyzbrODk8DItV
sU6rY1A7DfaeDpCzCAE8bbjYSciEElR4e8PJ1H9wduEOQukHf/TavqfX54OfDbZPZfjZMnkG1vVq
6KbvplgZ5kB7SSsLe8/+hgjP++F81dibgaRC9IFiwe+o8hE2zXbBByHlD/iiOkX2C+79r3GSTsMN
JbbbAJ0NHiQIHAGMl2ZnTTDFQvcQBUsUm+1lHdtVbcmXw1jraQhLc1xvo9fZA4aRlS6yPEtivFnM
spiAbRTwg7hiwWIceqhe3j9w+ivt5LA8I+FYeERQfbWaZeTRi9n4Py1nwM5DxNfVMvEmKDKeU26U
5Jl2UL1mxq1zTyelyAOTDvDJSggJixJxUe99QYDzxSYB1QCi/A30fLjdv3XY3CC3FzpmxSRkImJF
yuMTkgpiVbc+BOPj2LoNHDYdMQlfQ++elS6C9P7iSPvtSJiKSgK9UP3BcyKNSBOegiYLB0x3pAPt
E2TaTglIuA09nJ8lRLXLaat6o68pbJD4VU396t6gmkPTI17H0p+plRO7sSMZ/dxrhQZ8kBjySRMn
sJUed2Srj+f0jh7N2HjE6999UhTZnq/O+5JU7sV/pW//vLpwGecoHzIE4NjGvJMqmE0rO4XZHZK7
e1OHPeNfZy0kXYvA13CigH5JmB/+htaPiRsPL0vJUQszz4H0R+GTu9zhXfNGb0sXx/VXaOC6ir6X
ZDBUttOEIv1IL/ClobrDxDlRX7AGTtUzkgrhWqGhcRTHDruaFLcfpBBUnTX9mt0mAsx17Y+acMYc
lfK4zTEaqae8pFd2FqjuS8SJQLgdb3FGS1HNAq8KPrmf1AuW2HY0d9hsVJt9tfVj1CPYWuSW7Jkn
+OeLpIRxlXHWkTdejf4Kkn33bbnspx4+QfRUE9uZ8/FVFU9R1YR9qkxk/FtyH+EsOUkXL6w6yufc
X6D7Qvd0xThfnGHwklLmN1Nb5PvlSdgqLWlIsS7klLwoeBOF82OfcnftHwK443yFfNhf3t6mRM/l
HlowLNeB/Pj/6aRDgiWRtDDspxGvUB4m2C1NCnm5oNCOAqvVUkREpUlWjqnAa46N4gWZixbwzPAo
MvRsOaL8/OdXXxWaJ0E5jpZ6qELHfPzgRbHYEJBxMkiPN3NA91YRgw9W7y3l6KrBXUpj13KcY6L8
gzCl+La55BEitoQLrrvicKt0dk75h/05nPRuAj6EuCy5BB0uAvX/PNGiEVNCudjl0rzDxFMQG6S0
KLOHAKAXekKVVwkM9352N+xA2hUKSAWiNxTQh6fAQLl19HfyP5D4VBsst3kFMt1JkMp6RplR2GBg
DhhSCfWmd3UiHilpZJ3MK3Biv8oUXXNvsztYE+liB2wA9UM00q/M+z3D1xtm/bYgww0vV6Rz7fsA
pF74mMnCJdOgMJmOasHyUu635JFSstxEGZymv6x6vYsX7D34CZsW24RvvSb3p2qbHnXj6+xSHZnE
lGOh9H1pktwOcT8MYyFv8T8ESWVQKbdRsZNPdDDdmr4IJHv3lTXuGGtUWaibjDSG02SEwDLJSXqe
2vacjBK1ZlDN5j7H11oCplrVMh+J4kvsqICYMBKlVx17qZLIMVoAG5R2lzXR+W7inslh7l1Dh+UP
GI8DCC4TZ0+nWOj8OiAzQVCEADRKgAIHfCmi8ztdB5fcwa940u+c1bNhYRI4hFrfVlztadhD0H0/
2gbkYDSTbjjwJYxExHQb9N8eNezUjxLRzNS3du8UGK1CK10wTbI3jWiAHcSFzWJ3y0/OcPAmsnd1
uvX9rXy2AqpkDKF8GsuhMHoBpE9pKpFNiwtXT8gJOgCBu3WuhXLrmD84danvx7sDf0o9prz48V/U
jLT2b9g6BECWWZKe1uBkesEEdTpFdJ8hvdFoj/4TQGqk31+SJktGgvhv6plQoaRYGl13cduEsN3K
syP4E2C8Q8W4sIGmu+gFfK3ZcFDkgCk3ppS2Ps6iMgn6X2vtQJy8oAIuC70C2TeB9T4qb/nTjVOi
rOQF86KtpOyR0F4CB2wlDzUx8qw3IcagOw65TcS9EboDt/HyFcxVZ5QKdFzd+C/INuTIiSzYm4rj
1imsvyV2q6UqvhU4MszTqKaLZQ6vIxBUZBybt53/QTYBW30XfQlRoVIaIvvnkubxHYmg8TSlw5z2
Fzx+zDA3wig9FUu3h2SUvgC+7yRPU66EMDSK0y6TghiLLN7zsOKr7R/Cy995K6NeoQuw4GCteKcp
g1lSJXjWjCpmJ1LRl1fPFRLRf3/dmQuSYanInIRTKcSfT+2E1c3GBOwYWuQLi8LwxHckm47swD6z
FUBEx09TrHcq0wVFHFnuFABquWG7tYKVZt+IBKa6C/kWpRdfj5J0ExYVATJT9fDFGsLMXyasySLD
3iG8zEfTMZhKi6pDazPAzmeJNasNyMJwT+PbXiquhnV/NEOoOnv/Twkmy2QzLuLj93c0tZi/JNXo
4efgEjV0OfU8QObF5JioeiJTaBs5KUtTvN/rHKF5qvBfrvNApXgAy9eI8+qyQoO8Ft7L70Fg3CMl
C6iqWkv6jcwGEjK+0FgU/VDLRT/SoPvSumMSp9W4+2EDtCPMgVBBtKHSAFt8s8bLlOGaFDZthz3Q
BL5rGXhYFOrrwTMPmcDgRlf2UuaENF2UlM2pceiYrHnGknF2SehPQ/Bzv4RefOjdTYp5QSoHze2U
9tLFzwNKLMvMOnRkk5B1QRWsHHC3dKgA675JXF1qUaLdrxyskVjMUV3LzAZn2zvPEmTk48hz16V9
vk7BkJWCntz1hlJWBoQ+OKYOZK9iCnW4yDAxIDMlga8it01fvdF0TeMh62/m5qXc4Q+ROYuUak2A
NChrydnq7yrHRbvxruwrcf8DdrfiqaxJSy3L6wpdcIA8fXOap3d7GhM8jxwtz16MuWZOeSXX6jXW
IFGsg1B8d8sbbzwz5f9hyaNMrYpz+5CqgDhSgPk4iSOBOP0x7jrP8sFJLhbzv4b7e21elhTDZS5F
Qv/iYmaDjlP0ij0HOPChcgRQm+RNziQPCXLDfP56VfV07HcdkmzS7St9fYDaxnBv81inBygPHUSF
dHSU3EIshWeMwueRIxbljbFg9PE7aerN7IfbkdqoPkOY3Vy85rZm+7qCAY/CiMhGKPV2xHkq2Cvk
1qlmlIaF1iGH2KYsDUhwwofkHmKP+8LvMJJPDdXBUhl4zTkaIAcuX2VD8tfmlKyz1RETX1qwGUSg
3xaaguV1rxcA4MZjWFTdR4/gzJCrVUhdEnZSbrKUaxxewU8uHKkHoxwdC/StY4f7F5ggxz+lC7UH
nvgYT38W1EI1XoAOEZeGOZ6M9O1urrmizSwa9pNWqu6H3RvrZqZQfC97LPjybnemmxyB3Sp4xCAM
2lzo5NGGR8I9yCMjKRriXQXVwdAwSkeIW1C/VZoHZgUg+bsze9XSTqJmSGgON90gO7s1S8D/lKB3
XHe8RYIBS6h3Jo6SjeSPBsQ66RN1crNOnBSdNie/VssnlT0Zb1t2Jv/tSpuZ+0QFloPdLjrsuY+4
BPsv4dXwa9t9fY7QfuTn3VAY8jeOoXWYCS6+0Bm9KLjEJa8kw6vk+PqwVx48U+H4tHMJmgW3cZhu
ssOVEMLuWPPKSbF1sin/xz6598NVh9ynTCjWsv8nc43uD1tIbrIVEk85mvWfiiB6WkQ+F3rJYvf/
sSlutmoJYwuTIqL9uEV7GQBT/FPrepd+mkLHuQIU/f8FaFsmo19p9Aj/Ve4pxyuhDTBpiOp2ssra
SdahkDIR8s/TvDLhT7cRE/Cf/9KfOL1Y4SOTCpZnqytL6zopzNUriz4fmgKkIIvTBqaXE51zvwyR
oNci+cuMyrokwIzXPqkestulkTKuIK1/S32CTD94NKQVUopLhk58XPKqX/74XNrxCBdXYDxXoYgJ
Dw81rRADZXffUKvbIR0w7bhOGJqh+WO030X2TUaCtejeex8tnAuJozid4989ayAjN987BQAbUKji
mGafcf4lUw5wi5EotpaKJhAuwZT3WpVvoNOMQFJwX+rqXoJooIfBV3lQBEUiTPR6yytwW5U5bAzu
8qYahmGG2deUNmdNNqWSDpauUt08Tub8RZGVbC82TORWFvHH/9WiNq+iTa69wSVewtBGAUDqLLm+
2bRJncIvzo7i1tq0w54y3Ip0gCQTWCFwxXWAI42NlpJuJVaUv8LOYy1P98ra2Uv0nniPZPJMJ2zZ
Vm00hg0sDlsNJfRa7xhapqIkA9ghZZYRgclxsjO1xLakaZ6ck/6lWCZZSyVOH7PxiOg+85ZWcbj3
Ut+1mjv14HNvCkD/B3M2hvcAwYEj72uFsw+CPvyr0N9LNr1TWAnBVzyrZx3EInykhQz/upTTZLBu
aUuFOIPU0webvgavO3nprlt8EK+MzQ4qO6jvT/UQW9wC/ky6/+UT6/RoHYbL4f1fsaO06so/C0r+
au6hJ6aHoLkH3TDQEA8VmjChKc88EYjx5prTl9WV+UkcIbHPyWexIplvWIoA6y+8c7adRc82reZB
wIR0ZTaeFZqzLdFeBN2puUL0jc/HD7GXEkt6tgVZvZ8ADyGBIl+pdn9rfxwiwrYftkOiVsUGLomp
HPANlVBscCjCuz0PXd5956yIZO0jF8/5nDTD8qfrH6jP43wSZVM4i6nbfRlUEo8eYqO4sIh7weHe
IWBhq7SuI2E79UqlneTHf0Wij5Q1ksl3SP7SpAzJk+VGNrP8U1c2N9+mg22OpnP2bA26OAe8DkAy
anntUBZX+ExvTEaqZcK5lgyXZruHiGHHS6BcPOT9FV4Hmf3yMFuKdV6Ya2XDVXwBQSPCQuhLn/yB
Z6xlA6gwFHRJNwwH0qytjO5eKLitilYZ39zfZyD7jE151d+XNMIjU27Vucx6PtawA4NmRZQRJE62
nAfylmLdP6Ev3ZyxHmz+sGT47AdVHAq9+z6V3RabsJM8v3G3KktPfGEA928iQtGc00pgmY/4YBWM
qGBmrONR5QAUh0JtOvbRBJdN2/qVZ+Ge4+hZBeqoysYa8iN0+a6RJyUC36D82kKTVcwYR3Mp6+is
3J4knNvKJot2z6lNyjrLSI5Q7rQJJcCv+0BcURWYURlDyqxbRV6EnbdxNR3XR31Owqf5slkiuOmC
cl1mCmJmyB0ESMOVPFAKvEQwtey1FAdxtnD1a4LmJkWuGPkAntItjLEb7W+3/uq0+8TdulJQ2m9m
Ukh/zXcgHEro89jokc9zT6yvEYebIXj1IqSFayOR7lIu5S0OnnoLQEQ3PIywAwy4sQtUrQgk7kIV
Coz8C8r7RX1nv6WFEn1CMoJoy+XzvZkvrbFDM9NBK/dH4U2wd3eBqfo7uOsVtrPdJZyt4GdZM1Yx
HkBGdugpiuZZw8f0ZzJ4b8XnLb14Xo6ORqJQyszzsZkc0kBs6uqP7NtPQj474xCKpDlAsWL22k5K
7xglEnvaoMfEG3qHWl07WfKuk9KLBz5Ek3GtEwBucEShzpcRqxIBcvKxwc3QPjwbTms5Lx1aUL/e
9ISwz85MK8fDM9a8nlQnQlUDr+u8beT0WtSdOAsRRvSvv7n0his8FMJzzN+qaoYVcEsxavF42dyI
eF+FRahHGXvW2cRwNWmYGP/YzZH4F99Jz8ZHkVUHfUnkeUWiaiRReQJTcMflV95BA1247N+WaM7O
k/m3N8o8sKPEIERnp/KTism8jmbrpVtcHHI1t8sdk1sEKPPQf/IUPDbqpK1Hfp71JecsOpiqwws4
ZlD1kqkVaI4M0Fl6kdrGkkhUWxknFIDjQhB7algTcGsGNLKaKJiw8wAk/s1yA9/IuNsJfSe+BFmN
vWf1Vdhyiix9vvxdN7B3LHdKMnbMzHSGHhluzOXxH2d4SefGlkWJHAouw+djFDrQoaSIaRMjGFqe
MYvQ8rt4lpTlYWo10l7QUnUDy3SIEhVHeMSc2mUhUurxAfvSFaS/hKl9koTU1D5wABUxzJfiIbkr
j8fQR//sKkfnm9Lwd7VzyiCKrz1xxiFyY4ly6S+NvPZWkcQJpGIuoR22GuDBZru3cpkDJrQbrkGa
cvAbHxTt0YZIuCNFsr036Aeet8crTfK3sOIMvVyJhB3VECFj20enkEY0NO5tggo9inbWpEy/mVsY
sl/T82/qVHkIbwPydQQwovzZ8Ivxm9nPTU8TJhRqKSOVmWut1uX+47NY2pgvL9+yFUvT0g5Yj5nf
m900qRraius7nAAT79IhgP7o4T7dDX1Hnl8+xVhzxUwSeikkl2MgyX55q3DHQqm3f4xtvYE5DpZJ
SjUn0UUNmaVYU1F54q4rMlLuAdZl+EMfse4wNrkh9XgyXKQcz7+ZT4xnJMK5CuaDb6cTXKYHKPch
cUTLIlMOSTWl0X72vGxFiMiy5scIU/PGwKpDlTNFPz8CI6lPKrk4eDWeqFBdOVHErZEIyduetg94
+pfMBEEzpkhWK+3GTKBDLNQKh/CuJTuXEQ2pI/p1lvfp31RAjObpaPEp4ibcs1IBDJTrgBN8UGZp
BT6SeqiWgW2jwgRsuKkHILRPZe+DZfQW6B0PSgefZTk16n72AELI9HD9RVrYRuvBXvXA32WRtpHF
pmmwn953cQ1zagHz0e/JMLasZFJidhBzfws4b6g3E8btdiqEXuWhivncMUEzE/EklrPgJ8IGWWXg
y3BFVn/Hc2Q+taPPTHkENDzaL/PCw7cxkOdwd8F5ktd/qXtPVOo/J2nqvg6UtrhdiXVth7iN4rn8
Xm3WF1H44+0FLAOgCvVy4RxToIs8Ib2Sb5nQ0JRAsOo+E9Kry6mnEhoGuW+C3UNROwkjwraMCan4
/uUWZzo2TxsWlkhYZzkS69kNULF6ylJ1imt8WVt1lLq4RTFN5SDSuN5X2HmvlTrUOOpguVDQ5JO/
DvMlxzo9ioZYP796M7IH7p/74MzSky9Y2W11r4a48/akWRkMQ/XslgSwPzqZfGrh570KtzGJN5rU
eLsUcrAjbkvHslpH8LDgBWehAp09NushwfoM99bMXwYqzkqvxElr+/4afqZX1yyxqXaXZP/6ay/7
WiRO+JJfK7EVsecYjPpjV4HRv5bBeR31AjibBKgYcEchtoY9Uloji5Bo7AWBnvtg5MCivazzAdi8
nr/xk8dk5nsnGgiZjPnK86GPmig7ba3Wb/K+cgpwe0W+OzmU3fse+nW0n4TZg2DzoihH1Y1hQZmk
LlJEPcTPOSGHUoKdMP8nJij8viksiUmDCV/VBTVzs1X3mWknAtusG734Z38+qBU4tv2SPsRMHGUi
i0Vlh+Z611hbxkaogguvTEHV4D4FXlAbIT34EC/FTJ4mMlc46xuBpvA2pCAs9fjoF2Fu9be3Pj7t
Kns4ew22eNKgGfPV4vxvXrJ53g0E/OZo1BZSZjbhuJDMAWxfHCtgv47iFp9vGAD87hCNn4DFWez3
ZNJhG1Pu0dTgPnZHIElQmCTioSjS1gy60gAY/dezXKWjP9g9PRaPotgHRkh5NMqnpFKdLrMezfdC
c5iglX0X+dVeRBZQBu1/hOxu3AtsL6kFKSeeDPPmFWl9ogE3Oy+4BN8gP4klYquaGK+CEbvH173F
hVH6Y7vSvZWEbpsRB1WXxh3YSe2O8BuTOV4NA755j9UFRPh0ef3aSJKgRZ0PjCE03hQiohyfmfOq
eJU/aFCspiC6T5Fnzaiw3pPa5bUextxDaLcJs9n1ezUxV42AZCRRRAJVDUgLVmuF8wGN4j1P+Lho
tEevw6Qt020wbSV0XayJaygIAGM7NWITNgCV471Hwgn5Ss0B8grBuz9yKQB14hijK3mlI4rR1C4N
Q/HkHDqCBbBs+NWlQzR0Oo+iuA4K0e44zXyhsSxaxDadX8XEZYGwbq14lfXnXFB0UhVMco8PBp9C
Ml2SQvxYmonc7SO6NuGLKQYbP/7aRqg8opk+tirUoVeLlvKQrw5ciLkFT/UB1R5p69diXbJDmZOY
X+YuxcrrHgDK15qbe4LqXCsO/JXtSZrtJC8fQ6YSih9eWTjwn2K7DGCFkkDfUm/RQcCQ213r1bNv
3mUtDxQREsL/rQAk6A06XerROgzVYH8luSJYuWD9azNLsdM0ikhWVrhpZC8ijACAeDhAiS+1bZ/X
YwuSyBzTRMqYxEiuI4vR7jVvAgNwhbpUcLxwE/dS2ES8HvpWPJOJ8OJnVY8jmH1qB2PcMeW0klub
E655aIeKakbAX7+uM4DmfW/5cOiiy5lOUlBo/nQi5XdaE+OdkWNRnIlzAYSkZQlXt6BHALR4kNkU
wa0rro/c5/hjKjKzSDQ8vH3hDhLELaonp9A2OnbB84SQsX9+FntQv+KCr2maBMAw1JtXEStLBKCw
GE1wr7rAdSfIPEkQ6fr6Wn/xeVjv8ckSbBDhWttAl+dEQYwbAHqBPvafMwO2O/j//rCMedX1sKz9
Yha4r6wefVwgZsNd+G/cU2SYg7Qys0X4DgHihouNO5wkVoYMFwcOBl6R/8EBBTDX6Htu9hHZPd7U
eptYIlt2tcEMY5rj7ZqEZ/Rwmj0Dv/jKbTo8YPVL2+P9RKbLlYjD/4cf+ptkxBxsrbCH6CEF3Zf6
n3U34Rz/0LGRVfbtE5yDv3U+JlNUI+GALEZCK5KEbc0/YoW9PLmeKULXo69xVDw/M1NxVRS6ILFx
U+0YUdeJJ5Ch57bjGIt70Dj2V2KHywxU9n6sUh8sNjIAMsipwGmAhz/E15RScTiLtFC6aganmu5c
pasvsanDEAotXrX4XXunGuUZYbSY1NmvuTdZjyThrNdnjnJl2+4tVhfkY+AZRIGt7bxG8PEWaxaC
CxuTxH77XGI1fN6QsvG33W/dhnmQLgrAlKKyVTrCKyD5yxpdlXhOfVIDIMh0RmYMpork6Gc6XvOp
zXKP0iJemH9cWNzmkA9OqbjlJMZNKnjpzmQMjwkmietXGVxlRMlO/NYpN2SoRwCD/vSrtFTTI9ti
EgzDwwSKBiBrRgdHeANNI9nhXEBX/Z6kwwOGsgoVajSLyB/eQWDLJonDXVL6K+NEup9aP0/ys7/1
qOAUa0MylsEfBgwpQ/4LlX8aigeThRqA5AMJikPIXvw8yP5/ZjHUrHvn0ybKrM/aMOq7Z0Io+bOS
gyMtWPxN/b6DM5KRl2zo2aalylNZyFY02YhDQ/+Q0GAwvffRUhCCVpIdBi5JwLQ73E7jynVR+XIG
Z1PX0ww6mNirF3QKghxaPoOrC6OkiYeDE9wnn3zqH+WQ8YZHCHm/X/xl/7I3z3L/tFIe7ch7lcvS
o0n18fC+1iAX8aLqLm9TPAHERTFFwOoWZkHgqZSgOVEJxrXV4lPEzdxydXQ0AnPcqrguJnVMu+bI
GpWusYHmKtUjFGw93ikoOjidNeX7RRbRiY/hCIzegzoTsAOjVgFk4MC1f77re/l2/tDAM8B2hmjq
Rxsq/iVsMYyAAO7/RR0xK9LNEdEK3xNCyFJ4WuCwnmB1SqOkfqlEmnU1UoNHCv20PSunXX+qJMFS
beEIlOrPgRjxFIb2KY7JPArN2ok1Hb7CK9zGDtbfj1C0oNzMgczRiPU1oWiVp2xqPDyYFd5+mcon
gzXwWY5ZZRJmcblegrrAUZma0Xy443SdP5IbbcNoYarxh7xdXwXohD5ZMpJx6U3AOV4e8x71pwqN
XiDZBi0oGlxjHuMKZF6ehbYkKvc6EJjdeshCn03jnxLmGMzNVSZBlORAcKLJCrCMnvCjr2fDyFXa
Ht47+E02AUZ0BXehpSVqbih+eyfxtVeZFy/ked7DgzREKXXPoSFsT7TRyuSKInmrmpZVOHc8HCKB
C8sqZJ1PAHq2TRRPEnMMJs2NiDy9xVpP3jUVMf8OOLwcpqzXunY7h2IAY/vbEKCglIdDiykdSk/t
SG0oI4gXJ08+xkytr+0o5tMXO28tfySsX2v2hvmHCzzX0EGiBlbu/9iTfW1PhSMZ9es/EDyMtzEG
X7sR/OK//gp2miUQdATvCw5/gKjyIMDgVFXVplXNrLNt5IjVF3UNCvXYxdEPM2x7cBPbK8IP4xX7
wZA9ap7+CgBNXkT8zlc9rXqcBNPUJX7Hj49tO5r1tZ+dnDOrSovtaOA4vEz4OvLL/pt064nclbE1
0RucE1nwXiFkhx/BY2Z5I+k+Cf9eUnFXc89q4esMEcIRsz+mhA87DJ7yR984pTb6UB/1g3H0gQfz
Mne2Im+x1qZWg8IrSmikl+7ATpnox9j6+FhQG8GkKDBRkMj9K9dXjHRfTIffhvUjFUnifzjucPzL
cUVMx3c6+bxVV8Sgo1XxVmpif/lB3ouyWGml/pfp6198V/JqZ7uqGnS6tSyZ1RgNS0p/fgzfHwtJ
W+FUFaUeucz17IRAlYGBi4xZdW2q+xEo7DqKzl7nTH3unS0LwoW/cZJrddnvMfj9HmQvQdUN2BuB
vWxvNikMFYsb//tpjPNHwWWuBqTS6M/8xJLTprROiAqwledmRze+Li4gT1mt+LnGr3iwmPQ24d6E
/IdSgOTQ+C9XLPE6CI+bmEk1B7FboRL5encykuneYa900vfwPYoxPbq4Cbo4d5q3FjQeHPZwwWEh
fOZJW8SfSw/nCy7fYzrSHnYWMVeRwai3LAzxu61T4lMrKRXc8XYl6gxa6SzMbvHs61T+wTifcsIC
rQGM51RqwQGSVoQB5uSKEVrxtY3FELshlxyMgBsi2cHNj8V8mtu7DSvCj8RLEu73NN7pg1i18tz2
eWLoKzFX8VshO5ijYzDYiZU26OM+LTsQV4kIxAbDRj4tfwYMwsOYBi+CUSLL+M5zu8hHz1ncYasc
L2R3FwgjWPAyUIY469iB79LhNtzZThM8DZOfAPinO2wAh5vAhEYFEcn3KOJrBfUX/nWAwSiFwzDt
VvQDs5OZ2BffkAAJ4Sq+D2HtM/ygriJBvL2s8Z6gXkiumi9mlfjCpsAOQzLqNrTFvWbExZhrh8eM
vSYjaTpSKPcPiQ6Ii9X4osmA26LZQuI3Exq01lH+GdpwLGHY+JrZfMcMsKbngGFL8g957/imFIaQ
ux4Yb4HAFem90hlKehls7Drux1yamClvEWfacidQrFX986g1/us/z20uRgL2rmj7tpK3LwipRbH8
9eJ1ts45we/1BM77UeFqxycgFvJR2QqkBsucEYHTLfPBzJxuhpOgk8jqTbDHI1cs2JR0qghatx1T
sUqLOnIs4Q/siDhlcer3PK/4TVqZ1sut7S0hxEba3DscXE5hG/fmP+rtcJsKaRvJ3rI1CdEjsLhV
I6UEm2eanH48Zfh3MuQiLYVkT74p6MAwlK0zDXfjXcSfeUFZ09QIfGUahTevFY3SQ9ID9qp83j36
df1MnCmQ5gFlvZ28XYPswyHr1ColXzXJzdISiuZ+TE94D8I7yhIQ2MidFalccFB9z3nG6s6CvsMq
mm3jKQ+DmsN16eq5CjU14Z0hpvz7BsKqmFdKaCqKwwaF1OiW31taZ/q6rswueZo9RkaKWh+Irh/6
E8f2bCZvGk92yBI1ds0g2/7dTc1HzpnlSzbg2KQu/XTSL5Z4Gqgkb/29JYJ1+Od9n8L3T+sgFfEW
EzRluO+xd+FLem8p6nZwWxDRcZGSm568m/33aziHJ0O/+Bb1Nk7HCSvxjqWelCseouQRnQjuYbnv
VNE3ThviDppcf7II4udbdrOFNbGfe+0gkQzaVAAuvyrG1e8/8pg6DR7SlGMCfr2iUlw5Zstm3F8H
Rl/P8cDQI3RpUzp8hUKGCI2Ms3Ro/DqF0ZAEcyVoCRjwd+42rwO6jhYiOKYqM3l+gvuS5l0Mn0Oc
O4gOh8z+svkF8kDcAQW5tMupwQbXSoaYtqeAcubD7FfYDhjnzGavSHzFeREV6bOIfSPLn37toNQl
VJxrpmjaXMr7wdskjCpFfOL0pF9BuWPYxyDpVpi3Db/TKNpVCfSAq7TH1V6ObFzixcya1CwmjekU
WrkM4z1wtpx4V/D/7zwalU3EuvE/JdZqNoPUv8j/xWizQadrODJEFIyOZZn6D6shnsL2BVpoAbrP
otujWwNIU0fbGnmG2E+HzAQe/ztS7/rt0C7TuZdWwr5MsUd6vFc7AGawTCZgUbwlJPUkLnwcDS/A
lOahGOAlwEmTOEoSQaIG4uCz/5X++J1vz8G109WYbgSMSWPUJfR2quWXxvxgEuLniw9xjaACWD4I
AP1PllM7FrCf+kN7LPECbPWKITNrrYr7UCCX+wpMo1yqQHeOb7JZuKmP1gw6dU8hsvGrovn/Tar2
OGx358xQQKe+7N0RfSMRKWMSCUAjFiPVGfjvm6Fa10KUEd9lvi77rHfwJWSZMmU15NUH+G0X1fG/
zCrffVx8cgXOLY77Z3bORB/tmQBQDb6Tno7mBDgInReOzV5xotD1t0KKllmXt/qgsMznKVNxIlj9
SPwVb0vMr6DwONaUa+Ngj0ZB4c41rcBc3r/ey2IUURvTgAxOX9olSg5VA61BNY6LgY4SydfP44ms
fgNMxEjsFx8xonr1ng/Xq200wUoY8tug6xFSLjAHRGTb/nQ8zKl/X1nOR9QkxOh5BxWY7sJaSzpV
pWkDqe57+WsVsfRaP9fAfbtj5ewhm4TKiYuVNnsAWey2W2VkIg4U+pNLqPzkCGiRlqgIybTErAeR
3ac5REB8Zpz5STXkjEwo0pijUZnU+n5RGa7qX9uTKicKudyvRrX43aN5ECxTJhnxW1by9VAUuCBp
iep7KW3GBxntovqvkQJJ9MF0HdvWoZy7EvvoDgR+P6pG+8+4TOcHf8OK1TW6GzBjYZfvNz1ocUKE
muDE2rsWHxl3PCk4v7+XdE/6MBOCkpvnj3pSQqTVWQGD9HrzZXq7xLJTr3tNXkMPcibjoDPtAB7T
e7FDX0Eto2ZD2e+xpLlxCGbJXPz74tGvqcQA6FNwyXHT6k2l4l/t9Op4KePHy9TIyPJiflwvZdEn
VEGEBeeDxayumyElSoDGIYRNVSKRLYvbgypQkVl2f9qHBW27jH2DslxU7KrSfR8KSEVJW6eCQrR2
rs0GbHPhK0NlHpefvLtZ9t1GXZr0RyZ+p63xZaOb6bzOqS6dzCsblzCSZnZ59qVQS3YuwnMU03Vi
hX9qGSbxUi51Mftp0YoxNKHTj5dwdOVOyGwQa8TX8F0zCTL1QiAzYojkcu6IZ5pL6W2kD++0w1+f
HsweH2JlBPCVWqSYZbNrQemmfLmk8NrnxRJVB5Ya8E0v6V0noh+AKkKRYt/6lprhnWIYGv/W+boj
g25a1v+q7aavp0CZ7ZLYKdjcwZp+7EBoth+3SdjXNCcWV6lo1Aw8E3J2f+6sljk6zurAjHWEZhCl
6b8bStCbyO2jL/INfJ4RawxIrU99uT2K+eJ4a9/w+qRnlD6sPkI5rp5UqRd8FOKEiPR7ogXko1Lp
Hn9+yNgtxpxYc/+efJZYlwH+gz4IqYDSy2HgPgDj3LHa8MlygQrCTT0HuXaBYqP12wsVkx1CJ1M3
9s9pq1czBh9a30xxSog7rn2jsCWILpduIkP1Rby73ngPYGHAWZ+E7WJtpA9YXjpsVs0bqPCuohsV
AulLpUsrSVpRs74j+pkCZ4TBb+qJFKVX701/9zvvytF36anI2vG27XYIivRB4lWmQubWi5dzFS1G
V+8PbayheJcHQ1jIviLbTgHOnmbC48FK4eGO+tU6zLckOevFyJd7Xywoa2z6+p0d64ik2s5dvVnu
LagZJMNUyjaPzaP9bnoKGPq8snW8xarbW7wLUvN2AKxoqCaPcl6oGn9grsHGXbuSBtTMsolT7FMd
G7yNO9JrapulseMBpIDuPxJZJFroWmwTrI7hzuU+G2GPZpQZTwqf3LZ8mRVaXewPuFjoFnCBsiuh
n4k/RUuJ4wq8v5gpfe4wNDYjpQKGQzO66pB+r34O35JyEj/xN3qFiRq+odIXGPgWQaGQLGCWtM4N
b1vNaKEYahRxnCJaDMT/h5ED5p5+3Cq9WiEBeCVAMDHt/0VXQaGBrwKs/L209UCUOU2XNkwz2w7f
2NIWp/TVn9JTRgRZgj0rYqXzleMesBL+qDKtXgvRo5yjIgCe5RqgFtQorJkCqonPseBXQUhzIBvx
l0qIgkZuxi/lKyinJzz9GgYCJQRjN0qzHTgiLgez5jowFPXL9V+Lklp7Vxf4oEvAm8Mx+gEOBKJc
LL51OMOx80tIF6Q6uZ1XkiogM//18sJB8GzvXUjlHcJVXffBNVt/WcBoTYO4SM/NJlte0n12WS+S
SquLRYlq24YPJ3l3ieonOdYsVKRCVi3hoDLss0jxvf4JooGXCLpO7UhDFM5rWR73nFnD6qXuyZDH
aAkvYnrJ8WuMwnAjizuqkUzoT74b9O6Zib1vfqGO9QNFkWccyzZ83JutRgmfsXLc4wfumZ56WT2f
LR1GtlSctplkfSi/sjV7jSfnrk5NOnX5rKx4UJHlL5BT/9zBbj5ip9pQb7pwCSFgRJQJpMxgJ/aH
0fMGeSpK5UhBGsQxGboHTQETlWsmm9v5vZHnqVSm+60loTKDy8NckwuFuZoL5gvcs+is3HENSlG0
ROxrROyHjtZRaJXmr3vGAatj2Is8ES+zeV8+xErlNuRa65/VU0h23YT5u+BH2Jz/oZLitgi4umCA
8Tw0AKho7SynEG2O/O6mnOky3QlxLowp3FqSCxyjn5XSmqQA9hmlKzEvKZZIZZjFzJV42hxA4Iwt
bjKsGOkrsdjhWwPkISrMIx6JN7CFLkRr12tU4uXEMmY0BP6MnpvhGlKMLuv91RCIH7h1VemaKErJ
xH3m1YFr9osQ/Xb+Z9Ggsyxm/4TdpAivrShb6QMQO1Rd1jOyOJUNIM7UkID4RE0Re68RMg05YAII
HjQBfCftPMZMeSirGsGTdk8AFbJX2afyaXaKcL7ttYjGhwdNXoKtAR03s+j/X/jaczkSEnG0LHLU
Rwb1O08pPqAbWxiB/JO8r+4H9b/a73V0xPN20ADkj8sondKqJjlzbkrKNAur/nZAjGfCZciA883j
W43lTBynI0BMeqWEXtVV1opRApTPic9xcfRykrb4KJ415+LWy7z8k7ykzesURnxGgnbDRSEMuuvl
ksL9HE1+qzqXwe+CJpXPYEU/LC2OZi1jw49r2RieW4GlAzbNOs+c7nOOXg6BSTsaZZ67PLqs7eRe
fybw0gf7/1DIFZt6AhIDWfl5g2ube1A0QpKoFmXD/L3VASAGb42mzBl9RVCGkeNjI2R/GKfQPwv/
HGlGQcS+GeW7ZrTTrJ0l/kqd2ukEmnIPgaXrE/hjhtbb5utHvnh7Qe4kM0zsITdejhk2kfpg3KDt
YIkhQRZBATXramT2ITTod9ZdA9PK5toSR98CwQiYIVThDo/cPCzJ2/Il4UhqBSfQfNFoI1x/kMrC
qapyO8QWMJ68MINVDB1ExVhN9LlpZdDqLAEbZ7/yoxguscfiDToAlNpsVGvbro7f9wgsJkRAI/23
0zyCW1eO9AR713v/WfqD0NHY43aauxRxPq4OttQUmB3uJUpHrJ8uvPOIVo7oFFvQYn4bublOVa9r
17Bb5NQ0GMXhtQ9u0iwZ+BvX6VCeyaQ7mvA3XEocxSaWNrxA55wK0tE6igs7avibNVbe6E+NFLhO
o5oSsrwOBpcPp6m4cEhdd9P7t7JPw7TgfptpkqRhdVz4aSbkyN7wEka9FEEchDKXF615SbXqaxuv
knh1C6QTEZVbuPIrJQpJlIW7Lfx/+VRr1nvtwp94gWcnCZ/5Yf6p1KXkMnTnfyR7fKhSeVflUa3r
9i6eu5hHkv9THFjJjsvrOprUCmFvbU/cstJdy+Jp6P0eJxOA//AC3B4BuGRrT33XD05oXVnmC887
Dk99+QjtJ9nPrwI/ILWWRwaoaONzlTvxby0G5/JSdeRSAjpJTaJkGsw5pM0pWhFoc8lFBbt7zpof
8GnvBF+qQPiOtzzsISDZL5yCrD+PsktpHnj8rf+DE9OQ6/KeeETfCEDJnCneGOdR6AOrp7md3Vs8
WfWMULvQpM9hK3vonUT6mnc2fVxJpj/mqstF4UcciBtcZygIp5I7Hoyw2LEOCGNMHoKTLVyvnc0y
zR1gHeJKbkPSdvdDurKRn8SIdrP8okCdkzJEdOdVr4fRk606C3ufgL0FFOI7NjRitsn1cYvfXYZX
4nxCBXKC2VL7yMHcPQOoVwzod0FED/i7nRY4/lM6yArgv23BUXbDoSbdTw+mznEtw5sctJ3U3GSA
bwtyGx9+ZwIY+cXIx24HnYXuY7LRPPtIW6V2EjUjoyQbytAorEdTj1qhqRYIJJ9eDXbgLwRBN1RQ
icEn9RDgQu0g1xZarXccpTf+YgqYdqBaRT9FTy07XM2054BxI3zga4BTFuz8COgImeoKHZWd/g8x
DnFgLw823NPF/IOmgJ7DGTV9/FAOoHUc10D9DWFbGgh9XWT3NDl/veidpDd2acFqkRS1oCg6t0gE
/0C6kZ1AaBu4TtRpA12VDnuWS8mJcCK5LIrTvZn+/PhgAvtn5hF0AsP4i9UK7zrtOZEDhSoexHvs
JovVJMB+CB3OMgmO/J4TFR/nrqHI9LJ6lfGM8a5w2ilAnpJ/ro+FImpVH8bIiN/9R6XMQRFIC0Z8
66uQuQuy9OKt29ioPCB/nzbd2OqK/4KvdTgjIfNlS1oW9U3ZO3x8sLiF1z8WjpjVNueQgYq61ylL
MyHoFkvKhau2tgxvd8yd0m2iw9FsUHMJC9/kEkwOMzSNbXVsVzAtJCS+4wbEkIxq0aPzYhBxIxJA
M9TNKisHOEZzndVgHsGQINmG4hlsPFx1jIoxSNZKo0FaUbWx2t19z7ir+Ml9JaykYu30CGmBCcgZ
IpFAQ2Pll1ws5wSvgweraEY242/qR2IE+gQ1WaOnBr4lqSfgUNDazTVngTL+TPJnXNFqTZmTXRSE
dHQJpm1+wA2zGvEMWSJi9qbhmeupqomNgaQIK3h25mjIkANgKphoLhymHJRUNNpDHln+eEB1HIpq
2KW94cQ6ipWw0OZHhFXtUYfPJycpFhjciHbfDG+cwdq4i+4tVva2veNai7abhCUbQxCnNiqQRW0S
VB3P6b1OKvjbGjFqKQ8hzLZ/gtVNoxXuQpO60IOePuXBPdYBNCp5pBg78YmvQoYcOeoO9wF/s+qU
1WRsPxTD0rCkvz9rZ46i4x8lTTKk8Erw2VQJ52ht/jVIfVVyLH3Wp9PZxE4jrKD8Pe1WsBH94HdH
s5ae56K/OsSJamAi8+wC7ShnWs6BoOXze2bemUqueaqz6Z1eXF03CgZ6nf4lrbFRJRPoBTl1Ibdz
QYCrZHAkXHuPr7EU7rQAayRhCS82ckjhEMoFVgfqkjffc4cmB9XNtAPcTetxxXBlNsXes/eA6RE+
9qtRE74oDtABMe5sk0FCijyxHLqrDgvKwbCFRN2Piige31mXwBcgEtsjZcFAHGFT/2TgSQJAUXNY
O3c5pqn1ghf/+4B853+kuiBb0/G/d+/AjgalsqBj37y3mR8l0p16C1Z9R02SLC2bjhjTQHLfUv68
x7NPB24yT+forIZbFsWlsUq8KAFzAkus0j4jlZr0Rflxul3PlshfwaEr8a+opMqrvoIKW1SRu8Zo
O5ZtgyJ6szbDrTJexnDgh63uYa+EzfLqDR9okHpeydgBNDqOIImWCrMcedfPiVn9X463pGjxliJl
g7mtU2FHERsXF+gXyqUioydkp5Ld3g41WSlmf5H0bEr2CNVzWECT64G1UI5hzFmFDbMlraNhspNp
vs/br+Zqd5Q3Q7lnzGvY1gs7tJym1q0R+3dPQ/rhK9ZvZJeBKhzCWLGfH9oY6V9o6jA7F6u0yYzp
8llZDx5O0fg7ztBFwkZ9mNhyCfpMNsAqgLpr7vsRFmiZXOF3xYQ+GrSJJlKOZ90/MR+8KVkMWjzq
7+hOPCAF7k79einkq14f7B+05F/c1t0jIow5j1KaHG2thGhsWdiRJIwW6IFlxzrwNdhunu4tmGMk
foknYtKPAxWIyqQ7xSeWOm36P8zbHqd7RF/IBspGi/xRITE8fNlt5qBXAWR3bQhFro2RqfPvdc1a
wVZTf8LcYPRv2uZ3pEPfJ0gJyrcWnpvwBOT5ui3KrGbAIp9huiKwp6tGbMvs9gtyBvL57kq0f8gW
ChfqpsvJwOPwpMERBh5OTpLL2oBATbix63nNOPsIiDaLEySQUxh9Oj84bufaqK5SBpy/qJTpvq1w
qhog5mFaSURk6NNxnGNXxsUBYx7fb82+SoidYLaBsWNVY7lfb3C4gLAu7KXzRBWkP4HhbHbvV4TO
j1hbmJiqPNS16aWWZuVtODfddHUFvaSwLSw3DhovxQVqL2VBJgWQbGg0AZsDLVfXSx2hcmTBdeYz
R7F5PXeyiWHyNSHzADFAFr3x5rIK00gKuo08vKWel8r02JLFy8fkLBnkkjVsvw7dpMq+ZJTKVJsQ
fp23Vz/Pw/zFnj+mxWJplb80uiSrKP8OErzRaV0p9uMpDf/ioGoC+UKOlGREqcmUpqIgaqc+7Rnk
dEmTwGNXesCIT+tBeUhy1Aek2zI+b0LVJ0DzrQpcACcyh1YPjyf9RYbnQJeQ3sP5nML1L11S8u2f
0Oa4WOuzz83mWz2XsJcFe4sY6pyL2CyOBQ8hE0jwmcC0on9q0NLePwRs811u7pKwo8nURvOgo5rq
fBYUD47EB7EXCaiMdZKro7dvE5xlHCrkZkZOSjam7FrbZ5Dm/8/tYa6pLX8P/xu6hh0xOLF5BaKy
VOjWJPcYGBA/52k2tvctFQ9O7OoRMax2DtMfLvgR2P4OrlG4SBbUrVBJfz1evE5d+beTO2hjowpp
zpgKInixrOmtjr49Bee4tmlDb36C8kIePN68l1iCHVQV0ILRM9EzwdhvVcGP0PvK1Cc9Sol2J8wO
Ue7A1Gzs1kcIDCu1bQvi+Q0qCs/re+57W5JlJiByhgX1DrO71X2qp7f+j8dCOenlj45KtGYMQMNv
xwW2v6tsuT0yIEdyhljmD8NEFOgJJ1qI6Y1eLecZufbVSZ48NR7di2IV6UeDMUZINz5yacUuKiuo
zrqvIjqGMsK8bsmIU0CZ6XQkDa/ICGeA4pV1TdIDY+FePUZmv+SWIUj6hVw4HDxJyvPdZwAtQ8oe
iDYSKDuI4Qmte2DLcU+bqEsOqeA4eGoAFdurrutStM1IECv1T5xfAwx5mcW2uI0lv25iXNebctJf
lILRKa31uV1/dMSNYz5rz51FanjnEYK5SheRa66wTctR8QV2g0cbcouLfPH2mYIVYba1cWsWEf/6
qlpWIRe5ZX27HWKMDSB13DFLu4jMvi+SQyobMRFS+IunsBta4uvGLKF4CfbvRetng9TbCQk5WzAn
HtS7cY5/UE4gbesI/Jvb06lRyGMO/6WInW7MyKfzTpLj3POCpncC7OOFRb2TxO/tvi+AOaR/7v83
ug52qsM1viyh/b74R3yxy6iYgCEsvAYGb9gylbZ8AsgCxEvhNM00KhQhVqZuQeYUCq4bOnFEujmm
cQ+vYuqobOZ7NyADprtNrYdj4GNPWa9yZSX5ih5pXGE+WzMnH3l0RXWDlFF88Sv4GqVlStDENzWd
5loJwsosE2wdeti1fZsxjok/XOodnMI1bk93UPJcLyOYmcZUlrxgqyYLDUvomPtAdCTy+I41tm4P
BJ5M9X3e1LC6ALRssYmY6kYcWMuQdFjzRQRT6RrwvtRa5kHGKQ/NfP6V1tnEtiGT/594z3DmuF/3
1frZUVcDLVXtrFb0Fpfw+Gfz8s0jYyQGdc1FY+LgU5aEBp0ueqNkvXp5lqC1Rp9MALlw1xL6q8/N
pk1G/MRz3J88+OT5rllWhBFid8jomXepkuSuMTKucNKq+UvtwwAD67UwDq33jjdl61rWLXmKaK5Y
a8f5ZX5xqTdPXxgcvvQ3c/chC+/lGYb8+nJm7UbqOp4ZQgoalFQJWQFSfS81CbYnHMzyh7TmCJ5N
7RZWx4UvTsE1zXb4kEeYX+GMFwWaXTBnGqReMNAzpbNEuWQPFv3lHodnOVU0vHICg63DQCgd8McN
Rv0SdOybBkxbNpSAeJ77LTCNmERax4n2zu3jwdKEM6yR69WzxiKzkMD9+DSpxc81757ZPl37nLdg
kQ2jlLJYq9Zh7RMksdqW0njSy6AZJzmNBgNrcJ/8+IZ8GlmN6WPTS9r1DdBLWunpjVpdIuoQyBUI
xeGd2s6LkoAj6bPQxrogykh6zKEK18WyTu1N/bjAERfq6QZCcxFDj7GuhG0dLC1rj2ObqTGjqik3
qO7Om7zOU+HIFGljxuPtDp05iXVdSiE4E+SQ4DwcSQs4AmBAebeE1yOWlidOEUjolIt0hHO/oFoW
KjW2ivVtA4tZR3uJL5KOkuaBxg2j0paZYksd5HDJ8MrVCktMEJ2KbUQ1NFzOVnLO0MXViPUsu4wW
R9RM6L7Ou4TimyFxxzhVenir0rd6UWsLxHQOYy1dfnX1cn55EPQoQTCWVKa1EKxZTth4M2eKb3+4
5Fw7mEBnG0LWbVyIUSFtTD2MbfGh4rFAWibw2qZqJk9EqlMKn3cyTR+WcsP3E3E/9UGLN70pSzaa
7DNUHnFFaPEPPbKBc1hfyK6dCztzKi37kmzHUy6VI6YT7PjMmk4FPw7OsZMrGsZWd4y5AckaI1h4
1AF2gbNyw4+zvwnrJWkxKQbb0ruTxkoCMp4jladU9EyjHwGk6ZIUI9hUq9WpOBh4wT0Bp5W35Sl/
XEsfG4WC5vQTZYimcPbbO3sD5K0l9jnxRmeq9A6vnyd9tSGSJe6fHwqNNsYQH+3w71+XjLvTV+07
UxOUxAJCw9FS6/7Y22NcHGKs/4F2oUxByEaml05QqEv+fzoGFVTcna7bCMI32PB+voiv5JF+lTYw
bo8RqDIjyg5qnSmx1DsNJ5YE/JL+Nc6eFjFFfh+05bdBoKr8KfoXnNgcIAzkFiVGblqFG3M1PLH7
MwSiE1ebAM99SqIgtfsS7JB6r+leUfPjQ7cs0H0jdBgNb2KyK/r1Dl8a3difE/oFNrjiirL971gi
cHHTzOlFxybkmfq4s7arZ1P8iIH1UdMbB8WyxKRItXs3kNFgfVKSuM5yDJrG5dW7XOaCjWaiGgsy
LeWvWBfNIzQxD2k7UIh0AQQ1CtY3xaeJQbZDKr3kaLkoTNSgkM3OwSIlSV/05WIBzwlhcZ3hunAA
sBoT75PrSkLAZJ5ngm11+GJ8p5fT2Gn5PIRE/XnhF5BmKm2OkxytZAKlX0311j4a+xGlDHWUV6Gk
Ia0Pqx3zS21rX1ohiVT+xKK3O0SyR8UbS+N1vE0E0VMdFz687e+ocGEhiGIhtrjzZ3aVrF96xt0I
pKe89WWxHE2+BvKwTIBjjVbFmnKtzFqdXnvfDeUuOty+LBHWRMJiB8LEjwzZBHM+6y1R7uON24+7
wok4zBbIAU14RplFBX5O6sldbpFZSh2qy4u/hu95YdGvUTvCzg+/jBIF1bWhOeVfdtXIvTdjEwlE
3FwJfbszN9O+9d5JipBEKSEpYHfF4JdvtSSJhSua/YPXXwgVoqHILrdgCeOBleOkgox6uB04NMST
/rBoUw+GCC41vo7CQOcjsF7JZnEfisQ3boWTm7GP/akznMcz6yciD51ul2iITv1E21PNBS/xRzNy
zAcC9MyYso2rkEA1tRGjP54zBErvSLhS8udEKxhhaUPAjxNq0OfNlVQg9z7NcZCgzu6FMQ6OjKOc
YC+sdW8QnuUyqBs+8dSJnLIJldFPs44RYuO7NFcK2UwNPb/XOvBOdEd5J/sI+gxgvxalcmgDlv3F
AXkB4//OLJiUZ0LYdYdvgSy6TcKwi2gknnkkGgh3/2LVRwmuGbSK5tvaEIXMY2/LtKTiwtUFy5hl
wdPQTQ5lKy1gOJXPdd6VrXKmvWvbUNk03Yu95C11flUl62yiByD4M5uDzruB2MRH4c3D/M6FdY6A
9Tw5NyJcP6WUkQl6Meq+2gU3p+RY5G5h6drgAQfP5SlJoTe8/ASYeshDcPPPrXeA7lvbPiQG8vQE
fBCc5KHOLT/aSvLLMj7/sfPYt5pEcEYM+qZlXlWW4a/QjTs6C6Al9vntV15oNE78WhjCGDS8v0kP
kcOLMff2lxAOkG6lX7ZHdFUSFuDogOQRKcYYwQJIEGnFDtWyS82+PkIzFktjtMQ4fdASAJ7wVhcV
r2HjNwg0WXrw3tTl2v8ohtOxsyQ4x8Kg0CZb3l6n8oD50hFlu4nZjpv4GSjy1Zzacv4J0+vFisxP
hnj/M74m7KAAQ6zpez/3l0fBCZ5GYJwX7yN0sYFFTzS4ewnd5fI4QXsICZwzS7E1R2ZET6gxWaxA
CSynUsumNfvxQZ9P2T9u4oCxzm5umXp5AhAksqNjDWy2URpOtKGILpfsQvChOTzQc8+d1H0sPH3X
Z6Te+cZ+x7ZsV06maa02VHBjJQlPJlleOT65YnViLh0QlPGuQ/D89ZfUQMC7taU4fEQn8aZBrEYZ
/EOtOk8FcHdlINuspt4TZg+gycwfazf47ggVp8QI+8Z7e4czuZYGmDT0i/MzzRMKhg2uUvWmWnoU
LzI6WHd+RGPDJ/gTopxkmxnI7+FL3ocZUCYGyJ3iUqfyd2aH6hP2kMSF5DN32yqY0i+XH4FWogCj
iCNQinhnZF9Tqq0kqBFjlyxCbcB5gIGv4bxic4lNI0N17KEq+mcWoB68FtRP8Q5Vnlt/oo/SnAuD
9q3JsWkDTNFCnaZLYA87q7yw6TxH9nDArTPfcvRQOerWh9vWTTwn/esdfGKfiv0WzTKj0GIYMTKA
W6+kKmb0DzhzZ58IDYBqZitVuaSPrXW+h81RVgQ/IFgoh5xdygu7YK2CJQrncyBOsxCJy9AanVgK
/wEUGsStdlbKHdhItXKqLAaWnZvIPhTqKQ22pes8mRs2EOiEZsn44Dgi6a+DdeXkcQJm729AFvXS
QCdaWS6xcBj65Lc0abYeoyuDCnaLu+CQZQgWf1h+DamxxSwl2HCCNshGezgJ+eiVkgT4vwTkljhC
+QR1Orv6MfqwU/p7ZPYUwP0QXBsWXdjspaUcMpqibG3S4kPoYcOWaH9b6CnLjjGNFgq+j/AJ+5QJ
NHl27EtXo+X1SInBKtXSJ/I+Y85j3tesWQjMj/na997q5KgKWrpGRCPnJnWBpPBpk+DW+j1tIRu9
kBvDnluUj4LkWEMSwjrjeZ3//38BmG0yD5PPG4UvoOUH50vpyz/+sZM9w77GOPDPOJctAhjgJYBZ
YwhEBQMl9ZCjKI1n0JdWUcrPhaz/taNUMuAWLYzJn4uigLJZNJnYBkKiemaOEEKMMauMQ/iLsL5/
bA92OnuCzj+MCtWG/VGxIK63AmSl2tRCePWLK2QqvZi41EZmpjGLMeiPAwvkbS4TauDdkg4ZbgJ8
RmkplqCr06M++J2aJHexUVI4SNlNvK+DfhrF5bU6era6QYa5aXuCXQIYZJydhUxH0YggVYRJcomQ
1LEyb58a/CMKmqjn62yUalm77UpaSbqcU2INAbjEMwqomsr9zEcnilvithKbBs/EuGP+nBb4STba
68/mx/Qub33x9kwU2Kb6rvJAjFfYBRFrQaTMX114hG86Lig0JCQDlWkOKGIHdSeBVVZf6NeQ8OVp
+ZAelTKo9NtRosKonxuVFxNa9QBNfwjnXCH7JCV/3eenpyrvYcEHJU1NPs0y9qkfY+RC5VgnhxUe
Lnhm55XlZYJQGLbDjQea+ilkTlWpDZ4ZoTWliVenHCsG/LAsLHue+7rp+fMWKw9Me17xPi+8zZSB
p9BhfOAb4n4aOSMVrE9AcV50l1n4B90P0PUvbNrgTf6mFa+1SjbbsZLXgAVLQQRXDR7XLB1beUu4
cgoImnSdIGOo622ORpmb6zosL3r4P1NzgH/ZUNa8enOpBIT5dZAkgZ8mw00sp+RdnbYCrg17ehB+
EdZifwbWcCtf5CV5fcG87qbRI7DNnSbSTzNqPNkqIdSfW4ATW8aYyiWrG74zS00/lW1uN2GXhh0r
CqEnIEj1jrU73mqazE8lejFRDPCqHBRS80VL5KY5SW7rY/0LuiNSX1KdJ1nk2h6bnzeHm6T+rHPH
D0B4Z8rIL/Nl2K1B+Td0+818bXe6w4fm5Ct7QfprxOL/sLeF97dhPBcGBlyjQuR3/QbOsEIR3ZgG
W0lcPN5EuHlgTIc8AmeZH6RDIX5CzLA/WILBDO/JEz9jdOREVufsw7MI6oSmujB3GorATt3wrtbo
/86HLCSSBwKHwcGLdngm8+lxb2m+qeBbI4vjpe9O2dAkpWDNva5jda1BnwAjl9M1xK+YQpWb/AgW
ikEdNtnqX5Dxz0M/9vwwJ8JWBpjRtirgBiGlHCKeyuBswenWcKFzM4UGxqz2HpsBSluoHxzVSW86
3Eqw0FuKmLyJezgc/K63S5qaZuuMCRRxXbcLZhXXYLnXuLQ1X701fxpj6zG4O06B0uepEWDhcycg
4L0Nr8JSw7+e5kZPCylYEP7xeOlbsOWmPdsCsGKVoQhfvRHsogFzLnT6Xnbe2DNGQqMlkF8xGQCx
T3Rks0F10xCeXRqxO0Gy8KUQ5z6FQU+742HuykLlBA5tYJI+iNFe/ew5MA1xgYGyMkD3bc01DxYH
vUpTHyQdVYdThM4WFTAljlP88tzzu+x9ikiCVx2BNd23b0xwdDQ0APwI5pfn+UScYE4uMyAlVBwi
bGB6Iy44AfrPzqrOdvoOVkL4rQutJImoS/5ZLOVhMnvsXgGaMVRnLuFvF7V/h5VCoOlVXD+M9Zsi
rEQzNj8Tf+wx5us9/6sH++l61J0QGcHb1Yk1QT83XtlqWD/MVwqcK5mjVzK7Qt/4ivvaYbjskdXZ
QVPAtoYzo4q9VIVAmyayExCjFq0cYxlGQ6vT/GLRxGzLFwlPgwq+XKxp0V9ynv+9J4+tacj9Y3Hy
6xIlLGFAySC8TfyMR2CVrBT8hS6n/5emPSxo7nXcOoCH71+EpzO4RtQTSj8B1UWC3V9fnu2pQqVV
X4HrIZAKl+YQE/sEr1Hm+4bkGMBt6Uz5aGvRyOkPZ/y39JPcwY9U3laN8EOA8E9fgKGnZcXmafY9
DlbB+Rlx7VVKLa9350jJcS0/h1I7i9meFToXHt25DcUt0p879dYcQWGRJcyj1io/3k9v1dP2nLiH
6Qbx1NJGPchEQEBYX6Yu59Gp1jG6/yfGg8tG8+TrJ5l1XDLVYBySiH+v1nUQlxL4GbZE6H/CT1rT
2KMitpf4QcvZBpx54Cx8bBk5ip5/ZN2hunvb18cp7wsG4m8G6nY6g9VU6jCdCg9Ytd92yCFK+t4N
v2CNi3UMf+VM0NHG8Y1ISt7yw6N7XZjMH3J2pLrVZUP+fhM2SL+tBepxG6CpJwxl30/sTzn3/5MG
v+oDmRPcgiDJm/HzzMs+L/xuDWj+nrh/rdLM78OQJxUM6eEKR4CXwT4hyShgfPPkCL8/j+ZOMtpl
2PTiHvWosZu/7+r+NCfi87ViPSopQdWN2lmhofdt/7t/V9//muCwheELEHZ1mxB/CLA9GUIfU2K6
hAWl2eLAdpb8j9vu8uQNpUdmzIFVJrqbv7vIKmHfW99hP7TKYRqLx3WCKyOp0h0hd+VovOQ7zBcb
A4AkqGUMko2wI6CPxbOWG9Z1FIAcccF0QEeaU+kqayqrzy0+ZWRzIXg711Hdfp/uHcCR9FEbPY5a
VcbMnETSoTpGXcIwf5yMyxoZ1l6GBnnVd8kMbowD6rgAP5Qkgpl0IqTk6lvS2t1E8ysbC9y4HHLY
pQfEAiyYY+DLjMTa8AUHp2HY6fPLE+JJZ1R2w5Ps4UOSfOztXO4k7t/4CUvke/0fR6W5iP4rJkdK
P1i5srMCYskPxtz2iSZ0hxVfaiupK8iS5NsKUwFss3CsxXD6YjwqGsLiQtvgszckPLde8gwJKJI4
N/epqkqBPL+AQJ5qL4rA8LXNGExoEifYA6ihit96TwPBKfuCcjVXZ0P/Ps5f/XHkJoooKWfiDTP+
38YduiYVR5oWekWbEoZxwIaXXrTVovCWi8aOQ0SuNan9LCgEhfEZ2TZJpV6lzLKK/sCa7a2A2rpc
SPBGMvZeZoLgMXI3zZPc1XCAWh3T0gin1ETxJRmbSa6mKN6KU8JX25q4zaLq9a5RAbXm7ds7wkEA
KWzei0KoD/8pVK3my8CJOPF4Q2JyEZhI2dPPxyhWibRH8C4neVB+1jnnFvEogJ9LWjTeZlVFFGzU
G2QpBrJpH5FIasOKDQtgKWCLjsgYibd8j2oSC7KqqfkaYX0/bbGGKGqpmxZRH7UMsyzyR/M24Gn7
Xr2KruylfqBvF/vqNsNGF0nLiLo5660j2tWr3zTeOuTn9LSzIgZt+VWK/lpqidpae3cOVGzgrMpb
wBpIAIGKCz+aC3QcK5EOh+KKHPyTCZvOuDHPq96rrixw0czj4Jbc7h/IGWYmIeQRr9MhUDgxhFcT
3FbBe3EroZ5OZxE5z3yF+yjll2G2WKA4jePRxepBxH1zmLy/GgGP8lyONpCYTjg3JloFu7zoDqR7
5aqr4MN91CCvr5pjV5CikwhvT3Zh72+bvAojPoHC2Gpb4trIxd9ST/jcrVTpNbpkOElEffJVtY6M
h52jnY6Dk8wrJnYrzfoEEUx7P8PElZ/LeiPHqZO01brIcid0quKG3qIlcVFMJz28KR2DrX9pEucM
4qTk0qaavK5r3AAOclNKTe/Flef2KvRbiMJtUq2Un2VFlcotRAXFBWPHDbfzjXuopIgkA1vjM69H
lK92VJgjYOMWAMvoj6+OSPSfqJ/WftOxFszPPxUn2B0EVThJ6M7h0DCaURhCtnQsGQBZ+DXGk/hW
w/d5UHU1xSqICr/NaFkT+pO9i61v6fJoLIuYO/yhSmAAvBtD5NGbXdHnp+Li2u3TJjMuhpjBXEfN
XkIU+DC4jcQ4v2RZf3Cu3RJEI0/NIoMBampNx0aFRG5p0CJj/QzsPwcWPUvUM/mR2xPsU9hcWdvd
p3AycOXlLEPGGl9SQ9xBPOEybcn5RmSJcrUvTgQD0sqwnPxQC8kILuf3iGlVlnLw4iiXAk7UMBfV
vCT6L87pXp8dZ+YtED+agy29v8qTLiiQCFg/fsC/6hcB4/jcjSYqS4s9uKvzA714B9rYs8HOfYXy
oEClPTWN++DCh1NTyUMk02PbxwlTbLvV/wyeQA9hobP+osMT0HuMdqgWHnT1y8s7jbJh9xMqjDVg
m5ahf3mlhH+5i6AXXiyDWp0FOS0I+0b1V1RLS3QZcdlGutSOSu9YOFuvjVYezcQExwQP6YCdV0Dp
H7ekCyP3izRB1+bFnNWneTDieQjmbDB+UkWxoy+ktSmBsKAGVf9ma+jYN5g2r6lX6+z6RDC9MJu5
9Ms+rSJ2Gf1CgU35gQkym3xwxGxyuS7RCgYQqVagDBL64GKeasCBElRN2RdRVpvuJw48z+zwgF+r
O21DJ1C9p1uf7kOFb0XZcmyOQ2DokQ4sUztH+cvvYH7sTkTCczozxNn/vHJn0OlyjrM2WinBRiXO
luHG9u0yPIefH5DGBXE7PRXUIbtdD2fv8m1IIW99MAdte8pD9VszIbJdmcxhd0cL3Bs8U8uNsCjt
/iS2eX1to0BEQdX4eBje5q7BGm9KMk3UxPz4qzvnDN6j9cMR7qVzAWZS9YKzG69tuhVy+zcphOzM
n9lUazaWi6rzYgMYjG4Y20skWymPo5rsLIAmGt6cVaqxtMdOwA4JVxiZhSievtiaheTKS3ie68Bo
mETQn44LIEtqrta31uUwGzJh3fCo6LYCV0sp5UVvEu24p8bl0q+15j2Z36TfNBmQwwS9/EYg2YUw
B4ofC/KIU+9Zx82I868MhrPzfzQDYczgZqT6yQX9z0WsRAm08Oi4/hpliDaUDWIAcJdrrWfoOHN7
ZBPRDWMfxQxd4SdVgBpd2Igt/atKc5v1cdT/eOmJ586PvVszcS4RWH18OYRC1IXOMGoQEoJODu7b
88aJQyAD+F7QAU/FnQ+0O38cuF64su2UF2KqCxKjDS5aBsznj+7jrt+yZARasJrCws9n7uHnx889
6eubKwdq2gEL5tpjpG41eImSuH7UdO60CmfhZDp7RLRdxQ6WkMAakPs9n2q27oJH5P1S+G+DYQbk
cJoOmIg/0klnmClGsx0P8TTpzbjIJqbE5bMrgtH3UUu01O64x7ccCVctBlC2bKjzKOCmpCSi0PmY
rNCTPMJCfMe6OjMR3RLzY6iuFbLgIYa3MYoSQ2N7KQ4KDcWQQEoHuEHk4DkvhEhhJDcM578VM+pp
OLzLwKCi+RjFd+FfPrwUY5QImQm2rBaetS5CHTNB2jWyG1HWq3hvIn1LHjIGOQYFQxtjm9xitYEN
urueQIo97EiHQqZwNzzj7q3hzPqQRJD2ak3Nm79lOXZzCKz1gEwSxPpRLUcCoSPkamHFuDrvzCwe
ftfkOM/4I9bg9mZLcP5bq4EvMAq+LT13Pk60VX/pCW5cKQgfoiWX73NH//jeEB6rE4A8rTsSVvM2
PqdR69J3e6w802p1sgpvkg7szCQVYZN88TA6OAiK18BHezb3OVcB5RF4wEY2kDXGaNXSdf45xu8o
40mFE2UkBJFup/X3Kyca59Fw6kH2g7vCdINvGVqIKcYzt/y4UjQywaA8tFBq1b7sgY8tmQa2dsrD
v0sKeFc0Q7JBIQRwoR59dnAlhCz5IqRiCS5TxgCILInI+XgGolUjNFkEUrumW8Js8f/5gUPDGyhG
Ed4za2IliONbUj1dPW9EqTnWOPUCs6sN6a7vQWjlWv4KuDEN+iU4aYwPInbtktqY2ecNWnhIcnnl
eJ4G1ob2YlEf4h5upqqGHiiuyiaWga2ohbNtNcAh2BIP81CGbwfYpPIRRVN4ulgrcwIoxK+DJW+Z
YETKS9ZbF6Ce4eM4cz++ekv5Saph01/Zsq4hcbQ/NzINMSb8wwsyeLHIsCnqrgxqXP5raJrjMvxR
N82PK8BJ2vkBuO77JtRk7caC0k0Dg9+cH5K+y2u+nNLLHPvECQS/VgUOz/znaCvbIxP/EbS+cC1b
RrunNT3891/aTlqTCZGIVvSR/psPya2BuP+swgyiVVd7lJxwgbMvoGUc9gOKPuVPnBd/F3Hzilti
GaV+zTZkpdFwQ0qrvs8SKJhR4q10pp28YN01sddBaF3MTu0hCGaQ0zSNURjNaFBO8PjIvFl7iOSW
G7PRzAEtAXMr40BCEdoWKDy2Cb0ADCDp5jzm9m8zmx9rt+ZFkPCJCKgtsFXEvnWY39gA9aqHUsyw
dx53aFMUnl0Vmpp9ZhXyy5/CkclXSsda9V9GYYK7dwvLlso77280DdAfN5D1J+fPj26tzhy8GP3V
tlgAPPgn2k1VXLJl3SBReq7pqW+6w74x6PuAORs1KuqgTTGxVbvgQrKzYR3a6IGrhbgmY4mTlw18
c7S4svc0WsUe6i8RDxfOjc1YQnbhqRvibo33Gon720rRSUCR5gR2xXxtgdjA88UhgyKteIU53kRQ
5VoEn9uaCcufTBCwzYEh6w4hzsiQG0K/0ePs73k1tmEeT541nPWvnn37LrEMfJyNhw9weujBq/lU
/Id+3LrceqEIfGp7ptDThjF10TDagvKVnIowwttSSeG3AajuF+YGIuvLq/03rCpFZvUxMijm/yFd
0x1dehrTAiHW1Q+TG8uAZARjgEC3UEjB6yKBvDVYayFg8yteAZseK8ASNVY20LYWdnh0IF+IgBAO
QTpms1kf5ZDHlbLlMFehlNiJjZZF02EivH13RrZJo/wJl3hSouYFZq7Aeo2e1Pq2DGVn0ehWVVRO
1smR9ptBBJiVBe2bTujZ4lkBcaYcK3eB28glyS3F5t9/djuDBHSEUURL4ZJ2Hw8IIgeHP9xohj/r
JE7mwwLwq1VDUFH+LqWqY4F7dKvEVJ/Jv4R3zTz6kfVwMdsl5qvQFhxMDshAyKeFuJnVtUjzYjgh
2OLd0vBe1vzFKrrse24WBO4Rg0wd5fAcrqhWEDz/hBChmmliliCiGQq+aw/RniRfiD5hA1TW2Txh
1og77lNugDm57JWuKNqFO4KvNx5t7qvtNjJ0cxGPhWa+tbsORn7lfZS95eTLRFGpG9CwWlEWEPae
kdHWYIHtn0BB6UbEdXiTR7DcY4+5x0jyT19mraKdVMIxp4R0ROWYUlqFKBuxjm6a0hKJXHVEdjVL
JrKyfJWVP8mXuVpiOpGiAgxkrG0zMBjyQTF5mpOSavdVgd0UWt2Kor8Vn1U7D3Sv906K6OaspWC2
BtvT4wpLu8Ww8c3dMdD2lbAl9/0zQwXOmDNYCDOIOZDRbT2sGFVe/PtMXuIKMdjF5TQXvlDWFRQW
aP7fdg3CoYmqPHTy68zbhG/+Uld78riYrdimFjoiLZlPio43ORiS3MyNEDUx8Q86fztIo4nDnCGQ
htAqFlARe+EMWLT/Knur6CcTgjq3By1RK69X6vqZIqKci3TjFITpmHRY86JOPk/ig3EXe5clPDMj
IrfMZm0MLWrGojAZvBp7taSVmN6dG+5291zLcCPjrnGn4MZ1oGZsy4nQaOQkJ7ZNTc9WNo5fwWiR
0hBwdjNPaiwZ/U8YOI3o4MK8xOOOXscNa0Bfc3A3rXzBsTDdqVfpJHWHlmpPtgsBxcruVXwcdeC5
KUsyyfS1KGyoKB/bh3YmFYLBd5CgjPRXXymlrY+BsatelUebzgmWPjef6WFbFjm2DSEdTyMedrVH
Fs0+O17zIbXXQYt20wiJVoLD7S/07/DlokvKr8Tac6bJW9M60JlQRLVPl4iqhcZz+Gmtt2iDk9Q2
Z+CbLzuu4nxETNrE/u6VqGHcUCM+ntlSTK/2siOS5+PaDNruvHzBzM7OQBR/dkSY+OQymC8wDqm5
EEPfsx2RSfdxoDlTXyh4zfj3jPTcl66lzJUjXrX9Wm+Y3F+BynZSJS/Ao0bnrO7K0QpVuEQG2tX7
ob1U1RhmJc38YW9Lg7ZOxYvUZmgynr+8EkL0Qj3VGNcKN5s+OtqW7uIyXfOf5AKz7Ov+u5T45VMi
7k27BTXDMGRueN14myovnw7WxNGAAxN7cKJ5Wu0xWF/RCZvQlxpZVXEbevKV0BgAFC2s+5HQ8DwN
1oOWL4G4XNXDCqkC/cPj06yXyrCXqqg9PiteWtwdxN9HT4t4rG/Vbu4BbBgYvSvGeSkOjfn8zhhl
48km/B0XzMgFLAzhKIPZqEPQ2nh3pWy8EDpC35QPWk67PJ+ZoKlGBpKHapiuGQNRHzyz9RGDGADa
SL1Zja0JKPvbasNvawZF84YBm3iWNsmQz24npxSxmknyn3ltmMh7cFvZ27fg6qt73ZQhL1spXUue
Qpf8vATqmqR+MyWdLIwmbNgUwWwPfqu2KlIyx53Dg0yvxXGwaI7gbakSxQMT1t3ZVh+iphdALm0u
8z/n+Cz2iiHt7PjzstV+kniUmBlTkesZI7ZGK18Ug6w9kXjPcikabSGpYjFl8Vf4LkATRDbG7eqR
ci9I0wutlSjJ1KGHRWYVSrpihTxkKUD9oxDRSFwf0gyMqdgQPc3T+hG1yFzjnRtlFsPA7F+VvxOM
lGJqBjAd+IX9z059icZ+shljR/ZZtPgyb4lthTJTB60US/4E7TthfgelRrhE/zEWR0fJDkWMHRdy
ZR6a52TkK+Wi4254fJTLilBvwD6x4ROwRnNngpojfeLuGumsR9Zzgx4XQ75bKzGnKhqVcE3QOHfw
qSowgpwhwpGBRqpxYkE46qy1b+GkWZQnamohre8uH/aFlaJEVvRojYfoNqTITTIhdAmt+a2U4BoN
fzIKG1nyx3OlDEZk3OTanVgtVzCD9Ik9jd64QM1rwTP5qeQC5ysOjlxG0KZmChqRA4z4UACI/RG3
6hfLeVn+0SW/uTehrV1ncjQ/5NjDolvM70193zrYZNvJzjJ2+snHm7fnMmyEHgEYlkwVnqu66WsQ
ZfQ3TO2xyWL0IWZnJvB9VX+iGkZ9JErwvLSlOyZI34vhNZ4avpr6Km86ekQ5NLOrOA99EzNcdI6W
jD0p1TtEnjKVxHFqeA6+rokRIB3v6EFPzZ0C4++chrXWqAJHQa2sA6gAXKb6Y2uAjeqAJR4vG1Sj
E/Jq/h4ROtv7UgfqIfRodCVa/QxyogplH/slG2iOWJ62bTA7JyqGjCiwAncs9719UHrNI0yExvdu
OA77WDXYy+BXo1ojHp9VjbhjPX/Iwiv81/GI2ilnBS1ADLuep4Rerwx0DPxWjoqs52LRA5oR2GdU
48d28RZ81ryuTw8tAqQuM6RanSRZFbo7Rs8H2dPrv3hdiyjm+/u3C/YOATD0TlLvc16fp2Ijh6si
zU9prpOb31GkFNzhJGyyhIsZ+z4CSm4as/T/Kc4xQKT5lLjlm4MmpLvzEStY8SoJhlWvVB6pcwL5
5JzFJ1Nce7688RtuK2O7wYyimSbmBmDr/7YdoSM97JNZ0IptV4yj53cSIDo/inuUmxPdU+VyTwv5
dDBHSmCSjTsnZFarmj73FKKr2AGguxdnnWU00o9qtIWt+wXQF09ws0XKrB+MNl9HIVoYZs+8DHXl
wczxun1WsynXldITqCjcl0f+o6YdQPV0yLsb/aHSGHhfVl3F5RbO6McFU4JsuGghfQYHezIcfyrx
czR/CBIGOIoPUj8W7BywnrFz2Cvg0XofKATGA495jR4fQ059HDNzjzS9ke25T2OtQahXbRdpQGDg
bSg9eGnsJi/avzNg7PNQwvy9DJ277EyjaO5YNunp5+ZTHcmqE0B3tICj1d40fhGckkEX4LC7tBO5
gW8qO94q1Q0psDjiCbWPah4peK105eQlJLSYqrZTh2HKGP0dQkZAopxexr7I8gxL0Rs2WRg7omUX
R3yRnpiwxKUs3qihzqAGo0FYGeCfRbyttkUcl6ejmWRdulbpLtmHiMXTHosa47FVkvLX1tK+xWkH
EPHh1lF/u36p8ZwMUNThiDBIHQhGyVtn1INyJLZMyBZftC7H0CvdCsKMA8bqLXwjZRBvJcqhHJMk
ZAiTe9yrvQu8ppuQ9r3vL3jPfteaEWKn4Fn2pv/E8QONela9A7ZOLr/6wHG4+NNKvVXrj+21kK9L
1ownLbSYpCURVaDFM1BLQ6O2Cd9KHccbo8LOhzIqpGN7gv4KQTQK9A2w5akAIi5SHzM4nYcYbYcd
D3wasyGj32lF+glIbSjgdmY+aqHv9yBXPdN751I6uygqly63y87YlKgjuQrH4s1Elc+2Ncb3BGr/
o4GEQ+Tnh9WYnrL6MHnYZXNDB4xDDou8kYdGZ+idOxkq0SfEtiOlf1QRmXQpmRxNJxAC/fNPpDH5
fM7lla5Im7Ldzy7uZvm6AYBio09FQqq/FgbS8e/LV+PrN2WU5iizyf7/BvaD8EZCG3kkaQ5WbVhZ
dMnhDUnI5MZhDR6dS7sZsZ/anvN5pUHr1YxU2VEmuBnUKm5kDodsxfPBJ6j5bSGKeisl0vmiM/cz
ik/P8QotwRhUsLDahKsKvGFOA3iTHAqg4NzzRD1ttUWPTIapurgR5jy7UOzH5ZEAOjS7iIHuIHRv
dCOtyUrPka6X5jUstZv04zrp4q3KWa/gAEegtdBJuxHIU93R5VfAx3gJfDubuv6V3kQ/+MFZHyEO
gj8AV5t3ARuaDcyb2k1eOjiXte0dFzrDL6+y/sz+RoA9+7HDPn0wATlB30dE7tig3mHRU/BYVPr6
Yh2qDjOMyhh4sEGYmMsfLS4+VNTsFLnTElMRPLzgDHUC9TkoLoRD976kL3/mkfViLoOAqSoZNDvt
J2iuGeheVGx4wAxWHDiNd7jTh1x5g7OWOq+OwmNgItDepL/8rUE1NVQ74KOq8TbdYaoOF9vwZWFp
haryEQKWxnzKDvOa8PvxWdTIT5/ltrXXiC0jto7m/JmdLt6UcbCJlrj3e/GHzeJzBvUCzQl5dc9G
1eHGArTp0vwLi4ZpF/FbF0trl4m6lXki+FmApxomsLm8rSVKL3tgKr/u6jhvb8KJRnwQLgiPomSR
IsOzlO59CNup9V1Mt6sD1sxZO9Bjp7kRIlJUHbmr4GSTlMwxKI1trQcv8idS1GmbufwxDpEfqifO
SgmCK8zG7y8eqfBSwoGNgD/zqVccouvkrullqa5oepbjmOxSnjPLTmyBZB9dx1nGU8UJwzG8IZ8k
FSntQAG67pLtrMl1W/gbHlu3JL+O3K+LALckvQfc0zPxnfZD8TZbmvIdb93jlbA+uRpMHCFi2TR0
EZooA3/22B+ReJZWEWgYfMV8qYD04lONiICiqsesW6rwPu4daXqLCMb1rrOlPsfVqj1Kgw5XlhVO
bdasuY2+cRIk98rtzvz4t2R0vTvPpg/rrGvywkzOadLr7/bQFyxGPrbyT9fqDj21U0CjG53YFhml
Le61xLy+wp4iOMT0KqGtqz6SNyhJVo+u4VZ70PtsB1fbun35w+qdV8vFxx+5rxtB2NPqdIL8ka1z
IEeREpkSSic6FXiUMVDweNKy8g+382VPoOKfTL79PsWOCfYjeEDkBJFLHv3/uE48Ql55iMVH761i
GNaZQ+WhK3BIoTCpzLIb2U6Ee9ANe0f2LVQZbqFim5EJfhkla+g09HWVOdQ6HXxvI/Uq31sCudWI
Fq95yeSr/C4QyGxrwvKt+D06rN3ca+oN16q207fybDEUrFMSPMbVad52687AE0QCCb6F4kle2fWx
b2pgBO3karcxgQIpb+CVn0qCDd8FBSr/VlfsqllYLjKW78j8G5wSuyZ8cdRvN0zxUlJg3PIPBbGI
uBhHhadQNQlHMmQu5sgWdIlnEFJr4d577iMsr/aXFp0P8SGmgl3inP7fQlQa7O/dz+hip6MUcMku
oqjSpU+3w4pEqI7p6cNXJGFmeE+TVTVPhA0Wn72+sDJVguAiHYUf/aNo3op54Oucfce3hbWFHVOz
LNppC8/VvzVX5I2DEekzk+dhx3JjDA8Jsj4XJvU7lk5C5aO+nLARZH0OCY2B71PE8D4ZdESAh3jL
SwocnkCn0/4wzLpCtBtyRTbcV1Ftv5IM/gY1BqrFhPu8DjDGL2ZhTUsxn+sTUUsvXw2BYGfMGE1j
5Bnu/LtFFkoqz8ToA7RJMVk8s54GvudsdsKmFpVGAgZ1FrOKKJTm+Co4t01q7yGF46MLeseqD8En
TaaDkrGFZ8mDL4A8v81n8vhECu0lopzIL3pJxqUDsLC6S749xTAjN2xe1O9eUhsbWmjC7FXq+FsC
0Cu95Q+iR+wT1yKFmsB1D06tgn7TqDt0VyjxNQ0yQbkEpGTySob8esVIXMEsmNcGX8TbwCdsOUPp
eymMI4pCzbrAdZ4zpskjnBjDvbG5wOxU3EEEwoeJpEYOP8zqXprOCcUaSurRlLdkkOLeiD9oYJm6
62fSnwgp5Nz76UA5G9yOb46bkufvqfqIemBFvKQBqCnLUPXGjwWGOCU8JiocIBDP6/WlypOQ+iQZ
Fd6Bj1rzdsyYMvEnBbcaUJ9ApTCF9KvsUtW+QS4g4cQQYkVTGaMWsORrh3iygX+3Em5YgpEfWkha
bAMvQm+UrUYu6YPx5qNrAjgFoUIGq3xPd7VA9fRvKUdLLmAviZaSXgWR+iKF6DdZ3Q1ZE5xhRJY+
ZhsY4USW5VIyTi3MpfCUKIT4JSU3KMYKw/C0kTtf7fmEiEFvHn3VYFetOkWlmT7eoHIaLfo/zKk2
tAq8//jhW30ytaG/vR1x+fNESG028KdvIYB8+9jTpCd19W4zIC6KjQHcOc4g9greeyF5O9aM0/gs
DgUj7PynBXPgewOAoRB5BNu/t6iXEW7E+zILq/YmJFeb5Qu95Ti+ey6+qib696tKIZHCUATZQsZI
XXyDgUhc4wyAvuGNrKMVQLdTiNLqjYRDkF1ru5+oIgLwy+MbTX2CRohj2y5pEIoIsWMx8ewcPqcW
NnthcavBVCC0komYgxt6xlO0VA8KLZnyIYZz+ZVbm09pnghFs4CZIIGlFEI8Pu4eYIroCoKMEfuS
T9LAMOq6yeNpnClibCZdKrouSlWfkLOm4T160s6nDtCpttp+xD4ix2AvlaXnPVRCrRmq9M+EOco2
jKsmYP0NCJ90vlYdxdg2gZztC517CHIr8z7XPPPhch+8Sgi4/Dw24XPRgFDI2+m6Hjxbc8EgTiGU
6lAbmuPw31GCVLuXRVjXVNyn8BJdJsOrkcXUKK+r3I2Ws6zcfBwkUibxCvoY1/iYcwW3wtJBtr8B
lJjd10m1lh9zyuIPUIdwyIbrZYNz0GMM+ozJKy9qcQ/JczUAUzmliFKzuy16eT0WwBgOWo6iwMtv
QUpqfXRUtRZtd+Y65EUbz/6/2+y4bT/IZbi7qzZefwUJcNOk2XPVBEs8Kw7O5c5cjVr8JoLwL11h
n4vEwP84UK45MH2RyistdEbrChYzlMJ81JS8eDwuhEF0b2KTSaoX/K6qnZKbHQTQttarq+X5qW6s
IBvX7kZHxdkuijmSZ24LBWMO/tiiQ1XXN1IngONaasDE4sjlYxV0rJTgzKgrteB2hkscJmoqK7QW
RFlYvHyxsvSe8zG38+5Hqbszua0VhNrNZxBQwvk2HRj8U1Ncbq6z+hboEKyQhXAcp9QVPFwWY1LT
DvDUQ8Cngq/V7c3geBzq5VKIssTWjGl5LIyzRz/3ZUeAbHBUdz304ziDJ3qFXv47XEzKrKOQsSty
Hd3Jms968REgquEcW7VKcBIJlZFD3pALYA7VQ5nL4gL9Shh7KpEQd1pb4xvFzG9JRYKUMss3PvXg
1t/xZ2+Z6GRJIgzsQsm+CNSwfMq83k2GT8CQz9DR/3bILyG/EdWNjNyjVF3xTcPKuZ96l8qB2x7S
6kh1BeyvN7+HBnPVX3O5tdZ/Fu+AMm6q5oygrrkV4655AwnOuFmJXx4i1gr1IqsDEsECYLwzfJ7C
r1mjNa5mawC9+OltJciO1K/YxdqfSVOh9wqtz5YyM/XQPwpJ7wNBjd7hktqN8JfooDnoVErGldQV
Zcz0dzTjYPWgcvk62w+XVgYwKDwsXaowK3qtw17k7v714CC/rr4eJn2cFW0Ja7L4EhvCQdAj009j
qLF4VdpvRNH3UtGycgDG6kGPLuWzCoOFQgoTn2F1u7t/GZuN1NCX7haC5gvW7YwAR3n0hD0/Ee4E
XCDi0ywJ8QQj06vXqWJy5aWrEtiHdUwXebg9d3EotV/lifr8S9uEix70FsGWXUOCJDwHlynU5M++
cklGaUNZ5lAxvZJKuCHc7cJE94mH05/WhUbUKh3BuY9x3pDNTIFNl/+lSgkSJyliUns1IdxoNCjQ
RaHc4nJjXTbDg61BGNz6sdByFCka25ui876p8T1212czo2WsybB8JyU8cXxKTIjcTncqUV2LBH/9
wcApxScr2vrWx1odTXKJ0AAMCDOE48ege0THl0pSaWYhJK2LvAs3h1VtCbhwL1DVr2RpGpot1phU
e7Z15UV9col0+kdPo16ofqEDBCcQxDnesa+95uozVWjMfrp9soQrxg611F9+t908C+LYbEijHUU+
x1G8C1AKp+dHI5iJwBwl0F59uoGFaFD59HSgK6T2CzpP9CUnuZjEfCgs+p2PuCulc77jsGdb5DU5
jOv5pR/GAUqenU9YEhrL7S8rKpIXXcBXX5wXYdyZVEVOYSAzFZGV0T3llDdDYX+JADIoroCK68Mg
qDFyuFikxGh0eOuvBB1+UjWF+nndz21vSKUHo6Dippd56X9Q+rrDkfW9T7xlj59GOxkC+0FKoH/0
g0NtYd3xcTQYNsqzoHnEX0k6bU5Si3fvDDPK/UYzLfizCrLIuDdZ7TTwgp9oL1tHVedBIUMdi06B
gLAvrytGpQY05UQhmlA2jQWrSHZFQAz6ZtrqOgtJCQTSaJga1mQ5BOB7vFGlTPIzEN3MqF32ncn0
oFHXIPwlERuGljjFrApi5f6Ekzcr677cE6kJkeI63tsDCEqhgEJTTGqyeSi3sBs4TOaDGlIB7HBu
EuAgnBdXImHzu3daj3GN9AmR3D/0skxfO6g+C9lt9GRl8G+rIqZBWSAMOVB+RD8FF65MearQL4/Z
zmWsM8NTl+iRBU+5Vng5CLshqeag0iFDnqfPsHE6lMTuu6yYd7mOMOOwFMhTJ5fUQS1/3nPK4rCi
Fk11pBLKN7bZRUxoD5CGt4eItb64isBPEsaOvPiy2sGx+UXaLTwX0cHYNCIefa0hhn8yGQKhDm/A
xczT0kIH+aXpdaUtaZHhXrBo0Hc3qHbvKQhtK7pd41KvDLPoYbn4rfEAQKMmL+jwp4Ut5DMsxoNu
kc6p07QUMIUpd9YZiH4O7xfOJ+bjcWtUTyBL0aKIF65/8Gy0B9GfODlF0rbp+HctlWgMPAyJQqv0
9eDO0deQVq7l7Gen10JcpOly1UweBTFhQIBqR9yoWc5ndvlJ8yXJM0wVnXKlHqYX0zcOeF2hY9KU
wg7JDgzk5K/ilyUZ2bmi9QqVpzX3gSB9C5Uf8F/pw6SpGDJEe00eCtkrRpm4THLUyh0alTOZ24Fv
R6SOddvhZAuTv4XiUEW26WKegE63mu3YnAcjAYkoMxZI3GmKLd8n+zs/8BBh2hspIv3fyyKmrbMi
MwIBrGR8SwoKlbP0TDWUKZcUsfYNkTpYqs1DvNj4NHNua2jhpBk8tpDONBH0cQXfVrTPKw5UoMnw
HhI0IwJ9biTxopHWCMq3BuB2i1aNXH6KycTZ4XmkvPXteO1eVQrsWLHcAkqKxLGgCs9c6CgOMAvt
cR8A554kfY5+MFvGwCIfym8q6lT3/igbZ3iqz0zImaFcznxc0F+jAVHSLTlMZsz3h7XwZFZ5qleS
XhA5Fu3QD5YUm1pPknkXo+eSqCyOGPRGWFP9yvJbs0z++PhAN+ry8CARcrULRRIxwt2mRfjPB7iH
vFKGRExIL8iLo7VeHH0nwsIYfNxCsvO+8fhYxjZzqlqWjRUiId6zOyDbc1dsa7qC6gFRhRhuH3S3
C+61tXRCuGt9T0PM4Y3dEQxY+wuAS5mrLcYBDP7kKIcHqQAHVyGmf0BW56EbzqusQrcHakHL42WS
90vPrTT/+hu4qckWFY1I/zcw0wunkRc9WfTObOjM5Lk3zs1tDJ7OZ3k500VI2Qq7QumPg7GC0Udm
qWIAEdfFe8WKa33gR4z8Q1NeudLIcyqHJl4ICVZR8S2AD5RY1Y7mAk9Q3UCv7qzXgfFdorN0ymNV
GWoCglqE1HDGnUuXcQZvydERu+4H8myPXFSnoJRHQGbQ1T810J5SARCnOCuRyyh9uKyJxmOxw5ye
C3mfOHgtMhgfXFBDJ0J/DjXrHV9DqsGf3IdyXKCuE9tpy1kixOGXFQUt8vNATjDXSfxcjm1KZsPT
I85KBRsCH8l99HcTzazq7uRtDGY85bQpeaEI8Uvv8x/wR3YvbOT3boAYjj4V3XkH+16JGr+JGjpv
2S6angyOV2tD2QSVCOA0cOeHlM5XtVoR8IYHhYbp+DmVq0N8BT5GMGORONUR07zWy5uQ37WLQdDg
xDDzpPYGHYW2WAWXHll2NRtnoHstINJP+/cxtHTMuajbrZY/IKeXEaEcYU6fkDTD5uvI0Gt8Ug+X
qTdY8BYLj7deuZgzJCArIJo0s1HT21lNAUQTGtUk2SW3EaJk5F7rwYBBbCCJpebeT0qKusC8QyHA
aQjmUb/yEMY1SvX9/+YG6VCg5jnOQC7lBdsgL48xD81dOyzxPNkEXJ25+Gd+BHdA4eD/L9Fr98Ik
uhcHTHdy1tWCqQ01AdkGaKDM9x8PAMViWxllNNIuXyR6EzoIhWz5MrgXvP5Y2RtyK9DlfRPlbme8
wz12FGweFH8lXbGvHm/jfF/O3flqxqjlpC/ExY90SM1zaaxMg7sgbPFA7AdiMUfsSerPglaid2DS
LdM/CSHvPBX9ZidFDyhop0vfrQRYXQxGeN77nGCERysl6ZJQHzC0YURuL/dsoxotrkbOI8quZYiA
QPOo8+Paqlv/IjKwLuQWGBO4puYJbyYW0X+fl8973FTUQp4yCdJP95Km8koZa/MiZg9P5vBuHa0n
Ekyms7ABCBhchltbuhSJRflsNJ9SPhUYKZle2dtOp8YjdctXQhnfkLTPGVYF1b/9xdTqPe+Aaf1o
QeeEl4VVT+7mYLdzvMnbqJi84Mn9d3JEQlkKMvS26J4F4trC9RI6blwMhcKmcK/T1W/J7AV+V9J/
83qum4E9GvOmM8AIS8gzAFDbLW6tGjlZ/mmqQGAHe8UncIdQPAz96lfABYjRUvTW0Zgai/Evll5E
VpLAd81x/8R68fhLih6GUZASSVADrtSAZqzsHEvhkOA24/m7U2FsX374D4TmqpvuCH8gd/24yKC2
OJp2tpN9mjNAnWRAtr5yCvr33Yh0dhI4efJcB7IsTypqiVayrORIMleSjkWJ8wIBnvUCS5f8gkHv
1N2oH1Ha+TbB3UNC5lKZl1GuSVgM0ryN9EmNlVkNGxH2hnvgVA9MKxJnNU6olD+WXyFwEvIef9N1
ykqpm+KrXCv7mJDBZnM/WIaAy1KnEDaJ5YjSSCjRI+z5OSlkyF2ggwWhoVAwEEIIJ+xrNF39mwsB
vPn34molw6mUjB4LskS2x2TNJBED6/+6+uqP4AHd91Hv8sCTX+fPcaRQVBy0LToQF521YUHpZnH0
5Gahxks6xBdceX9LftLfTy3NGGaCG4pIVysE2tUToOe+9+uwdJUzTUgdoknpfgLFZ2QVjD4YHnpq
gs5bD+eedcz+Fy4vD8h4zKDsOn8CgIHbjX6P71r7bGPU+sbjsfVsIwVkahXsGTzRTxvAz4Uy8KrG
LI/Hil46aqqb90XCwwt22l0rZMOZV8ZuTQSyhXG2Ln+22YrWyb7OtEVgqXCf5/ArJh4Z9S5sDM2s
6CzCwQT9Du2+DW2eQqof6RG+Emp/+aVDQecVLDls/3F31JapxwZSlSrK37disCcosn5jN+IoaEYr
GgjInjIXO2eSKOscUQ5dmmK1CFW+7kh935vAv/pU503cAsGtUDKL4M/dr7Asaelh7hU44GiwQSAU
dmSZFgSPsMWzBQaFGXH8obW5FwkZE3e2AAbWMJUWB0Wd1CBcu7eptay9H8NxKfjSmkdpPBMyKjv+
UbfNQsyYZ8fHra4k4rco/Fum3SRdYR0euFstvH+1yDzoXBfOuZsMJWnVCwBb0sXZL0q20XNTxcXf
uQvBdvV6WbNCwISpdVUkGYZBMVETHiUmbQ8+QDHQYfCIvqJBccxrCyPnGOIyCazKHBeyOFXah5zM
tHtioe1V6K+ul54/7H+NJgm/c+lZ2YLuvUQ2qa4NLgOUmTtcN5a+GjPyl8X+yS+YgSZnj/geY2aw
dSN41UufU+nvpUyk3RPt2nHDi5yd9SyoUZBKmSgR2kyKb9zZws1Y9kel1BFZiS9CbxgitqsjGy50
G/wpOwUKoOWU1Ub6QS6IfY+iCDNmYcD7KW6S8suTjibIkUsuM0qS2htAbWt/YGnOAmuvpQzpl9Ss
e1m+ktfY5Q0RfBN2HfCAb3v12DnzBjWsfPHe3tEAbFAb/xPAzuA5TqEe4D4X6ZAw9EpLFW0TWJ4Z
yQkQvV4jjlFbdM8vaf98BbKqh/Yn1nmS7w+0aRFp6YF09SkFBL4iGDRIcfmukbhTvJP3kmSB2wwQ
jC1LVLgwYP96xUh48UFdiKY/VyE7eHgug8xuMH64GE4XMELblRine0F+16BuYF1DicVMN0j/tani
Mjd0bKfBo/YKcBMpyKM6Ecs8u16hLpmm1/H5LeNigGuJ3MjiJBYKCb9+7sZAZ8tOSY9FzPESl1ws
F6vm3ziOr+2fhKQCgDHH4+1ZROF9QonLcCoX6Be/6zXfYhcD7N5j1oCZ1q2j5RqJOPa43mA6yVKE
yWAqneC5SkJ1UumjS02N165+T2wMfjuEVKvtU+1vuy+uIWJId5Qe+fe1uzK3QKLIhL+7+IcK/M5x
245M5wTywcs+lhTDiLvkSBpopodvWc0mGgecglVD9cIr7fu/edcNmfBhGYhdUdZEHljZfJ3WonOH
NsxI/K5DQuo2ZRs1LEVygR44Oo3TIoR0zlVgDPioajgLsulHKuG7NwfEFZyJ4hgj91X1p7Stwvy1
57yIZrKZKizOz2qpVhHn3j8Pt6t8zIJFdKfSVrKlpsxTi0JHH8XM2bL4IxCMiWfW5jgOnPrZE1yE
DwZyWd5XD0nH5JPzQVVFuyEDSraoMk7Jh3X6It770w2l6Pa2TH9rpI06JDeppWQtfEIsRsz/40Nv
iR14IoREhPnOlAuyxYbE99vvviQErEQh14NM+eqxz6FGILx9Ewhhhx9jLHtjtqcX4wrzm63MGY4S
qZ8OieYIAtUMHauxYBE4w9N6C6lyLs8C6AitEbxGJqoct9YRLZrZE+A8uQX1IytdCd/W3xZfFKfB
vSL2fIPDCa2OuTTiL1iV/fxFZENiVXPXgwLvXLoy8URqtew4tpE61iKN2/8fRk4Xl5FLjunVTeLI
QkOsj2KUpY+f4PvJasyduLbjSWPYMRAh5mjILEZoUpnbQrlNZeSFW4EdIIGFrDZAgP5/k+tnxMLs
BfxABpqm/GA7iUxbdyJ8nUkWm6Nh3UyX2PwK1bQ9KyjwGErnTFoi+0A5LSQibQKG1vZqmF9DUgoj
y1wruplMTOhRW1+NKblw4zcizJG+z02ES7/89coSDmnD7/Ca5i1S+p0ETdOOIJxlEskQ6oY+To3l
Ys+oF0hPVDm+GB8EXGKH2scTnMkudCkBCfLnx7HNooEvYTqXBe03ZjhbcbMonTd2/XlKXy+h8G29
bfAFdidfbLkVbkG1EDexFIHTUuABa6+CO6H4eRFVTPvFDQpzAahVRkPIPlr3lgPgDTa7M/pHL0An
nVj+SF7zSvE0qhe2ECFaF3XPtpbQHsnJL2D3B/wJ6FbVAC0oBXNC0MY2lUoQILIhbshg/tI1+x22
0K1m5DxQbc5C+KaR2K8QPhw0Qcx6gdTMVKd+we2Ce373ez/8uIASI+5oHQuqwObQFD8Xuqr1WY1o
qCtdg9/HgtsLnvnL1YnB6W7NJWyM6xulU/xKgjbgWgAxEqRqTxViWeh7+auo8GY6kUB0FHyFNnv8
6veLC/ubiUXn7H9ZUWDbdr7eEquCMJiMv9SshcEcGSOYk77nzOSR7Dk/tK6HkT5V2VB7x0oU+tzN
zAi/qpptbQaL6DpVhPMis7+XQ80EnQOPbHrMuCjhTKTsAIRqeVmQYyw060YPIgdsTg/VDXGVwuBd
D31TToWmKF4/iXNcNhedz0rGErCU+WzQZvS0phvo+HG6vGUob6E6YGwssfskexJ9XvYTfF8i2RA/
UD1nxIisMh5m+Z6rYuI4WVZRzVtE+BaP7SHthj0aBnoqVfMDRLGQhzRx5IWSKFpW+cjEGbCzUj7O
zniHjgapU6WY5xggfjKikzSZ8+r+5NvcpO+6BtaiG9meSH4CXzVepJWv9zN5mkt8t/an/0L85nbz
/X7zbgUkWV61nibsa7U4vawIh+N3RWZRKSAxP1YJ6aSiV6TI180ZxkLFcOSHzx857bX4xbgUi/iR
vfw4s/xebzu7WrViHnatzFH2Z4bAcJaZItBqIdKmGBuz5xQRlvx6vDDLMM4D1MIKylgctD4W+4yv
NA7UcQsm5HcOoG5J8qHA6FX72jr+HvfEtqfZOiV2rBOXNhfpiBg2HyUXqk84CIANVWdDqvkFyU1I
B1laDIeBB7P0HRVX2zgPqYQfY5vBZxXT7fX5t41VGjaW93nGiVPT6MSo0DDApbrYih+a+oMIm7Zc
gTrSdIi2lW9bp6YJZPTY1Pd/MQAxwKA7+cMrGYkuw5EfAqkzXHK7puROlTsJZVxuQYQOeKLpXAqO
1xPzYv5ZhR5+Raf5+ESDaKwz1Q9DcSgauLxGF+OxbViWHJe8S0Ga3DonfI7B1oXBqAr4Gd6Mwn7T
4mjZ+Ozzuya0kB6zc54mkc3w7YIEpReolNKYMCoWPqMgkkIS67iXnAVX2Nrv3otnPwwlFGxW6LwN
Rt4v5I6BMd+7Rw8MFXJX8ypLe8MHYVUbvdTdThP10stwuhH3OJiJZrWVbXm6MkGFHvcIMVmcd6O+
NwHv+B6S7j0W5X/z7aj8+2PNSwhP6/8PQKcWIFvBsoKdD3Ant24FTqbCPj5oS7oPSCMwrmF/VtAd
iXIHRsqI2H2c+9W98wr5aw4lfz0mjHxsD1l/g028UvEqNNSHfU0ESg3doi/KJrFvfIfN2GR8jMSD
GV+VaM7I1er+A/6cXS+fUWrJVx+hJIt+LN/+oHfKavi9VeoXNsOP8uj07Ey7WViMT8pHjQHkhynK
TzCNhEKq4qI/sSCunBbH3yep15OpXGTRA+aR1Blt7zmBQXPSiI4Mix0ItNsvMDkOP9WCRWQ06eht
4pMa0rgknfnooR2Ae363QxUj2VwxWnpH0MIXAmcZuqv30L73TymAWPmDpNUWDcqkYIIypu9BsXmT
bNNkXqKc9lMzvR8wWBb+NMw6hFriMzT7t4QGWX9Ta58+TruA81VmUCC81QfSwFFQa3nIGQMOJM0L
Ij6CJUxP5ci7PzHgk33UZsumhbrKFlWdpaAr+KILhdsbufrz/+VxGAK4OkI6/oM67nRZ9HgQWyGM
wcX5oE09czBVxECyBE69dgu44/dNE8x4JWmznna9cyziJpHCJkUN7A6/xeGVC+wsWt+/J49yZXEW
Aav0P+Hj7jBiNwqkJLgvqVbA20+fucn5nLWUoCog4cybhnl5PggFfIiWcNzN3rbMa7219Ce+echS
SUbJU3pPoVTQYNEuaoz89kxhL3F9/vvLrW4pihKSRUkuINEZrJRBDbZmzIbURUNUUFbTzd9gi0/R
geKcpdM70U+4vAW2N0tq3nfpWDGzEJVlzCgN3xYgkRvgrssKKWFKl8t1wDz9Wtl3kxtVpJDsCY8j
sI4BuSioSDlsm8myo49fhHxeTS/xKAlnpOrw+REgHUzYe3IpLJkBmGzNL5AfDtV5l72sPUvdTstx
6Va6F1M6xmqo35VVaUrZLsaoOLFwMZlRoUNvy+il8m2EpRwfUWmXeN/q0lgVzIO8Mn47wIDGGSCd
fuIrZEds9XwZsewnHJXZGeodUQr8UH5ae3w7cji0lTXSyEyMHHK8qjm325UOea2U9or1c+vcNft7
52lLNyUs8qWCU4RSq9skCRxgoxEvWD3UA6UKCzb04qxjQ4lydUo2xdaO8Oxwk/fE8aOsQG38I/Hl
f687oVagy63U2iOmC91pCRBsvVZC6lXfE8BXN+R6GjJkDkWspRJhyJQJiBtOpZzbeZ92UXRMBG7V
dksyEcl3Xn71eneTpvFNN6aXfUHdh0D12BzAW+6/LgmdayHKMnnEWV0quz6d3XJpCJcsQiQsi7x7
xWVsePm95v0wyd5wcLvPk6Sf/6xFBcJdT9SvENOyxAquydzZiO4uv5qxaphFJpdUZGgVBOgTjHFJ
x5ljJmWgEDP9zF/DsdfcIB2cENxPmub91QeI8ql/n08eYB+bdcrLy49xA477+7ig23H9IMWfP3wn
tgc15b+KzoBBM/JL27SbuFUCnckS1h0yWm7xqlSJUfTtOuWh825YQqL8mlmZAR2mP3Mc5sNzZ+Mm
hem9nb/QJZu8xbxDTo6IMx9fKeVqLKP3fZRoKwIc+XBYvC5UeIzEuqtkXR+KhxFjFsUzBp/eI9ro
p4r+hjIYCkMPbH9EHAD+GvDyXVHKeIFKbwZAWtHWJhtK1bBuVPMhNdUYvI0+wWa382oi3yIskKS9
44qM4parz9HAtmRBTIyAcaV9Y/nPFfjrdPe/c5pmGM1pIPmpCTXE8X7Tvj2e4C+yWfN0h4j7Zt0T
HaFid7Jim7c4yoem7xNPJ/LTXhKUx2Q17wIQCRglXS5r7vCsXiXRzb26uUdo4XJ1LyReACXfNpZi
KRq60+vlW8YEXk/U/2kjNQqcabCo5f0VB9luLBpBxjOMEuEOX8MkkYG47mO4ejaN32SnGFuupRyZ
1qKqv9v72NkZjtgOo+4rrSxClTG3dJEAZIxQBCGG/0frh5cNu2YU+KfddpIDOilGvNgZqu2DOvJ6
q5oy6eldwM+3VQuHAv7zGVC7XzcvunwQz3YVqImfqfp/NeZG42NCtQWJ0WLqUB0vSPJSi32VDp9A
vE6ejk1PTxkhUdFeIBE96FkFv7jN/yvF+ec8Noe73p8zLIrhlUrTRHLIyacJQq/R2Eli81C0+Fgm
431N+Kyy6ZmcKlUG4dWtoBj83PrjCvZi9q56tYoF5B7N6ss/0zaN9y0lCJ/aDe2c+6TVk3FpsQdR
FgbA6t+jQdI08y43ObpeGkBVSglgoG4pfNXQhV4d1BCmEzs+762XrDdfhC4tTlw9v/sISdipxzm3
o3/hI2eJVVBr9dfgumxG+iYyHS+rZOulxrC7vkpfuSnkb9TuEiYHGejyuBbAOS00Njhzy3J3ENR8
KENVccDHYRXi6bq3bLOZprSeDogceRA7ExYYS0EzHhdNVXBDJ+nB8r4O9+9+invPTFDDyhq91V93
/cpOXy2BQOcl2ahi2t18exlPTkXAqY+pxi3GbOd5aWTMCz0izp07ucFPVI4H3hNwncR7tVOHOvcV
pbLZtdVzI7n3+dulE07vb3wa8ePzvUtkIowW09cpgAWDebrcx371ReaOuOlhklYiZTwTWLknc6Wi
5kMytp02363NLeWfkFGrNuR912Kpj0k3/emcyFH6m/5rplVRFeM8jV3qpDXwlyjw5I0t2gqG78c+
9EszUtyGitDsgvzDIaxqlCpjWTvg3q4TlYyEp7t7diXK8aa2XZOa0lLBgrOndTvv8yzwYfPpPcyi
pJJw4ybtYmfa+5XjAO7V+5F1kS1u4cmYWxlkAo8EANO47UUx0Fz0onL+GCCHyj5RcJhhpAo1OWqO
7vHMwqDrabRn87qsawnDld2hGXEQFCJs9aBm5UOGn+8De8LYlXPqPVqPPKPeBR/tbBPZwWjq9aGA
4hA2JUFN7ApnrtD5XKH3ZuzXUge3MJsvaqiQOdazFndQ5VTM0jIvmGADSns1iF7ZZUq/DIrBrFQa
Bv2GwvYkJscHnBBYYOiTp9+PXuuXWnQVX/3YFEtbBu3wI0+SfwV1GojEUb9yhpS3lpysgpjZPkPh
QGOvCg2ZL12ZJNGeCIg/LdB+PAXL+zdgSdLB3jJL1LhhVHLNGhofE+kIdHo+0Y1Pf0eoX6xoESBo
P+MbcaG1XpWAQW2dHvwK9i6zJqNZEKR8EM9n3tNDD+4uLftNa81/FlmkYZWuIqjYZ5nnVkQ1iDEo
+QhJn2n6tQ0wST147xGpLRzff/y34wir8OT532w2GApsOt+IGJKEfqaKEY9eJzDPavzuhltgLWF2
ZKQ7QCBSx6jpPEtVHFtpZlqGwk4sqGg7uS4+/gDAeImnMlMDX8egRSv+/mSBkXFcoMonsd2GOiFq
etSuLT7sPfTVOgbSRqUKg3IuyBuG560tYjL94AGyBZohE/8RcKJfC+CYxr4nPza7hqcDd9+YHpqu
av1vR7Dm3Olubh2tqG4oUOnvrPD/axLDHuvViAGo9eYVXg/SxtyKs3ZnHOyPmSKhRN49pzSS39kX
/ewA9DuyeWvO4EsdoF6SikHE/lPBbs5kFbMvhFZa8+k1GRtETnpvbDOEl9x7CSbAkzReOpvxu/u5
WNo53bzfBhBvLKNF6Kk7w0/Llro4NXOuc20eKir9FWei7wRlsCjtmkKsbVg95ktstLEVFTJqCsVT
Uw1LfAj87Cxb9LAKd/FOTTfX1N3OSOwl4kjoyU45alWszTqoXFgu1G9nuqOo485So/DNbivwiBEu
yYqgjxH4j+D35ACf+G+jKOawm4Zpm3lX58YeGQuUdlounw19dPXTjJ34ENjmWLveN7M3BEy+r6ZX
W90N3evAj5PGc4RQyE/Zvh3efoO7EAFyAf5NO18dx048/p/s4hfFgz6k73PAuv1M9F+6AgCRAgEk
Gn0v73DclOXQ1sdsTe16gYDbNtsp/KzBe4UAYxZnpavWV+B92RoNfOkeRcNSTpeRT352WCin5G6c
ng3mQ9gpWxxz4fGhc+psSVDRolzSEfH5g3jowkK8SU7zrJRGiv9wIAfD4rs+dh2RAiRh0qxFJTLA
MhdHhK+fgydNllELzHC/qsJeHyM4kQhFssSyxKSA40jBkS9F5ICS0b1nlZTwk77VUbXJ+TZbiNdn
pA90KBob488qBLOxYV8yiHJ7YOATU+v7X/nPFlQbos/Q3BeQoDWMjEhECmR0nOFWNdVIDzP6xRGf
msDyv3bgQrlovf/mizha5BV6P7Lc+RNwxTfibeyLBOzk7wNCS8y9u5WOWg8UURH5I6cp6sboV9MO
CK2CM2z7khm+FekDMz4iX3rmTdvAbhAqPUT4J60wLFrZ+HUYxkwvzgsCcnG0NIlj0abg1goeJcqq
7d6OAM4wBZyf5Hav5qVe9TFvpWndpWr9AEZV610Tiwz+1ZsYao7rdDhBxyn2VZ7+MHIEOuB0Zzep
acrVRKtsIqMcYfD/RZMZpiahAUBoBr8WvnwHRrinOrC10WzLiqE23ZN9jafw00hyHMf8YiyffiMx
+uyCqPDeCliLffFxjdEt5ukEo61CfXkCU1N3Ya0o+NydHuFBOWyysV0DQn+GTU2Yk8sjJ5riMkhH
Su78VxjuoWFvko8Q1MmwiFSyQwDqUrZbgSfGbTW6F1DI4XBKlXPff7Oswuft7s2reL3xOYmh8FNA
vng5Mjabur/5wbQTn9wuHad3y5nwbHc/dVJcUDKiL+VaEdwLGwTMMILat9UM2Lj/cB1/J31bshBB
wT88UaDbAJ6zh4nHO+0R35y/Kag3ZD/8Hj56eQLJpvQdOmGQR+TZl40/hyznhpg/NPhCLHMFvpcZ
CW29+uQgRp3MzkK0Qo3b2E898+x4RuStO1GxyrNZRytkCU/2RhR6EHln7PAyQ7YUdq+DrhaMk/wK
4UTteqEZNaCk6Ve/MDYaEUl0AJZUydDjQ9ugYmzHMJM2QccRgkmvjyX6CZBUB0em352hfKmYHb6e
56FJYBNXRNRDXt9hXf8kgINQj6X3TTA9scDsHeMWx8TS1g6zt9UFydvgwszAAWgRWq65xvUnIKwx
Aan+RXXayXiklTw1NK2jdeIzz8aWmrULC72z+E4keiKxlSwhkHsLCyMrIJ5PZ2io0uA9C/F2mBbD
YXwoMJjX7j1ZBG2Votsf4MBpL0khJygniUGJKlGmFVjFwo7TTG65dT8bQenWXC2+x84XZ6pt/cf5
lEoqrPSqh2J8NEDG3+Xem5R6AVbavaAiqUPsSPEmZf3T0DLgXjZSq+5gE66wvgGvTtb5Z3RDrrTT
2RkWokwESDF4cMJJ4+8Y9n1lJGVpztNKladms2nQTkl9fRK4UgIGYW5OyQXfk2LQCFPMq8bb8lky
EN2oWQNnBVHsBGK+OdKGWtVzc9TTJXGMdzAKNNZrdY21TCACa63IaD7NCcZrPtO4JqNQ2vVv8A+o
UH2tAyrTSq8zvuR7In8Va83GAPQQc7yDPWCUMUBKzXGScazEEXuoyNM4yBhJfD1eTrS0yzui/VMz
Bnaq28P4feKEFdtbfk4dPs2c9lPVEotxKkR8zHHVhMJOUVGawnXnPX3NHyWWaSt8D3XJmdBMRAJX
8MCJ/b+RVBGyQAxtIRA38upKeVLlqnoqQj/3GFUwSt/wAvB90DMXWyAwL5O4L6y7k9xRTwPxFfoh
tFOWMteGOnJb/rKITAHKVLBk7u142MUuekylyhIaBhHKhLsnB8WZayq+4E95fmyGI0uFZzG5/eyB
X+2f2ZbB7K7yq9z9AmREHc4PrduDbSVPpuAq1Ktidw0O3MIXgmpKopgGpcBUvQB8s+lIP5UK2/4X
Xt/GsXMTO7knq5ypIqVtB8to2J0O7EvzyQwTIc+MVi06yreFZPdM4IyMkl4sw9LJHjhUfQXg4bXM
M+CgXW4oIqxae7Va3r4F/XKTu7PNMh+IJnqG+H8x1f9IioBK4vakTKo4SQ2WWbxI4aJ0Yk2FQcUw
cCf1NAK7JlvjFEi70MRQdtw22ectYbAdOm3HrnE8Egy+a7cK9S6YbyX7HXcWsEn4leCM5dyPbdb0
XlAsigsRd7c95D2lpT1dS8unNRMNOz4babKRKCqDNuw06U/FecuMVRIhJORg/vamwMavELGvl+JF
ymjclFpgX4LrLoikc9lQjv79aiJeIglwal3b/Hs8N8Z/qsBT+5lPomHUkVI92wyT7VN+0HFFrbFQ
Ztlf/wgEi4S3R5fq+uYu57SfJTKfLxqQA3PsmDJU0txXp0t71giBssYOLvj/cT53bZG9P/B/veVo
kYzGU9w7SDZymjdOx9cn32d1k/OhhzVv/UcI9nNrjcb7pgllvkPUOwfaA1N+J8lcxog+N8DEq3YM
ITBSPLiIxf4OLUBJydwR2i4FPWpjpX9LEgbbr+udePk3+SLsAVX/XPCuDLXxhF5E3UKM0YVYjjvc
G1f8uKDrwhOFN9g7X/1H+cgwG+CwpnrlVzDoGLUKghMAUnNkwWN1hdKEbyCRYlJnJXXdAoD90QDy
VAWkCVuB4rKOEjMTvaA/bVO1HxPb4FYl7ueDm5mXy7+WYUrVbkvygIGEKUXgL0XS78f3B1u/sSgb
0qPZWEH3QjZwAuX3lEBEckbMHPgJZ8CmEhfzk3WOn6OCg4FaDs9lRu0WMGtHnHG2UaCZo81bEa/r
ri1MFQFVfK5uyZTjQzhvArmMH4882FpCRiCKnsrrJ1+nYf092od9T+vMT3ilOAJ70frFu6zdsOYf
AmXrCmoPUyctml7IoPE1q91H0Voa0jnIQF1VL4Npwr3FybE2a6KGLfETB8gkQOBNkuk+eKBqorgr
enIh2y/wA4mWMD7Tvx3eF8+/dNiyQpiRRR055zjpROoyJX21kvIS6Qd5y7VEzGSSPqRGHiYSrhf0
UL0O7g+ImMWtaXLwdOKcooeJ9UeqatcNevQiDMqE8fzsp6wzgRLmmqTCsKb/6SEEuHls+rlyOdg+
sDcfAK48ykYMIW+O4VyU3TyjWGxm2oa3loFEUfiZMRi4g+P21iZIrUrx8RZy9RjnMiK/v5Hvq5MK
k4X1jiT2NntUTmkzCpr6foob+IuUNGUlfsjLxTrp6+/DR1dbsYj2BpnK+xGPJ0j2znJrw5nTwOE6
slrHIISkohdARFtwhQ+Tkx9IufgDDsuPB5QbiEYNufbsrXZAjugMlZLZBlyjl12SLYqDyVLpHC9q
Znz4juwvYxCQQreuYhdX8vI1TttnovGz11NW1ci98/jMTxpMTMwwtF/oT2zEr/quQQZpNqBhgdqF
ouhArV9bc98dyZiB3yjoqvXWJpEb9rUppECu9NJoayPHElI0O7jUs6sji41w8tS2OcMzgCDF8wpC
yXuJqo7ZAW7iGIdEWLrOHohGW2Uz+6twDd5tkVU729TxcJcbA0UHoYtr3CW/UkFJz0ufYARa7s8h
deqNz8aM7Uakn7jS3hjiEsT2J50qLbdOIcbNEhVHhSzvIWM8wfVSEMu3+LNQe6KJXCuPn+yf7btm
Ruwdm5uzkfn/4F3OZngkP+Q4vKLt4xZwZJe4dubqn4eRiEr4dPLI4AjQRp6iP67yY0jYOwSaS2tn
rDpak7lAdwnsWJtxtei2Qnx/WgHSlHeZIUSzNAViL3fsKp3h0QlT7/q9qo/zEoyw78ddJAo7RTcm
9HH1esoXmdy7e6MY3vM1puJS10F5bN/+xtkd5qjw7UEc6OxZqU2Dh7THWYeNGXTsj79m4y3xsvlQ
Up0gDiAfAuuhSCdlqnb1aIDy5OxQ3bmeSBgAscw6Zx8Ulvsm4cR+qZ5BvnHZNlyt6UmBiW06Msmt
Sq6lh+8Ssxfeg0cI4GQkk0DU/Tmurzd1/oL3VMXTMGyViIdsX0pQkMfwJw5ibAY+OLEcDzNdecj7
cgVdx8jgJklajuu2wZ++TSu8fqXdnE/KAAgn0wlVy7wHwdCw0DwIGw+GabLLNOXfny6iXiIww839
VKaKL9BsqCxnukfZo7vf3XEafnrFK/1jSYd+wAtTH8yjFNpGRyGllVLXHOy4FpNFiRhLArMGkQbE
/4evvIXr2P+aUjb9T6egB5oEi4GOYHo8vaF6AD9uIf7LIpPyT0oQMxtEJGheWpSVOWzVxpa5HgTV
jnln68X7gYKsfEKWgfZJN/439SR79ZZ7SHce93/dmhlqrPGNRa2NLe5l1qlrX/Ak9F84/fap838c
K9K4GXdtAtTYg/ncHK5QiGucjJTg3idVacQOZY++cz0bmGccegU0q0nnBaVDMEa+2+XxJBrHdwv4
ybciuUZoovY6KgH7KWaxiuL+Ige3Nzx0Mefr6zd6DhSPZsqHqJZzmar07/Y/3ptQ9+FLeM0K1S6c
6RLtF+K+EpxKEb5rIlyLzroHG710Mpu2c39xWd2/W9GJuqa6T48wdB7x8NNYUGul14WUMm1r9flt
JUT/7b63xvp1YKGt39+zrV69dlbaI5rLGbIiTYtWJaAZ4xHwrkrucUccrWgSmdLCDWGhrChFaz7z
7/PymFJFcTSaRtS8Xe10Nr5zgrqDPkf9iK90LPVWQhxKaulPg88yOB027jguXMuQZCdEEJmpqQQ3
1bfwLfhCdAlcNYrw0NAO2RxgkBc0s3Qs/rdeWcpxmohKc/BU7s+Y7Ga3LzTxzyjqSRADihuVVmyc
uyNf2FzZ8y9H3NMDzP1Nz+xnM38OrjJAK1cxNgc0V3QLc4ASqi6fa4C3OPp+iLbggWTOBZyjKEVH
sNPCeHaUHIm4I0o6VEuwPjIPwq/i3GUe6CJucccw6EWLSyg+xnVvuU0ie1ceTsNmiwII95Q+wSFr
s4dla4Hl2zGvFpDwCasagtmyMJgiwqNwq4n81zVkBLd6o8sT+gmzFVqvgfvR6mqRnbSPfSHLyy1M
QNwu2TKLxyXxUWwIf44buV27xXICRhC5pGty3my7MlEd9EFJLvKgncMpQ2moms23mzR+fRxZ2dXT
TkhT9V/FSfY1Wdg4PAPgOSk6OHnnu17qO8vJwWVyoVqTQHYRnUGcifIxbhg3h/p3vbg3clZQ1IT2
7MDAuIKeqwbqYjgKTI9s9RR/07HcxjrAmZ5hG21KaAmntNQGg3mGYTQ/wFfrd5HB7D0ffhiZVpV6
Cf8HD8/BVNuiuajSaMkV4Z4xZgebxPB3ePn7t9/LPV+Om2OoUsy2xgSr3rPsH525ZAPMPMr++TXn
eSYcZqRjCBo504RgbHce7Cz6ma8gncKFlnszcbs6DjQF0IgakTYVJiEyUHe4f6xH1mBgiZ5gxoti
K2u/oY5BSx/PozdOY0Sfpm3cjaVjJ2iIavNw3sgLtQyi9a+XIbEiSr1WLt8xaoQ25FnbyO5stRtk
xIBxULrbT6iVB3UbkctmloPpTREnqFLIjy7yzu2XGbSglA1LpsHCJwFP6bZm+qL51NAlpQCQcCs4
oCvZ1+IPW2PR1hVtvRD3eOqVOBG2EFTHnnT6EDDuh/iW6J757pRO0YzEM2xqmFtWAIneHI664l8o
FY8Ch1eOwUPHQlfXlCO+S51IYT8tu10Ad5ARCl95KVn1u40FctMoftQ3dWaYtYfjnlg+0mhh44Rq
Hasqi3OoR6sR/svmK/XGMwKnjGequ9q8uTKMaa7DJQLUDBva3A1BF0sTh5Lui5/13mlhRTu4E2Ni
puM4SboG0D52PP0+rJy13EQZ4pG2qukRYxTlULWUgT0nCakttTaQgvayDyrvzbYnIhjHZzotkFpb
avbty+GtQC1UIJhXrkpuNUP0etoSb8ztxiB/c0ZX26LLk2rOAJmsO6ehX7b6XS12v8E/4Tr4VKI7
XYXSrSwMXap+m1g6IH/oz/ySvy0eSQzKaHxZhAlDeVgouNUXYl39FDoDWtD0dLKEghWQOiORCS3S
tiW+5wLuILdUmvtckgJdDuiC04aY1phSfNMDbjfhdPQUH8axq6dd/YMJVJRcJqwEN6MqJNLvnXSn
nLIQAtYKZQOWZEIkKpfqUh09VyZvE7Gym3APwbgt/64eE+rZyx5ET0BUDyY6JwF5MurAQs5ChFO8
25yZeIx6+PJpdjvBUHeW/q3Rb/nWACnVJswK5bx83Fvla55N6aHroYp2c7x8NfVs7SRX8HuvwBbK
g6XvsFc/TnDvURDGTE/lKQye2auQP1d/3wmklykBmE10wY3AjfgsWZlRTbq2xMJYVQyi8pIr6D/K
P2AmQHEIFdr2VOrsP+ydfuECtjsIrPgTQ/LGtlCK9VcCdgJPPDEgZw3UIvZ5IW8Xd0C3EJFi6RGh
Kzo/W9HHkZbdcPfJPxxOt/Il1omeVOVikPVU6LcGDN2NZVVE2UqCgIuJocv0ApUSOVdh8XI3OKUn
SCr1IPI6vul0S5JWmYndtK7MISWRVT37AOZ8BiJtPChoIlJhBSw6MG0zxMpjUuoCdN3AGYX0SNqG
aNvPF6Bj3ksrmwKy7CFIh/F3vvG7CtPTt0bYax/QkiLs17tgA3DuyeiQU/Ub+2ISlKvypO8hSRPc
J2XNOg8guVLNnaAPanMahOFqba9U5h9tsocxV6cjryDvL/Onw1tE8gqMvxpmtQwzIgpnc6Y9+K1R
8DA0qtNoQ3+SjrB9IxyG7LOLwpZTCIs494HmHP11xasjxONmcXM2WZ406snh6gLdc/m1sazdNQaP
YbQ1RL0tY3KClq4vaQ3/0miOxDEVF0bZ0Cpok1oCeN7xz3zNkLvrJ8wLLIwXVKUfCDoYvrff6HmO
C0RoBg/jFyHqiGklgl0hZj9zryNSb2mFqiAGNwDfMgXQMlgi61y8F5EVc1AyCk91qncYvmneupJ/
Xb1fzeHY/A+nnpm0Ipy1eBVxE1Iy51WvFHBEjN61ST1+QRlFKYTVbDvTHd6mcpcwRhilArHpl9lp
ygzMP60Cucre0/ybPwit0ZzBJcv/ZqoMkEDHfxvYCahwt382183xGaxsPuDXRzs0Q5i+/cqH0WQq
psdqgEDYpo8UxIYHxzI3nRjviDYcJYiTODADInaDEabYqPkiDJQLSkMZ8Ow+6U1TcprmwHSUfF4+
Ayul9KXr2pza0fr35UEtonk8s27Um3q6FoIDt4jSE1atOx8B+NmyQyyE1EY/0qqYKnLb6P5bf68e
v/2LkO00ispeg9Kiruhh2k0PGwQQNBapgpRyAKtevQdwsLeGkmrEm3qA9Kw1micVw+yuazqR+Lg3
tDAOROVlgtvwzBjFkzzfXdOOQokvgxjP5ClZNbi+zrYSfXgkkmFocYN38ZPJTYXiiEdIzD1DTfu/
/5raGVx8f31vu8Vv3saDK+TbePFBn6lh3xocXyZzyMzelsiirzVq9kNAcXqpSd8uAcMAM914O4bH
4Z5xiqtZGmmcCO2JCGiGZ9kqSHv5byNy33O8ELULVE/3reg9hyADPDWuRCi4mCDvlNgtD5O/AqQw
XhMZiLuOvXyGQR5KqYxQwlCTUPlxlkJtiBeDYoyOFXqpQCSfF7ZXFtIIfO1vqga+Em7ytUq1DhWd
lQF6RlRm5EqUkAD+8FBzSpm2oAHpzNL02kseQpRu80ixWxgt1NUcAlR05RkjQsIJPBpmt7zfsNoP
Ues0vRgHGJ/JM/kXjmXcsOGojoTIHEBqscWmIOD4gQaAeYQLB/al+qAy1zYIbFGgrsFkNQQLG9ht
dK/NmQjRrgHHdXQH+z5NOgFZLM8QqKCuW3Paw73ssOfYi5VF1iNiqHmum7Uw97fS5ytimBRSqJaZ
Eqwp7nodtIT1xVTJLPgdfiC9Chq5PLnuNiAL5K7Z8eGeJsTlnz8XdD5cGDYTjn7DtnZg3Dow7SqS
JyyD5TMllVAOwMsiQ9XUx4H27RN3mEwxZ0PMllkCBDZiaa54cTwD+7Rzmws/TrLHX5H3IiaaYizW
MqstF2y9g3MtyWfaGRglsiwGHfrEEUWZrWR8psRq6PJLyB4V8rOTXbyQ1tPCmeyFkBzA5uJS/Vhc
OdWKvjG1fart+Qv8J8ZI60sVY3gkwJ6OLu+LRmpupFWNK4Cnf/8krluOYdhsAfPds9wBIt4lT/2z
mhavNBD4l5oOVvju2tHUNrsewK2KO6k1Sed5K68XPBckdmtXKyGVefQmlhoakLGqUMxq1ElaPtbI
XrKKSxTITFxI4TraCZH5vWLqlfZjo0T0Wwvj1opQyXx1z0eN48ttwYgQjtkdJ2Ve3X8jrk91FcMg
3PbnF0RFqqdOTLvFQaMZvETId+7m4pgJ0qPs1VCbWuzxzRVYNfdRSigR3fHDnWpPnpRbGmAIRurt
gUEDqg52oTBOmJHHifG1t6hcCSBUR1/j3qlEnILalEjHcpk81wuR0cfAUehf+eEieHRAkATMTZE6
DItE2KXIM9OANqjmw6L5Qk97UDD8fn/7pRQs2jnFPO5PCoziF2gpyUt8VEvMUaHWUoHxL0KuxaUK
gj6QlfSpQ9kgETT3Q80mG1155Z1YfvfNZHHtEYtzEkUAAKGn62va2/Bv/KEGPSfg0HasgBJ8fGq7
HIkR7Zsk4RtmP0g3S0a2s0MLecg+Mto+HuOntm/KnkQVMSRMxJQayz+MSY6Y6Cvqbd7pnSi5dAsP
BmaVvZ6GkMTmF56MG3ZiY71mhn9w2qzF76szdDQGMoHysvmPbH6sKfCIfSWQGaJBwvV4k97TZR20
0CGdUFFMDt1Mmv6U68sCw9OkUkQ0Frr8+F+MDXau+klgt2xzzZ3vOzgJRPaUx1nCu1+7qPxkq5Bz
wOx5GeMQOs6rY37R1wXgStezkkKgWGf0d2jtnRDwx873CLFsFlIQG1h/tlCXzScyHc7VF6Ve31sd
h/g1kU4ptYS59Yw363z40H7Y94oSLTKN1fEyuC7RbJdi4VFgjCIHUTf+kZbY4PDg7+xOrsMWU44Q
V7Za323H/DqbS7sGL9OLADbuMdO5bDyI6ftWRZbk0zb6zcFaF65i2dPgV3EWfVvfD956LdzvMLm7
HUqjELWpAjFtmSS0y53VrHnJ/S5eDn8nU9ISbCN6YN3FJYzKUVxyhqK7Aw4QsrrYvhN7EnsctHE1
XJjKvzNy5ECQycnbAp343tLb3GmpHZGJ6Z5Do/jlT8CfC7dCUCCgSP46MzEOJQuvAjENGNSpwhrN
V5VSZucDmZVP6+9jNB6zy54yFyv2NgbOpemnUwef1D5Xrf5VAcyny0ZYcD885GZelgxd28OA7I8x
uTjrrK7Dvr5EapQjoMWURVY4jbrrc5O5M1yhB7n5Qr4iBwnNI6EKRPN5tK0WNtA/r/Yd/KhZ1MM3
lQBo/Q8XAo0tX8lXocNjiQ41oWbw29nqyVjQjZh9tb/MF38dl6EcwhASRJOvlhBfrlMLqX11ic/2
YGkm0TkWI7q91qcObjvZsFnVR4myQYu8LoLKz3kT1hGnQEXks8WU6IAm9fi3m6vX5wP/rrYogv4v
ZZyLr0p7l5RiNFI2nQH9v1DUHhcf4bFGpbP+E9Q+TVgOcZqQxRgHsC1Ig4aXtvE/6ZQ9VdcGfkpO
H0UfuNowiQVe+LAmn30+8O/yxY/uVga1jRheHlZsoqo2iD3zApIHCmJzV1wgZHec5NhFwArwNjdJ
jqQRLetZHmpJ56zcprqY55isfhs/hKY5F7ZCsHyhf3lDGO16Ia6cOimBm9ayu4+Wres0epSpiAFg
yVtNEd5ZuQa9qHb4oJ12yY9VDyLIX5VAeNiLzi8KSk1w9qHPxL1H5eTrbFDNgROCLBvRavOUMYQX
sH+Ilg27ktfjTRfHAsP/kwteRS8qQNi+WQZdqAVdDz3RT9h/Tr6ktz6NwlOUUQAIHFQGiEYA4ayZ
u0+bbhzLP7XBjWIz+QqjemR3ZOoeAENxGeS+roCGtZK3OS0Vxl+ewv46POi1dn+vnKidVgHswMMJ
aGUbwXPNebsOPazFJ6Ve5tj5YdwLO0b02Fr9z+KYaP46rS5k4wZKNSDVjn8FxW4jxhMSHZY95GLa
Oqf6df+YuivP7oSSoO4EoXoNtssWopq8P6UXhwh1z0X0x8vgt0no+ruxgwHL0TfAbhPmM4yFuu/r
xbLl3XF0uL2ky34TUTohMGjSPSIHt9P1mMf+8S0Vl2blxjQxDF4vvHAXaEMEZiymAhK2moUPlfHN
VZiZqehIiCVVNCv3+CfXDbn9iiC/uNiYqwNtvwq0XcBlAc2isLLZUHGxymJaOBcBma34Pn6OJysv
E9a7K007yFwHrgCBAMxd0WXv3KwJ53Y62rUpwOFUriiFFNnBocHCgPFTeJShAchAJ0/mRbbZeEbt
UApN0WTfl4qFSRcSJ1zIAAsxvLlhXbvby07nGBa7n+W0V5ZMUYm7gwUI9kAWyXxMwaGBX58nAZSs
J5WeaiCpoB4dmubGpqGsBdf25Uz3B2fDaImuOzgDQqUfoPg9rZcGp9wqUD7zZGl5bScd5piK9apu
+gpjuPyjfQIPngV94Mxh2manX1x6c787QkS133dexuo+pdPKKG9zziLLv19JA2XKS4u1EYi8YKMh
7Yv4qMNr1EKb16ngUHSZ7fQJ7ihUrXUP3geW0aA3HjZx4rFBacm/SiPpGKtqS4QODACYvCTP0KuM
srH+TKOFRLSPOUXNO7Q396SUSyRgECEdAjf0MvCfXYhWsqGor7hgPzcF7kOezcEgOhjZ+FqxLgj+
XsEGDnboG3fSj29M5njDTUq+9umRwB4LIubnaFDAS0pjUdNpsq9NkxhkiKdFiW9n3Az4ZyDht9w2
scrIhy4p4v9/5J+PIBrDtClVsBsuwspbqjYO2OQln7EBhvBlEhutuLX7muoSRpRPVDDBER5F9Ogz
LUEU0hPzV9ng2SQejpH/InFIVUNc5qlPgYMCQ3jCgxPG9bK6yq6Q9EOVdum4zPhWS3hIQ0mrnoJW
kQtkbvIuIp05VM/5XYSPKCBqiagHnLFYA/fIozQk7tdDOZj4QR4k0qL6pwQ66MdWM5DfdcIDcUcm
ydggro45MdbNGEe3ObCH8XG8R7WaR0FO9o+nIm2yZwZqnyHyU+xTe8I+5qnerjPtCgWI69K3GX+u
ymbfiUpMc8cq20FSoElVdm9sc381vb6FVmJxX9udBD4Y2ZJpH//GEwmpgUuZlgBvYr411yLPm3WC
4t2RWtWKiVL9leMt13cSeTvFt/u3zT4jQiOGUnHUsB31cWEIaBhYhQ7WpkX8aKlLSgfBJoVfKCVi
tGyhqi0KGAldUBt+uMu55twHI3Q6/xJL0n5eDY+zpNzf9lnz3SoRnIQWCZy1DjNkdbOrfiZhE4AA
KVSKxkzwKkQF5gwut8IugxUmAhC1n1dMYITIaA85Kr+/XCzlzzelCEmmOuKi4mHcRh3NyOwHeTfD
BjKxKk0K83EN+lg+FgKM3jUyZWAJRwLKmgww+OLJRakNXCEO9WzDUMQsmron1oizGXCr52BfZ9GY
TyadDy1VuJMqb7L4YOwq1LeHmzHNab43pPv2vtbDU6BKftlRauwgKmbm55Qs3z/awjU7BKkXPzmY
9HQe7BbHQM7pPNi/dvrFYMmD4+KPHRNeKH0eqk+YhI8afWWybvr+UzvanDAHY0QPHG84SyUwx0Mi
/fCCaGPhHWKuUrEJxsCjWOgD5HEilob/l9QIRSHRcXPJFAd76jASL3mJTpJgVNOmF2a4jY0GQh4A
mMx3LRNsmBuDvA8IjHkKaolskEvX12DOFuj6ked3jHS/bSP/6qdPZfA+0V1usVy5YnOFXUTFMj9P
E7R0X+RyBAV95bwnwGiiXZcu4+pactxt5ELOYSeUZUTUAnHWq/pk2wo+i8RBfiXHw+TJVl/Z+533
iAx2yMeto+N64qDSBWuT26usXBw+ojQJSP5KHISCLKdNeaPA/RqrRFrNN8TgepPUtISpQbOJSNyw
jctBLR3xdBtV9EAS4W0fdzgZPGfIIjK1VzF4AszOypTRcKzve4bYZ6lTsG1cUszTiCg8zV9zq9G2
SLqP9avSjovD0mCMAQmPCapwh5rn9YUR+wJj/Erh8yO1lB/Ln9iJBkcekXps3+ChKx+Abcfef7p6
kMQaUiA4/lnodrI1IDgvVV4f47A7wE9SW8gbyJS3IuLzcaibsvHuP/rcBZB0Hoh7EWnpMT43Ixmd
42IDauag1G6dhGpObufnU/8rY1SKRHhULZO6UHYb13brF4f5JCn+LjUKi0PbdqGw4BS0xEK6DqYG
vmxcOneybcNVUEQ6LttSoov08OUn64iq1zvuA72k2PVHX0u4YIb3PLC0+yMQ6NOhY+WNzFnWsCBo
lJGNpuwew6mbrH5efGKlQQq0faefsguG96ZsaHDabkOQe6chXtW7tpkBUTb8SDvFuxNIOjJMbIIy
n28caF8VVVGhiFMbWudSGnxxG2WhFq4QO/mvLTMF2pSVGc80SKeaFGx5yzfWucYRm8xiUz34rMYn
d+LAvcYrbwMdtvPxixtdDienMJxlyjb6pDPfwyofkgRRMyHQvQO/QC4fa1nRir2qYRE/7Sd4OEN3
0rzhwG4nyU5BBKsm+GUGKV81n672cKr564En/sVpLSfGzaG0fpOcjVGITd77NYRXLAAZOPHAFToS
D8pFPEme6lsFjwwnxA1ysPUFtmiTOkvN/9zHIdXw7C7Uc3yR71Wj9WkpBRM+ZxlwKfnP4WpRlUQH
2Fs2JMCuQ6EKQRI7OvyKuhYn64W8xsRHY0R2acql7GgWaRr36XrLSks2/kPQG5p+L2PRkRILyv2I
mlaLo/kw5fqbl/6MiWn0tfc5Vfsrkemg8ekcOdQ38rJQ5hiCNYdub08LwtbbYdvUC1/Z/Q/CELa2
m7jTBW66favsgGuR4OTXwddiHQXDpKYMndJAV2Y1Az+GEoJv8/d9+B1lvrXYEZLvJW2nOSWT5dZc
62OL4aCzrer1pdMlTwtTsDh68/BiDPwdNrhQ+4v3QqK0KDNE+NL3YAyPjEBunzIc0RoYhdn4jKkz
bgRPDaUzmiGPLWvtShA0vWL4g+LudhRtG43DCat1ajiXRXr46cB91lMO+eFekWTHMdpiyT75Droc
VvR9bvvzOG87pExau5XdI6oDhALNh14aOj2DrJDO+lRW63VA0Wgu7pIXcNitVr+CRtRhZ8VE878M
XbsckbJuDR2cV5nuOKpwtS7VvBbiVvv+BhuLIyCA+RVHRt8TpPxm0UkEMj8X+HO7AxmF8FvFXC7K
hDV6JAA5GzVbYJD1CWunKDx84Cq0MUnNaNVKqa5Yg91YGlg9I2i4iXwU9pO1Z+ewD1n8DrS1T09L
6tK6SKzp+ZuU3gETX1QYiP+yt9kTDILZ9cocOmmQALgLn9ymMC/9eQhSYQr3/2X1QZvHCtOGN1I7
xwCqzCekhJ/5RG7GwrvH+LVBNYMH351KDzf4hA6Jmx//XTx0eG0UB4TJF6uzQc7SHuYaye27e4ku
xtKfW4YuWsa4Oy5dmgV1LPtZIVkzmjrLNCl5liR2dIBSky2lag0fY5XHzOuFFaPzpaMISFc995eA
E4hkm22DjD4kzUr/J5uqREO2iXXJnHYM1unX+yJvDKuKpGok/sUmx30mVGj2uhvQ13XAYwA0rR8F
QIcDAM3TBDqx9e7eI1Q5FQgFEgFe5uRDKmZ8qA4yDiMMYDhI+5ylKginriOMIKoQCEnrf5cOgSlg
+MkwpV728eJ3tVwBiukOZfSRf+Qajd2+pXwmPp8Ggmr8g5r1MFRFWY9RGocrpr50S+E1ITCGGbr1
ZnUKIS5FGsUtm9qqSKykUg2ALJNR5oz5VaiajOp3ZT0oE7wFRv7eAFX1wbfFxG9rKKXiwZPIDRnA
ixh8hydJ7z8PAzyYPfUgCAsC2Ql20QEMWIZDRVDAOR0kf9qKjcX2E6k29Byteahg5nyzBikMcc0I
w3jH3yshiErkQmxvlcwJ7ipYq21vW8YlC+UduBHx0ZMRhOgv38E4sTcn/HxNmvchIiTg8VM/rTfW
EFo8QfZ/je9A2zW5T2WTAffnKqPqFmV8+/kgjdouNbGRWB7piUtBAutu5RFW+kGJfRBXwlZoQ5JF
QmXpvOT85Hmp5rX+hxFUSFtCqsXSiMtMQRC9IPWkXydxFoQSqdU4F8l0hTPjXTWytJkGuo9uctwv
aebM/Op7/HyiqEdWOfvMqzqdq7yL8TwVtN+nNUJ0f/btzLztaF3Dg36dcMEB7h1h57pHMIgAoDID
+3pyFnKp1L4gcFdjcX80LdVe0MuujSjl1IRCw39oUxyQH5J4G0aIoCZiS+FSdtCd6uP4huAL2AHJ
laN1WhpKmPnU9lZszdU/sUrX8JwHcn/FrAPXvV/LIg9/0hqPhAtHV8IvdkWVHRSs3QxIXYr4NjyW
8OgXxquFPyY7OR290vHwL4hLRX94xqg8ly5xnzPlSd6hC6GngOwg5pHdUqDTaNuPwEx5pXMxgkop
ovf3caxkyDo/f/sFB5EVtCpVdnpOj+X+K5DAfEjHhHM3CoUWq7EuKkkhjiOtTUFkTfRJrifCTdRf
eN3/7NeELdSI/KQFAoCFfIA8zvHVy35TXRrLhhLdA1vP5+vvoOa9Xbf70rM0E46LHrWkNTc+pWfg
bIOv4au/WnwVMfH2QdsIv6RlooSlny+/KN+SUGlR8cfFOJMsXHgXcq94QZoI515WOX0xCuqkUh21
v/r1oPag5UzZo4G9gSgcA1QoG8cOw9niGu3KRUpYhWdRQEBVa2+Zg/tnFcJbetQZGe+U4o1LTKFV
ylPbpKHTKVgjShk7/Kqew7kV3Y5Sn810dZ5Bx1dZy55BY2/xLgp8WE1SpQlaAvaDJ5ZHYwFwRMe5
JcqSrG/CiMyRfx3I1q4Er/nZqzAzBgiWXWHurtV0la4xx8+RMt/u8bo10TIfjG4FZa4FuLkFvkhU
FgbWuaUyAnJV+0ijIfc/nPyk4Hf+tyYt1mnsScvVT8mqgD0C5uKzrEuSfAmybiqncfhyS5nS5JTk
6Wf+KMD0yCeUckfFPJ6hXr3miZSMQ2c6WGgwQg5kJ1DWXauHn6UFGAV0+lIFv+rdr1U2HZt1XTyi
161YraZAifJPUMU+LtiwHsvYP3mi6BP8u5fbHlEH2yVYZL7T4uknPr83lersqeuS1E0DO+ptUjKM
moFT86SjYrBcxjBkjDkAmIEuQ8HVlEGg6FJYUuYaU9dA0LBSQIXjYTRGVYa8NbcKQTzFYIMplooe
WbSjh93fQaXdGvUtMeEevHQZD1CVKhWvWLzG8grbyIMrU5tFUmuyOkXFYKRQY7qjkomM0DJqSVjJ
tPPpQLN+4kTI4yxdbFu9qsrO/GA3tQKmUoi5FYbL11kuwnb5NDl7FgEvsPCeZFAN+qoVFOP3uZcr
Zjpr20emmkF7yqf3XNwqkNx0lHXWtnoB5LGLqS3RwUHj9zPbFzjZRfxtpLqpZiNaPDxuU6AdQJnS
pE8qVmvIZzPfNbt+V5hyzeJksiE3rYl2CsWDLujoUKZoIu6Kd6oJdtC7YbO724/Q9qa03t/Da6VF
z/hjkQnzV/odrWzNN2DKFcIbb7oLGJIK/g33EaYnUYeovwPmb3nzb88TZ+0XqwyLzOQF5k0hAr84
dUd/VSVzA02Kzquhz6f+QZA4YuOeEw57F3L4ppeLIw5UFFIdlDuKQ/W7ylzYyPesNrzA8KztjspA
nnwwl1h0s9/tt85EiQ9k40nba8yMf/d0o7QjHkk7BEvXq68fL4Yqcsvm+2ZqZIbILiT/GeQRVeqk
2gJZLVnSNpPqTlU2gRJa07aCOiPvVbIpUpuTRgCYtZtYqeG7aTedI9GQGbziBPvJaKJP6vHYnlQI
3LID2w2CKKQlXyWfDLT+uHyekGM7OSfAPifO2ArFa479FAC8pTzVB1uf7Z/HDjtW1EeKjgLqk5ZY
t4hnRXROcwnlWDkPfbtNmGNAK+h8KZz9hzOvnby0Lc/xjKLIiXchbQ6OS0pVnSG2UVHPeQx9kw/M
IeuOS0KEZUNF9ZV5HLmgfM1MNtbslCzc0le7BKjdWRdEBk7ZDqGwpqnzMKZ5DYTdD6inDzBPx8Ej
VCU9Js1r6mYcirClBVmZoElELn7IZe2aOkh6z7iMZynTA93UUqH6G5Jysi6knH1lmX3+asUKHrdb
OtNAm9ah9iPI9kzdaRPOu1Umoc0+VVBuChxvy6CXvmzjAJRwZqp6pAF/0948qSOgRxenSekCeDa8
3TBTOECUD5iwYiWzELcsByi1VxRYcXSz+tl1iX+dnwmVPDjV2P3PVie2b5l1Ppjqweif8lUb0RAy
byKSyYR9gdrDeq3UBXg2tkkYwat9/Y4p6kiLTyVUTxd5ntu3cVHdsP38WLDsXoge1D6Nki0JCzO+
v7DdtzKn311mtzz8rEWqx5eUAZD8CinkcrNFYBgMiadVa9Rm+mbbdOJ5/7uIl6fsAvLOKyEXwLnN
/ZeRJSVs6lEXn4DLLBVAbKpc9sFrgzX1FlkJYAPJL8tplEC5/EhY2xZnlVp8rpiHRJQTyTKjktAy
CEfBwHxVdru9hEM53KxoKRK6uDVl25/JogSaJmb5iQbM5ytWJNoKTIZ1w0N1f9Q4lAbhHK3Z8Tz4
lTskTItRPJs3X78L0Mc+H7qLVYFX77A06LlpxKmsGsOdp6bxKQ5CoLsadcnTCf2DpP5bgSo5QWor
JyuMTi3Qxwcn3XbIAI2guRUdMP7Khrht92SogfY8wbJkHDJNjX0Hp98UZYziI9hr0kvdlLTYBPun
rXPuYL12Xhhn2nLJj5BBRcMt8MXe5vEx3XIfkT9bmCJuC5Q2YVEU0FATHaPhRXtOaG0++v21EoqX
wN35wPYPjdgnNDc2OZS+mZNEL7C+izGYwce9hAxUhZ5IR3SKYW5CRJ8xz7/AeMZdoyfy/ImhAbrZ
I4a42CZA8Ap2sL9ZSOd02U/X0vLB5mOXhcmyEN1BdtbblMeHIQ3KUj8IidSdvXijsTAyYzPsv1cL
7OxrEx2vlN4dQ31I81N3c1L4FYLrMyuASPBX6KBTvl0JWfD+mGGLsDQQaqDulL/7ovJFfHRyFlzx
NvBmTalf0PaqAcubb9C52G02A0s7X+zde/5bWEASy6WSrHEaTwbFV6D8CB8RfZTwkeztwEu4cnXF
oUvNRuETy3YP7hbrN7bjtbEUkpZfslCFrBKywZvMR20qrRjnU05JaP43U+abvPsZ5nRN966lkut/
ASf3EI3igSe7hin7AfKdMh62H21uTmK+sLAlrSYYKmk/T7jFRULTirU47Bat/VnQo8MO55hDvfBi
r3UjyORZEzRzx8tLeKG7tOsGa4XES6hqC64MHblUVQthYq2j51s/ZIi3KKMXX1fxn/kFePVyXQYL
MWQAwzZPwRvUoF/kOb+7I+DBxGXASRmwXR6B9ClUznFxd7kyjAb8VEObNhAmzvnS3DGs4LC8/13M
7rDh5HWP3W0uhfwtTw48MkycXQGvvKCG9RPv4egBYRvfaLQ37hpL0baGNmdqvfg8Ul/GJ3KFowzX
Y1AgTWW657hQyD6j5007VT/8xP6f3RIWRde5Ecg4TEFYUqbEnCPbNkezMg+coqfRiR/Vy4Fj9kJr
dS+pn73bhUkpPjpgsiTZLdnMYsc7hNzM9hh4J39ZE5yv6vFTzD4b3N3H5keRKihFQ50/uKqxUaiR
F3wm7RKSb07A2GkATJICgxhcxPxxbY0FLw0hWJhhQq7gIqH24jMVPPdD4MbwJx04aKGi46M4aqZZ
oF8K+iFsZv+FnnqSxhWnROHi0eDDUczGrxq6sokd7DoxCHp/l29+1Z7AQl8xGknXDwTw1ugsIAGw
dHiG/DU3Nqf+7Bx05nLChp7kXck8yun9KiRawAbBV6Ehka36kssCRpqsPshwyE0cDy2U4/AVmJ/j
DyPLckTXfTCEqB5b3XQeNxoE6YuMQYk7SUdY2F02v2blOlUqJlm0+wnsnV54Gp8kCdaiLd/PFwNX
RzhkHTzumblHIXBB8M8ztuGzpurFsHPKb5h+nwsbDiyWB5yDBO2gqxrwo5wo7Ko3Z1sf0hDb3q4/
vrZEinNsuBLkX2R+cuWHpwfSfsWi42ws8WBXtU0v8PrhuQ/3PHgTubYh6enfV0XtVQgeC2yZt/iM
7UU8TCV3d6ZLoR3PVE0OEGdWhrrq2bzQRa/dghCUac3ajcExjlh4uwy5/9Rdterp7EkQwA/zmBJC
IFdhCvOqH7CL4PDscc+tYKgzNjgM2LM77Ev/sMRURdTLGRIclLQ8aVjyjeQ8UTXbE/Zof6jYDBU4
cNsA/Z5G29VOr4ffL/pgUYV6wjfeqfionQwKZ+vbjhIsZsyZJWOIyM0B5hxQU8QQZAk0MKh0fnT1
rzVqZQG4ghqnISXfKPDFrkS12Fc3AnIDN2Q0ThNIcnOqvGNM1b/ouyLgQGRGlcDBmq7nIW9WUTFg
f2HH1Q7fJoT2TrnTA+F6t4EDNnjNQa6jfRzB5dRuIcwhE51R2KY2pf5cAQm9wBYbH22W215llV50
0D9xBAHMysCXsyCnY8d0ikCtYWC8Rh3J0zXdybcVIg/XVYbBkV05ILO9aZ0HKKmMnhgt2bstbUkY
1M60SoSqxI6prWd+gsPyAgiRe93lr40OVc9IvLdOJ1FAd1k3HaY0NuUmh2RTQ0HYAbsO79Dh5FEt
FdGyLrS+u14depUoIleSJVnQq+dzHXH/ysplzPu5/ZcYNXD1CbV7gkpPjIZVxKYJybLgvpye8rcl
H0RnjHfJcYgagbVW6/b4RwJaYgGkQTxjO+ldIS/b3wVDpBa5d8QBpbc4FyzvCLiCCtCdJteDyKpa
Hn7B7OwaCfkE3VFsoDH2srh1jOHQZoOcbDMAgGTZ0R+54f7yoEBzhym5LRm4cjIeBX3xL0bh/1E5
hGKlps/EWPcYfekkBJIS8JD2wQX3XtidgYrV9VRU0hcYpFh+J5HBnjO5dixaWrvlYIf1CD1+jLsA
uD3aSr9g42DFSdXTxwjTjh5lMTq/Xs7RYFILfe4Zn5QBWj8IJ/CdUo6uQ+3CzyXWAdGyjV09VcbR
4WkSlzhJ72NrRd19fUXjR76o9ho2B4oK/7pBmywAxOBUFQDuBm7+nscwsivCmRLU79nR0EqDCl3v
YXcBikZRWEXpQea6EyXjWB75pEsl6VkRWCpE/H77Z3DUqD4qyzEXy00iE3MeH+6CsRIqXeWZH72Z
OJSENan8yIb0UyrzpJ/ainq64xvxVfTRMcOhgnegRnjjJJTWBZUy2S7DKrTr14Ymq/Rqt/fGhJGt
N0MT7ak4M3575i03B9H6tK7o0thN89+zdXd+LVpaYDUv7UqDDoBL7tkY2aO8yzR8crz9/STOyOup
QMru0s6lJwp58JqyktlS6aqc0fjbnP1nZjbtVG/Haic3PoJgMgZ35/NV1GDSnqPs1THWLFXVMM/f
JOvN8ErJn1Ma37iONKpfLrRMfPjk650tUrgBucB5DFLY4UJi3SgvZNcil2uUPsyaJnt/DbsXjKJ5
B40DV0v6NbJ/mljTl7sffJBcglvfQ6uMzBZXnEYO+qdP0mkQlIxJNej7fqFK34P4dgYR10fzM6Yw
wzyjDJnLikQZk91uQNRANFByVYILIXJXyqaM83log6xrEARongX5mI0b3IBA7XU4CQea5WUoXso5
BqtaB/zcAZu5IROPThVtaUVQtfebTf00Oa40rEuanVtiY03fD5jg+7oyhN1ye/bzBKwPWd5oKnLS
L7iu8NixRQ0wWKFmkjOyLzvAWKa2Q6ETx6dDQL1eYMUzsSOby67MrwtDF+AuLU1bQtkx4ifzREol
Y6ofe0tWH26kqAKq5/tBiWvrk/nKIDF4t8QyENU+tk0uWccfcCpIjWDZHFh358+vQcpVCQZhBuvJ
RNw0OR+MTl3PFy5FTI5l8eNFLtRYcabaVmYtLbz2N6U3J5sQ6h8Xh1cNJk98qvXyxIEzB25OtUhU
IlHLQc+jdV9F6oHxK3YqzveEEHbIChoqIw9OlYEX7fUerL6R7V50+dAn5qoma6WxVWKrgZFGiUj/
ceg8SfLcjlZR6dLnsJXVxP1zi6xSKuSs3Dza3n6b/yyklLfAgTjC87atGDtSKIUzy+6MWhdYVu0h
+D0U2+93fstLRk6nKW7+KiYQKs3Dz09uGPuKLZJt+TCL7knzCoG7oacTMW/Up9ykYQ37BhiQ+Omi
YG3gBw/fCpocKsJs6dDXuEGU1SWSAS2AOl9QIUlMMB2Jq1+5wzSKsqfyWasZx6BZ6ZGNwG/YrITG
sMEYl0IqquoAzBNDmv7VZXO5ncETIr5i4+CUoSq5P0Fh4xDaoqOeW0i0Y53kgYANcYG427YZaIgA
iGZRcnkmktRRIBxqY7ttVtKYWbyYihyFrUnqoBnDU1Jm/673TSYqArKsQAAquw6WwLdsMdFa27nD
olObvwvU7rISqSB+g6n85+8OHm/JscgGAmpBslo0IU8w1vue2kZtTzMSnj2sZDV+wV7iUqRvKTMh
rwXwo4eRYZatX202ujV+Fv4T4iVyWZNgC67MAjBUQVd4LGE727aRLop3tBUrMWUjgJ3hIzRzbf1K
T96rp7AiEteT5UIXHTLSwxerbsGQa4Rkx2ePVInCcy1S6bUr2coXSK2Df+EZrTI/jt2yVOSzZXuT
F6IHlyXkahfbwJR5poYHSTzsgFM7fa3uNxrP+5t48Ac1gSZHqwK1ofa7kl647TZT9FhddwnglHue
K+98biG2/Nl17P8l13OwliRJQZf9U1jqli3x2ZVSWSixyF7zvn2mRvvu3i4yxSSr6vAUXN1Dxmrq
kVsG/hyeN5dUYeV8kp2SjAbt+JdptM6yOSlWUcgPfULLV9kevspDyXIrWJ63QQz1d24g9EbZCDUP
QAJCLan8zyCeHF3SYnxnZJsHzQaS1bLO1gjaYrF/Sc5ekskiTbPxqn65TJ38Cf/4NL5iLPKfGl5H
iCW9ysiIlNc+d77aZOJAMYzqtMTNCVjaU3UL+5I0tUZWPGFUU8xK9tbkhb4TNdMzW4c3Iea15wPu
G2yXB6mzkeGwouc9vM8jYdab10JIwPWyvvK4VtxT4fcnjuIheSRO90n9Zl2Jkb441GYIi6e9YdSB
Z9SSc1ga/WZpBgE4NApfiM1y7Z87Q4i5kqG8/jITgNKs1eh/fSxka/SJf+yqflQ7zTTrHsWlwDjq
Fw7gu8fpS7ckzTHp5a5QbHtyoqUzdEXlKvmWNG7L0cUrenLkTF69eUdYhh1pMUPTc9C8PYKHZoll
6YljJtyEwXTd/MXc0sCW0q7rvfSxBKeZXh/GqXlSd01YJMpfc2lb/1Lx5cv35AvtSvUVEvMsz4wx
4xcwDYhQqrrc5mVlyTsAWmrxZFM0HhUnOajMIEnvo8CJvVeKQx/qpsMoe7g6TtYAgdt7NW2nyb2Z
hN1rCSWOH9SAXBrqUT4jOqDywdCQ5qPMHgCNmEEv5inK7MTiTnqQEOYBXjp3Obl73Y9RflapqusH
krIxpj9pVDBhW8eAVdyco0khRscMHrO3CXWhR7Khkr+nQDmEwvmGESFStrXIUYlSWyjIgxHsNlLY
RoGuGOzlPSSTHd1izSLUUY/YZrUlMAX9Czfo4vuEhpiv4AdkvRkBoNfdg3Ev//W0ZzJ1imF/yJFU
nZe6Oh1KoijqOw2WfBoOu3o4SRUsiUObXsvdT6ZiVdaXvPRkaP9CgFO1SGPwxHtJVhzBHVYML40O
0Z9NIKUSl58cIgdd/fBQXmBZcOT1V0uUuU7n2Rv0xpBuK20vvrB1KgDnlGPVr+dluvjkElmIIrag
98LKPHTd/L+eAUk1CWcdVOHI1JYYQnHxYWh9d4NLrSv3RXL+5DR0PpoEJbWG/G5JSNoYWZZ7syCC
w3UiNgTHRJItPLy15/xGQvrcoUp+nOWZvn1aEPWLvklk563U1r75FHam6wyEJhLG7fozq0OVBq0i
y1LEnce4yedcVp+ly8bRPEC1Y9kaWCS9Q2jT3GoIwqdLrXiw/k91xqI5/lrISVZro+6B+pM/U02H
Sx8xA2l0w1GL+eU778ZcPOI4ZJebhSNkqZEhYTAH9sE65Q3m/5E0CaQMI/0ZyTvKh8ge1Bt9rLxA
tRrriCm8LGNsJd7TxdXAnschrCSYEcMj5xl1KRFFJ1Z7IHQs4gluOWKK9LwOoa+mynV2YZxE9HVY
OPLOiSlIWIbB6bQcMDM8lDidJhubLujWPsw7v26TNdF73CWCzH0AFCttIBz5gcnxobsRmNR6PUCI
vpwBejQzSRRixVvA1yIgeZR+Ug8EOwBwDP6i3VXBJsw4iq90NbuVvZBQcWfWQvkCJlwUZPDg0RKq
LmHeZ0SJw0CvHEgrAS1tMlFjblW4zQ+BCXtyl/Gy/m9BYHzawJWS67q0N0rO2AhmAB4wH8SM+y2J
YT/P8JPJsplOSqhU3tmZSX0Jq+oNpju6h4d9Hk3v7vaTu2Cll85Eq7pMJZG69uyGT81JqqP2twCE
2sooMCJwGCjxWOg2TvquXDqD04FbolliuSVh1PRJfZo3RlAXX2RL2FQ+3Sls97KcOghOxyk3khBk
5xXCre1R9o2z98gYIgdiRgkM6HnYq5NB0jp+usu99hfSOWwgsbMa8RbAgGHL5bEidnIWqfh9vEiV
3Fq4aUWnzWkmUlcigM7W+7b61bzVgUPT8K0KiD1HqOxcBI9FQHo9NWjP2MtQ0jeo1Gh2MDnlAErC
0Qb6pggmUDrbe5Fjti0uXdZ4KQ3nsGLai5UGF0JuYnNKXA8DcFqhgX9PuNh7gusMGtm8XfHIUULB
kuN7845qbgb+zOF6hlBahIz7i/qjM4iPHPTAGGMhn2n9y98lJDhINCOnTF/vJVhdx5iJpLTuDbmY
T9zzzKQtWSVPBJvaGMZys38Ciu5TH3x6DiQQoJjfSo+tMB1Zww5OQ1h/mjt5yhgs5VUIW8rtJooJ
bB9oKiHWxB0UPl4UC+MhoVr/Zvw0WkMIu0N9Fm2YsfvYqCpSPcm4lfNv/dswscBIozsmhXt6xm7s
mwDnEmqqFJk99/Ogc9W5dyqbK5uZcOTLeRuiw6ica1Uqv5t+0sbDSzEy4Rwl84S7vOYtp4CuHRIy
7+S8jVW41QSBle/NsDhjvm6USg6WyoMN4nx9Tln+1NpGINm782u7Z6qfNOxHp8gIMXdgtwl5zubP
OYGLOOXhwrNghqiNnasmlaoUuJlehKpm1HApP+ye1br3MfWJmL+qo6AzhhgfUaoWnLBKwpVLBf1c
14LTKQpi0j3O6Neo1Ttsr1H6OVO8mRveb5dwLNkEx2nvtgjTu1Y5MCRUplYNBMveHebWSrWc6Z63
LlSrziSDM88wBLgvfmJ8czUvQEqENcCfssLYmTxxKtm3eXt/mEhOdxh6Ho6UDcsJjnCpzN0kKitp
+DTf4Md3dYqqBoaBtxNJ3UaHgbMf5wE/Gg3I//0s3N1D2DB1AEfwJUd+N+Ha10BPEiA2NOt7PgI8
qEqXFoWlU8kOgJ/V+UVvtSx7BiJXVEPDHMc40g/GhtWEEmxsfL5SzEX3Isco0TP3Fv/dlRv9gOy2
fLg28s1uyKmzgSnth79TVqC5pXY8L4q3kUvbGaUFXZ30iSWj8qkEr5zxw7G7pbl/ELvt300eCZdI
ktDIqXRRPwBJ+Vxl3fB+9NRJZXYd3+pDY4VsbV4SkYUvb2ZXr07yMWiqbCeJQ6HRDTI6D2iPmhtA
VdFqeizlismUyv1iYZ4UcCcabQFxoU4X/XLTusrwhpQSGn+SQfQsbLGJjssD2+sjH3L5r79GZ1Iq
0t+4k+dzRbCOda5Qtb0AMYd55KDZZ+Tkrnrf620U5D+nWg5wZLVZXq2kPcNK1ar9GzYdS8vftgzk
olht+kUzYRnxMXe7LnmPf6ypE9+sjrwyfTD3LiclJP4IjXXiVKWS1O3EZDafWSumr7ArSPT0tFu0
2s+ugMiARmob99iGRz/2/DgwgOmakrUmJNJodSwfobXNiHSGYevI0fJyfif36dHk39fbP4mTTzyf
aqhBrLs3bwW6P3c8hjol0GeWnFmxpNcWuBaD3is4trYCZ8iDba4JOjUA5vMrXDxMrUQ5ORSDc/iP
ea1/IM0f0xlXdnduoTT52nnEicWIVeaFQOx5XQXfrrNmWXsvnhPRT587pybZzpUKtZwu3e4X1rHN
uVqmKa+26XEvtCuaS702BpEnGUZrMlZv6wX/HH/W5FkBxoku0LRBL9l/dIlgb3nNCazZNGZY3H3q
CxMYsPz/OpgLkoFcQVDUFCHxjEuXBMEVwBlXjPUBQZqOOkdHKqq8NHLYtSGjeSlUWVsC9NZhd8f9
kYYhMCF6q6xXoqudjnEOpPRzPHZ4Lns6o1dbB4d9bz3WlTiitI0vtxB2kNmIR4sJWRVFFCbt9v/u
uL/K2yGgH2x2sphwhcyDVLaVSUuXJyOsUZxcJmqvX68knemK39IFg6hWIoZh72xfSTvfnpWJdcCG
7TnQfxMHNPiH9sox/9gzkrtSqKG/lQrYeFIyUBjrqj9Iq12KkNeQ1J0iencPNnt/b5Zvioix/KTj
TbPkNuRrBSnW5YohJX2OTv3mETTknw6AR88GB8qCY3nuEZ1z/iJkrBBj76tJex6LdO2JZy8SLlky
fJta8HlewegSqy67TYTQE98vk3T96CmTr8Vz49QhiabA8BPzZEjY2TSnXjcbq8rtL9XduiFzkHdC
DarRTkwT8oSZwxtfvMBNvbyZiZhSYiBD2yAj17rzlWqlQDvAVAJniCrXo6CSw7UP9QggfjFYgA7w
TmXOXFHFnVcBL2OQZnMYFu6tDE1GLPAfiLvPf11YGjhtPWJSyqKQU3/5w5qG8jo/bYQcpEO7/I29
qUtrv8ITtQ9H6sDX2Fc04U8h3K+FcetMqefpdOrYnY6yGL+8e2m/5sb7W7ah08CMkdyHXMagbtKl
gL4zhUtoscu8DwS1Le4zi0YqZ/zGHjEKmuQZwMxvKzRVppLy98xafcytq3IQW7wx/z07tpCvKCSB
2bnf+yi5wFrfWlGMTQk8LFpMSNxzD3ebMFNs3zsRmAkfOrFHCR2GLKug2BzAZoH32C1CKlICoXdO
w3UhPilqxUfL/XktCR+HYCiC74N6zC1NsDThk3I9DsjVGcRFMKJKixPoQk3Rux5ZVOMiCoOiFQ0o
lSaiFTJ/nGkBPU72S+TUXlSQGkX0YswSnZVX1koASgQUtntr5ntsVblDJ/hKcXldb9zEwTbccTJg
L2gLMf2mgGt6oVUAFsIMjEQjK0Chk1CPLp1aMZ2ar0u0THr84WoD8mbsgaIe0KFdte0W0TTh3Uf6
P9TdEcLN5lhaRPbhUL4syHkOGpxqhrznS/yAFjOTMhYKUjnJu037+ECNO7hgqQvzVKS3BZ6qeVJh
YH+KEk5rbYnjQTP4eyU5qAF43XIC4sxJ6DFex7/h59r1dFR7B6VPjqdHmurGqYggPSp/r+I31FUV
zx3EgOw9MQjuTywuk9CUtF81t02bc7ISw4fLjL84dehDbbnJ/ZlIfx+lp088QUjf4gR7o9z+CI+W
szuAx7VrmYOwDIYLOVmSPE92KBbySjb4g3Bu21Eh+zo6rvi51LhU9Zov2fY11FPegWPJRbDd0p6R
yXA4D0+Puvc02/MDrO0p1xQGr7LjICkjD6lKgm5PEP9zAlrU9TgnbOuZalvyuMpK5zom2G8yzm21
yAyDiDU/wrc4bzv26DgXpEIqeADOl38ZJHtr0Zfjsw9/UqR+O1In1KMKiHnwF1Deryk7uJR0SLQA
KwjIl1D/NbThjoCOtcBND/+Uoso5zECN86uz9QpjvLGT1yhs+wl8VikFNhDhfER1z7Dn+NJpBl+7
c98k1Q7Cck6VqZRh8y01X+aT6FvDGWereYFHwP27sqPITVKlGq7IeRYgnawC30jqjMWMdtvLqh4k
fc/eEK8fcpU5IHVSbxykqi7Yxba2/8Z9cTqvZ0nGMmybFUJFdPvpLpMev2Q8usWxG3IMsZXZeDMP
EX+gsAff281sbWMBMpRQx4R7eU4bmLkOSTDrfJSZTvI9/ThueKYK4UImn5d+M5FMNdZh8vUY//Ua
4wAgSQHWiwfFerPKLISG5FGfjmQGi5P/n3vSIfzMOS2KCfMCXuI0x68HA23ymnhe0X6U9uwm7+Ia
tkEv3p+rdBq5panBL8g8HJCilIBYXWi1ncLRMDsUwm7cP+vbDfNVCl9qysl6xoPqi8Gqcgv14GlJ
nAHATjoTFp0e2jsgdJIS3uruZfgqwwI5nI3KkIhJLeHdZo1acckwIk6PfoYN9EDCQN3YBKfqDeVp
nX1x/nyr4jnSgspPmhYU4sD65RA+9nrWsTV5sVqPXjYPMJWSbsl+7i4leUMSPn04PV0XlCzj6GAb
QnG7kojQ/NMaoQdlaSi210Lbyi0THcHDP2kJewnNfvOpwYj2F9OZadS/CYfGyS506DMjJwyYwk4r
wKYnaMjXv5ipn23oXzoE053g3DWzNEByf/3VRGia1euOxXqAUKh1FwYfFXsCA/aLTGGVu9YwsqZ1
eQU3L2+/CPj2IV2eGCBPS2NQSDNxlSzgpIODdDOpHil8NFf597/6+gXB37MsoHZV63EIP3lkIWVe
Phwo/c+wI8SBhmkNkeRaQg4nOJhM6DpDc9S9Uh4ZFqdZANRjFDodmRjs2pxkwzATGc/yiIyj0m7F
OuXDN+KORHaKdHnzkirfgsz119SJCW6DwUMWW9nFrcOlittJmFex4dd7Mb4Gmsuf2pXlPpZLybQ+
QQgdSr+9cDgIMSIpN6V/n1RZUWP5PR1LOQG1BvcaMN0GRs4fzYpdeMQLZRgKwJTuqYwD7yhJeSsa
vz6OOBLq6voVZpULdfskp/z7+kkN2zpoXuF47HgAtwHIRhzYOWNlNwEN5wRIlj2ihq2G1RfAGay8
Vukn5GJwZIZoYj4iDMdZSlTtVSU8j2+SKNzQyeZ7AcNxErV+R5RLoJUm3BplWzC9URtogY7grU1d
cBYH9yD0ouLrWJSrbbfyJdIkzxCr7ZjKqkXKbrlyTFhVmsJ8eLHCCR/3YYIPUO4frpEJCyn/aFSS
blMX549BA4le0Y3LDz7vuSPrm+NnUZQkwDPGSS7GxcDmBnUbn5tEu2g2RVmpLVHwQ7i3AFWjzld/
8ilHQ3p7yrJhL3HgUi+GgAr4EC+6ZRwlKJxGcgJyD0WdQaX0oD4chkTwS3ePm+aFWlGqjgdf4MGV
HH0ohJy5iHfMSPsMH/rBwnulwIT2QZd198pvCL96u1bVevjOo6VlHOxxOGBEGYEJeosNpipab9US
gWxAjVe8yCKlcHEwyc9ZQ7SE1eCWK/duM3RG5gDzme5G1TaFhsHgMRCfvxNR1IV0sqfHf8bibPti
dkrY2J8k51oBWRK7orFIq3D4ZmH7eRZ+wQzsMBX/7zNbyJAM8lf9syIQIEw35Av2qPRUtaeUNsjV
xUOm5zAXNqSOn5VBpsUqBOX8d0VHAtjTWeZkkSwEFrxyyUbQDZsZl0fgaVvNydgV2uUNbsZqxJca
Pmh2R8b1O37Wt+HjFyYUnBmfPfmczewlZlDwT4hCNuqJavu3YDO05+zOlCiGtczSxCjxwBiw6aod
TVihMSN/irIjwI+NTwJwS6wdlY0oBN3/6Xjntsk+sIGl1IzVX8NfwMoIrL2mC8PjaLjJs6crUXTV
KNQmIVSGuE1p+fN2v6CwdLkm/qS2Hlc+s/mGPLHtYiWrKzemczXO5LHmaewTrYjFyc1uF6lwRDSI
xbZAe0w2M1NcNag/l1aS2EKOPk+rj3QpztdOz6Hkr7cAsDOyiVN5mJ+u+mdbR7tWkqfZwd7zMTBp
rAd7BtU4aHRZBAFOZN2x7iTNwjiJ44XdsWVi6Lw+E2i8jKfx8LafyRWuejnARmHq8hJSBNYpWSm+
BXCnQ6YpjxiodIun0lPXm7zC+oW04bjV+xM60BLg+IsfUidPvHKb5LhlNWgD2RW9s1luAiQ2mLK2
Ymph+PvUWfzrz/n2XP1vKF8BbMuSNgdJ6X8Ck96O8czncfUoUrA5HPM/y1On2DUYbAmxXmGaHDoZ
3UhzESGBgLoM9UYKWtntEVfGDMlcqOFXvPWL7TEb3RQVk1fSdw+Kuvn5odJE1tafv8Xkhvj6vK3z
WyUgEEUm5y3qH029gq1yaXdXW8/UVhjFErk/1MUT/6VzhUAZOD+/5qbSKULajL0LiuJ/QHE8l4Ng
kQs9aARcLSIarptqu1MY4HNkuv6W+C9MhxgvnsHoGXq9MVmOVaidvHHThoJjSU4xZvvA098bodj0
CR0WG2bEn3C+R1+pTOfaTkVJwFVCZJjAhgxTUcdIpBtvoRkDVUBSXRkCT/LAU6bQxnvun0z9Wpo/
qM2AmS8kyGYkGgCOEet1gx59KTUo5SeT/wPnXRz38E/3FoiQ/TFtdAJCcfg/NgPBIEelX9PsAXV3
FB8dZS5NOyzCekW0tSjxfG0HPQ+Fs5X+i3xdN7TfXSXCuo4emkCJ3csigvIKoy9By7EHYYOT52xW
LeFuuJ7V/UsfznA9HOqRo0ozhchnWiszGYYkLAOALNcmPogMSGcuBolELnyVQRIauA3ic9/sE5VP
uFte7hJfF3mjV6SeEG+XglJnBO+q4EZDQxMyEqPeT+485b8A8IYl3cuIwMsCSm7FI75QMSY0+wXI
Qq7Hy1LAHxqAiwChqHnyy32XUUW/shFBUGOXF9MrTfXLEgwUQOwrRRZvSVp2SI2xyASWFxaR5Zph
ApiXU6nybrE1+s+0nUtT2JfXKu5NQGsvuS1TU3+JJzs+p99SKJYoiDirMF84MjqCZxbHbeJwmcNG
AGgncU3M7lUY7WepAtcU9fHJ1U7j38XrhAbaTS5d5p9Qc7ZQqz3Gqv/TkYNj6OIRDCqLmaGglgVG
2vlh8btukYIqQCKB6KlxSabySNtrFbtAQ8N3wEcPaxdlMx1YAtYF7Ednrfcs7X4j3ovPo7mrfpQj
KJ6qvmP+O50EP8TWUfOCrvXsa3wwn/VARXtileXayedPncheEkPhKm6wppC+dM0sYebPG+rhLjqL
j+MK4+KI/MJfOGOpSQQ3HE6Zlbn5ebuMQeCpbfanXSX2LpMJM4VI/cHWO9fLkGeuEzHnspFeokrR
eDy2NuxlStgbB0JnlJdw+4tlCytccPpVgIu5UE51e4X9F7PkdFj2AZ0EXFCvnhMTtW4zId2/nQjb
N2Ps4Ii1TVGjsQL7jMHIIVB6Efm0eX0uwxDUBjPtTNLvhU9JQfvwIqI8BOTP8leSNy/FDTV1ZH7m
Upba8Am94couSGFzfuGjEVkRJbOTmv0zVilDNxKK+3XqFEqQuXbZWT0H5LdshofiA80Ab1qDEpkF
RiUeZ4ZkzhtZvOpDWZSHxKY2Vgc8LTh4AZcDTtQQY5bpEiFTAYSpU1eqeji8R/4tHY0aqwo7r4lF
f/RgSCdvklCG73PH22IDg+8Rns8zvo8EccUGarHkkkH4Wj4wgWIYlFQvN7a5NAZFEzjVNNruFhKu
zEIYB/SX+cITXJ9snFe/JQ9IZ8GH0KieDa9ZDXJo1pCcx3uzPN3ipfVZ1EhdN40U7NH+wIAP61nR
3rEXuEJBXIoAaU/RpjeOBckXk8a1y4OqQwCE+9wWdaTmOKBZWCmzuNdHmbOSDA/3lD+3eBwFfm05
fbZke6w+GBsrDZOtc5cdnxuQOfu2MXQYYV5Hz4DzSlhp//NhjeWeCnrSaAEeJYRWh6sQxusbVf+L
OqlKYTVM8Hwd7oT0CLZXuNfRMi56HKPUf78HgOxXfNCHfW5A4v9P0VP8GjTRSkHYIod3PyzAqvZz
5sNdf8BuNChOQ36o6OV8qbt0Ux2CuHadKhAZedNiIMq4GauKS8k++8qdV8oLdMShVEUqOjE8rukY
5tkrpjJznZ129l1IGmV0C1YHVxwKYhCrBAUF2o01dbw5RbgaH9I//YXSJY+FJXo5dJ9PUCp0s9l2
aEmqBti4dQvZYVJogfAWGBBuc3DUFYT0E0NsIenb598evYDLYV0k6bqIIViRN43iwbDsZIZ/Qkjz
w47IPBZlsGptbL8m+tZLdhiqvnKNFfR7uWkjfa7on6OtWenKXSdUwYOLOGjJFmVNVAE0guWrAxUO
Ya2SaO4Y6l74y64CvG8z84DeZ1NwWy9bnHHbJs+AneJHjvss0t36vDhrsvaix+CZxyu95+PmX2Cf
ez8lBO+JP8ojN5j8H99EL2+bgexy79tLegHmWRUJ0kNB/1SJBJGBKpZlILKxuiiyeR6Lp+Wny8AI
TdU3nd5gT7tiIJb1ayvWXaUoQYfmldOuw7e1UYlDVTGq1agCYy0tbxBr+vdFdDsWnWtgY813W6Mj
rnTYAIJuQOVgQW96ARTslm+BRqw5bbwU1f7SRfuNt1UyKY35mkaLHKUSpkk7rXWJevDowZp5xzD5
b0asaQ8XomL3kWsn4HsceguFE8jvJgkTK3a1Qewhz40wQEWid6SGafv3dQg+LC0bWEqUzRqJ1ahm
zCZ9DwxmRsivlpwyg2UEtKkTjMvyQJDnFCtoCeMxzYhXzFw9qJHWuyhYkDeIpatuUDJSo1XyQ+ST
sMNh6VArSqD4WNjbiUga6ERXs+twCzGBQBnneHnjyBQWZYIpt6D/BAdgxhupFZFfF2quNZ7I2xxf
2P7AfcUMoJ8wOcqcT6HH91wEQSF2siMzJNwss2pXkAzZ41beea3Sffgfs1RK7dCuE8zQAELsA04l
r0ASFd9RJXGTbdNncYOAPIvVLgsucKHX6PuvVEP0meNn+yX+a6Jl9Vi7pAdxkRIS1Z2Qjuiff+0E
6AkMAgqBuXMavC2ozSX3RVbJY+ZcQYF6B/itOCZw6lP+vD5ykka1QuqCnIy3kHOX2djAsb+g07q/
eceHOIxw6/cENBlfYtap8NiEHMpd7DDE7/UVAWiKHqnJMDGaBwhbf74wJLfRt/YU1D4MqWfXa90k
eLowxt9Upi64FygHA1oQ0Fu9EAGqeiNYPkeiF6GaW4BYRMwfuN8ZwDAsa1M8fYK2ZraBJSGyGG//
CJ35ULwuFcuKFLqaU4Q15fk562tT2Hqez5WJD1BrobAMVYY37h6SUTNCO4L3U83tB4uBD+glan+E
MrrNn+/gZRE43HqyIc5VxyAvhW5yLxOHaH/opHtk0Nvofrx3dwONlv5puHcL/JYvnBwZ8PI/Nj4G
bn2wJOlS/ruuSDG0cLXFU/q2nGxRK2LfHzsG20SMq0QrWgswxAjgcbnWe5TcHLCXA/4JC8nZX68f
X33Zn4XyCo6sFcbzJXekaEsJPruq0D71ah6HNhZO164X+1d9k+CyVMt8OsspTbzlVRp3AjmARU7s
LzyG+EsJYjEQ/xKzE2Y5AWmdfd1I07N7/vh1auGR2RaWxOJJs6AytphuuK8tdPDE96DvtrqxVQnv
/WpIhcUe5xe1WUCXfdcHOxymmXwXZaWLbRIwxnQSfNqOSJulUKytBa43v7Y0ia0CXoPKgRJfVDFj
fH3MF/szW3j+Xr/97RzH9ROhYKzr9fGe2fOOlQ+RcTPgSRwIx+eC1AzPjVwc3hoxumknW6Xjh8qb
zOmh6OR+g6+s01x+1jSeMEQRwqjdAmnfR5pZW7C1FU2zaebjUJB5Bg5yTyqB40Rq/osBiEnJk8Ca
/JEPy/l4CkDsQmzSDCkQUgY/ObtR2kpH8zyIvMTe5oboApQKH28QTcU+66vfCD7/2Dx4vguY7914
lcbe/nfhohb7hwt/9rHTOMto1FrEg95mWIt7wFvQH6Azxn1NSLJQ3XU24UbaWC6fDCQGChxPZQcb
KU6VHB4Gz1HdF6fsH2Cz8i5v6v5dMvcTpp8dp8FyVkTAYwDCrkdgg0T55tDqmzCnwQGUEtHC96PW
2VKaC0BGOjziIZODHSiWLxvF37wgRkUcPNGvScZ/D4i8Z35LnqtJ6H8gTvvJJAmiKS1CdrzyWH+h
+vcg8gb5mOXBB4M+RtCbqbriXU+3MtC+SwtiFK5zoWBa9QvGwt/qF8Rx4PoeGfpJRvXnCAuKc99H
64/0YtLv3Og7q2Snkt298pHacSW7iM3WzhkabdsioRAJPuqsMkG+BO6qReCNBquPsg9zRRAouMdt
RNEzxVRcInZmUTydcLIlnyoIXFeMIbzeRr2hC3i45m8bjt0xNshMfRw68051CzpVrHTIWvsdNM6r
mfpSKQCzoPPzepj3Ln78FY4Cn4dEQT4cmX28gN00n01Drb6cXpgmo7uCbkFVdM7cOjlPfy/YuJ88
KV58FSiJHVAgDU+fGKX/ot41djsmqYO/Ub4PG8JPUNCBENE82fVDDWh1sUqVgVoh6HLvds+auR5u
njKV1cnghCCIU00orVlXwtBMYXkKtPZ76mTi2KdRsDSp1o3lUET+PgoxKmzKIc6zsJYrdkYziBWe
XGSOcFpv1P+Y2kMX78bUKCL+PpBRqDqVNkaFwOtTax8do06r1gAsqGNXZf6yFxlMhqw6Bqwas6+n
wv8a81YE1d8292WeFjDi/QocGk0UQhUual4AbNn153TFRoxS35cIDEPCoBosHX+NpbuLxYn688uL
OLUpOw7oicl5WaKwPAUcy3ZDD99B+4pOEmbD6u3qfPwpWbplal+YFPvuiXmju+czOdW2Tm7gH2+a
VxXllPctABC0DpgaODGYF3ZeQVrPd9/+OWZo88/6CIjZbeWRJvRyA18S7rBJtg6jqMD33yHQgoJr
3m+amvIcTkDJYHaeFYnuwGtVPH735RwDgJsk/dWdU8IsBWej10rd1Yhs6P26PyHRHCTi2rNeWf11
njHFSt6h48V4V5muXSffMy/G6D9WiqBAtf0xCApYHZ479S8HiXL8YXTcpCrccJo1sBkUpxUfSsOb
dfTBEYxQn2mDTCBi6Kuuu2oKeozFTqcnrbGUdDrP+RAGYBbPz0HJuZSpco8/j7q1OTzpkYu5apVM
uSM0Mn9DD6/S6zGo44dYTOmBVtBSNRXH6ojMiw8PgR0/+eF9IXHIJqWGDesJPfAP+tjg1as4SBCJ
p1bpZo5DpOXMUSPmNnEeRQX71r2a7o0XHpbne1CrkOkFLNxb/8LPipHnr4MMc5ERkrkToBCXQ0nl
MTQ9ndX2L+h5DthkTuaK2Pm3Jtv7NzIO2xiNvVMfVBfpY6SfUQn9xOIjgPT2Y7nentK8BowW+qiE
S8PC2BybbygEjagzJE2p7pbu7l+3z8KLg09k+m+2esDNQy5K9/Lsd8uaQzL7bkO3Op2GtloayL3U
b3+gqP+I2DtyFoReyK6jbUkrlym7ep+/Yo5n5Ru7tO8qw71mh+5AgqM+U+LQHNPbJ6URAPAPMb6d
86Jeljvi5eVjBCH8i90Ze3nKwMvnF3JKp4oP+ZcLxW9acNmXEz6k4hdbnuAWrYtSFF1qdJ0C0e+W
ySu6cy7PsQQAUBVehPhml1vvdKu34sWHNm5sbsG64ytUJhUk+J0vNGwiBB2IsCT2b7OPenEgwpGB
6UBadOd51VkxduRsj4dh2kLWR0tEYQs1df0LaAz7GCuqtYsnX1TI2PxvcmjTL3R0NBwXXRRy+gxm
kPr/jLZ9gElZ5lEXEaCEsiNCAHQNsJ3bG1l/gIbyDN9kBGwpUSiRCtvW7E/NUCAjDewXASDEmdJv
RkpdSDKeQ3vYoGjwWfA/P6QBtjTT3zvU2TpfDsgkbUtVdokeRHMdBcODE/oYlAodGkDEixEHNY0h
O1fnFiItz3wlB2eavJ5TViK8Boc7FB7kXshD0SZXunUrEGe7nxVeEvB+of/blvzOJa+TCszNtGWL
3Ix7QLRxVGHesfpbYywXpmaEtWM7P2mXs/+A+vRt46Gq/j2hU0zRqf5rI1J8i0xgl8QxHf5Ofn2J
2bfL0SpnjZKgpjd1RCJvMcg251p1aS+GpQOjC6wpv9Lw0CofwL2q3kVMIbXqWHIvT5zW+xFnQNAd
5YKzs8sRIFGGwq9MGOcCBFtgQX9bfiHKdUj4tZcqDQdkWMkWvGNBZcbV43Sb9ucGch1R9nST2Ety
CM7rgz4UYTBb1iw75scRPuOoaA00D9jny86lAsnfN//pXAXEbe/uEXGTAw4bp1bVp2OH4Cksw3TE
Zsba4tmoUICHHRdVJxcA1P/FGd/SEdWiSijwkSbMNn1FXypJ0vyt8J0A7netZbY2TSwhnKS4Yutu
bjvRKpcfkZxZzmL29nGC74mfsfda2jKRWOfyjYcT0x1XLPpgsc27+Sk5gn1c3jl6ZZhXg/NT1xy6
xn1nw1s8SMRBxG/lYY1CH8+xnLmDcOrW4KvbF2xrOtkZkBUJZNfP353MrgSR0ao9Gql7umkpHJJo
xt4IPINbD0ofRp7ixUZnWJ8dYsX392iRbWXInCBIEu/oTzPKzFV0Ulv2VHIayeazNq5KhTk8HYka
YV1XJgCnf/cJxJMQ1P8nni7tVAg63Q5/OVe1vNFR6vQFwIfdEWmfl2OmG18ueOYlMuNQKmixYb1M
ZiLfNLF89c6JykzYCdpgpY7t1wX9yx8spTFt7X/UiGgxkW3G0WLFk6/O0gnOgiavCzW1w6CgdWI6
wRKcyIcSCYUiqYQt57xvFMcxkln2KpBkWvVhBbadXlqXXtHknGGIFX7qCRK8PsvxCy4XtMdR9WCU
VZjZByEH51G28yUh5O2VI0dkANcQiYBuqkuc3xPR7tVHZ/hOuViKj4kdE1r+3gkJROffB5gy4viC
MMdaQiF6vkj96puVYhtgcKO9w5KHKfa6qfJbW9eZ/kEwwT7gDFdCH9VRfbJi3dHjx6i0cDGl08kA
sxY6HPA0Un+tYaFiBPm3pvvHxM1PRVj49vsOIS3sJeHF+QoYPBzjNZ8VmNdeCuG/LhdjFU/w+EKH
GGASmnVGWkxCjCDUmSg/BMLukI2MsOuAhiD/Cavz9W7G6lDfv49Jb5Q4HXFpgNfAu5Enq0QRIrcI
dRvSggB41Rxoqm7+tKBvLDmNK6kjOjOm87LalhmEctdKAk/vhUgu65ijtZ5TWMFebSVZ1xmOWaDe
wlbKyMqxtgLh+SEp5fjiZa7SvV8Z+9d684jFd4ZB6b/Vj4p8XjK75gH0ukBNYA0y+AfDgMjO6IxV
nBuHQSEOSMEvprsW0AnEkAB3+oHiNokI9aiKxvyEIKMaImsc7NHQeE534c/M+/fkv9aT1CU044PD
2gI3lEgcOavvo0cDGYynz2zEi9UWDpWfguzgxUt/i69c2myZB3bPffF3w5gszVwmzOzDDn13/25y
b+FfO4T0wWfm22BHzYeQkUBPF4hyK7ghV4OPVdjngGW+zxEh20gSze16eL1EsD+TZLoEvNGadJGj
bVD/B+LP+STh0NRHb1x+KtMdRzCMAjtckILVkTMcEoV58G9JVYUBlCkCPiO7xcV4OntNHi0E5/1x
ZqOVSE7p+6Thd3ewOPcJHwWyCtQYkEdjKu9iOZ+k2ydcO7tsQLcjlq9FOOSNtC33YDpSU/FzLksk
dBI/7Y+6zgnwX5w0y04FKSPbrCOQpim715wgAEYxgRT80M69Q44XPMQyOphpyN04W50ocVD7Gai0
bs4DyMGl574RaXjJm8ggNQlEQcthovB8Eyax9UajFoW/smMj8kKfoTn2RJYGGozoo9eEZhdk47ez
ZTseSDZwp9/lQIqN/rixGm8RxIAMB4swLgzaed1ntRCue/KF+c1X484PYO9+jjKLfx56L+vl9qFI
Y1/lkVDvW9tHj3fTbL53mWX0coR1I6TKeihh5Yr9ke14DMv5Y57j8AbDB5o4KTpaxnBveDPz7WdM
rRZXLEX7E5ScXf0zM+CDcAMydDEUi8MbxAFcz6XIlTlglpb9FiBzbLs5B5gZRSZOPfut7JCoAHsg
zbhZNxwGKV+oU4HhPiPgktmz9KTT3dPvTJL13ot9qPQFSWoAIVkVxAFARG5u4pDSFeM5BY1eYh9z
Zaxq8fepq3A2/dRwxCXB2SVXn0lScqngslk/hCnwRnsGNSwTQMNyRRT19VT+uTUOYoInWPl55YnJ
zJrBzyuuo6JQkfFt/OC5k9aBgcN3dLbyygFhLBTmunVWwA5VVkzhDsohVygHESXBBOcY4DMVNG4c
+b7zZuNT2opEt26pCHC1NJdXDVYw0JqKPgpftb565BOv8cTLdF678p+ZPvcsWiO9UhV41/XMOq43
6PS4ysSjBoHjaXBNfYOwkk+Qi1pDVTrdLjsSk4W7XtrPLWFrWF4Ix2EbXd2VEize5Sq6NA+Oq0w4
kGKmXFf8/zu8omGfq4X/EgELYjFeZkuu/HiZBdKLUlcrV3nuXSf+4Qe4IW6a3NvZu5RnWiv6orMG
rnqCpGm82cCSAtVoqW8jFSBIDc3A7OXU9bh3u6X8WulnSCNrG5tfI20wFxsemXjqaoTqlTdbuCwV
DMpO/vl/tQpQZl2xAlXID0gNdIb3ifD2vLzAUjSgRHVRn2cCO0Y5vACw3B4bum7LYcXyxbdAfmoq
hP57TFEeCsSssB9cIUs9QUU4wsNqdeo+XrjUAyt6+Ddj2QLH3It2bsYLVIsAG1h0lLZyN/ovzbDp
X1KBLl2s6oEleU2MmGeDJAgtOlqjDb4k8oubwd104FVXO7P2tKuFA9eQMXvlu2bCLBQWB44WhhgF
gySKU4rivwf8p61EjsJGQSI/Qeqed+40M8fK2cY8xskshaWx3F2DvlkXy+VTKnWNfRBnLiY7bzgn
7Kzctbk+NFVf3sWNmJB4UuCYTy2Vi7muXZYTn5xwij7CTvR/R/xXKgPnTYdoHZo+EZe+qSglA5Ex
JBn4PK8+JzBRj8pFDzVoCn/olHfwMwuJ4IfBqNYxmiGYWk26X5kETY9wqIdAX8GVU4UQwyogWdnC
6KUzULJpUSVMx/y8Qr72OJV5BiaIp4KfIQGaIR1DLVM9VHY6K27KCYOYIvr/R25zezzu8+y+M+wN
VPrwNF+4ydmhD+SRjPYNjPos9MVavdsAVZJeSdBKKasipT+2INZvXoCifIkbP5IjRyK365cex7mO
ZcTUt8Vgayiyh9BlcUK8ZzT8nWSUfRf7KFGysP8GRjzBGPc4wGc6JJ9nHsmg6sUKra7htAa0y6Ij
Gy1+V2coYDcg65LN7xHPQeygwXyAZ/uq1G6T8Kv+1dqkFhYgSAI0yFYHk8IdPnEF+xixMto3enUx
oakLhLPR+0LuMspTPyGf5lEc/NzxpgF4Jg7cIOYRmsf7MivS4jrNHkBWFo+aUhHqWCJoPQhnxZ1L
9XMsss1kUkMAxIz3cXSnd5/ZBkwdmoNaEY3avgslLatwePU0nPosMW40elxfQ66dredA9UplFo9F
fGR1xvGo+kbwjTa/GVXimE05IThW5QxKG43XRf9V8LJhMtg2caij7mJxf5fs2cvV393drS/SNV8B
sO40NswTJU1rWKQ9n0Gj/2kgBNkGtmIiP27JJwpNoFkivmYjhrptmdiyjU9xLtR0aXuB32GNRNMP
FZs9JLCBCMKkiR4yPEul6SGR4aY3H5ESeb+Toqofio6oFMyWAabV4px2sK6KoxGy9dtOW4awrRs+
o6aNmZldhb6suJIw1A2Ks8LIgZcHHIxLK+Rpx9kIcRW4UuZBJaCpO1cEfL7quPdeqMaJ19r7nHDp
8BDgOaA36b9LY6P8hM9KKNDFSaNrWP1T4Hdk2C4sv7mXgJ5A7ZLi8E+gL5v9Tc92VZydPy08D9Zs
nQsDMqkRp6fmaXv0BNhjP47I79GuUyLVanZin3aXEvCa/OSkdINn9qIgp5reEVhvChP3jeX0+GZA
SGAlU6kr9Kz3OKXZ71wwiJ6sGA99UrnR2wAUvY4W+29arjYvfvdjnQjspcg0TX4+ZpIqkgQYwIUU
TSTIBRVBZIc3tHf7CpqPd+wHmKizq/3/GKIPDn9WIqx8cjpM2XN6PYEWhTfs6ae77O/qnGcMK42P
pHYGRDhL3rL+GnnY88ntanw9vjZ2+H6p/7IXxFtMgCOPkgS+MypKUIiR0xCkYiNeHeZ/za6aiQVS
xrh+GmjX8ZVX5VwuNhRxRV0pg73MOEyFujWUxTkBvvw98RdWmfolibGxDj+oejkWWOX3kFEThOal
hr/FNZ1ZK98r6TqjLhAHJI1Ez5JAm4Pgj2sroS95TCQLHTWx8Rcq9KAXg3X5IrXe5fFE9wqBVKc+
tbw8P/Hdc4dxwNs9hxkO1RuEqM/7rJf1qrvCytQzj4xvkMMBXMRQ/C5fD06CCW4ySqgcYG4fgIhH
HWk+LDw1yGSFlj85Opwr0bbqSmQa4GlD+qIhhf/vYIr8zK9SE8fB6jO7TGCWXLJmdaqCiBKFrqj6
iaJloPJJPWzQj95mqUj918uCTscpVyTTluZ7PtIZkYfWVJxGR7a+3NuWDGAh0WIyeiaEj9w7hU/S
o8FDyUdk8dUs15O3B8FoL5jjBEEwz8K+d40zAmaTNlbpHcPv1S45ai/5zVUXb42qPpTHrEFpERu/
oFmuIie8rjQqfHlA6RVgCCWeHc/uiWeMRHStvowLRKPO3AJtL9pRlncpTDiwghv8s+Egc20B30b4
ZKJh96zaxdmsABFBGB9Q/a6nXiiunTXE0hFdwP8zOhBWYzOg5bCl+K8VPSaH74Igt2dMRkBLR7r0
XlHh2U7J1v9dpnnRAI8wn9qCQv6dYSLERqfjhTXAJEe34hdYRJLUMglWfc1FMwoMbZ48brSYyrwg
DeVFIzuc4W76BPlHBrqcQeQq/hpCKqH1dJnVtRCTf0GI946dTnrx1n4H6wb8WasesSwPv2sATAKP
QGYeNn2FqFZeZnmwEdyBPzQQbDUHk42DTlpWbZ1AEELE0kO75L/K4Rwdfq2tvl5bUPIEeB2zEEgd
SCIsgc7h9gRTMnTerbUaT2o7seViQdPtpI82KdignqgPGa6ZpELsf0NXLZLq6LwYb56RGsjjo7cy
pR565EU9THQldmEGtmcnW9LN6di4MMtEEoUCILD+0sVG4kLW5YL+tLW9SvEGOGHO/oiWQ8F+mOBo
eVsIq4qfwiT3tBSfJeLH5ZsW/1YCwWeBLo+z9FTqJeB1GR90g2LJ67LT4ZrXVcQyZLXljq1yz7ds
3IUnoAyahf8aVHJxPenm8LNeAK7gkEm/+XM2I/b8791IC0KeIjnkqZGfcWjEwV10W7JWVMtGNViO
XD4Qx9Ho2Ls6d5IbGg5Xgbr5gLV/O0i4JRs8/dW715J72nSiC6VRJtVCzBqLdzlgFVihZRMkqGfV
xYf/Gv2QmgEhfuGPQkTTnQVYFmSwqtyB6hgyUuKUrpWpKywfym9CWSZkSLzMY19OSr/T0pBOLH0Q
lMvu9p3UvCBZQTGhpny4O57v/Z6uKhmCwRr9h3woeKCxxVmaU/C8ny297fqQfV9m/CgMUWheT1iT
dhRVO126ZTuZzgcBqXjLtREhgnhmrbNNIehvmV8I5rmoGNTUgDWEosCyqJkqZE+Awsy04vmt+81B
PqM7g1gT3DY1kt353u7sJdXqssamk+yqhrh5UH3+cVd5Ac6s4jc6DSVioFff8oDReO/gBQWsmfKf
fbltswEuBxZmZgw41Qd5GrniTDmwa743/x/YLzHgbGlX1jpzm4F6YmEzp1K4VHaybem19j7Jjye7
e97HEHg28nceFRTq+lHRmA+DfVu0qgNNdM29jSPsF95C7r2jEbLhicg3iP8+65+oeLgzyhlgf8Y4
Jmd0hDZWQcNrSdYvv4iXX428tVmOs9Or1xq2pqeLXtCcHAhYyq594kS/hqla02vbsIZH0FAVKypW
uV9cEeqZJxAUCJ2A0RPzWBcOpWk9GPIQQFqbscex7OZR+tdBaxycCRDIgAThZxTmLPobBgBm7qWJ
cDDOgZOniz7UUEdk2uzhJ8kTeWvAexT9XT57YvC3HfplsFC7uO3UI95NS9GC71qq258xxsAD0pkJ
dS+MphFdeVeC4jNpHzlSST4nPq8IYoJSaMKh4bgev42W2Uomw/1fXYg7IOiRLoXTb0lGVG2qgXOn
ysWx2tH//Yr9l010IE1/sPDEwnnLTAU/oequG/rGulo4t3Y6h0ZpnlWMt64nz+Hv2++Loe99+OWd
RfRVglgIxTjj94fno73pAxWV5BycOlubP6CWmlYqg3o4Y2eypQjft3yiBUqLSlNhrMzudaNSlFkW
0Rlav3NhG7qkwB9EhJo4P5qnZt3n4Xkzsqw8sdo9Yb+4P9OjG4aONOOKxRQNoWZw6/B3GGL3gDA7
09LFFEXG25jYGTiNQtZUENj/lfyO7m6DxNehMJVm1TSDSdi8IEuzBggGohWUqBF0ynNR1yQs28Qu
rg4gINO2fpfFCvLiwBBBw+9E03SZbUTJ4TznAOIz7Mn2mI3hoZbNAFYrX9DlDBNiI6+MzQHybPWJ
39jQ5bWoucB+E4EKzNG5spMDdg2xAW8yWBYt2+05n41ohnZCfNGK63ZtQ+FI+OhdlKyIoMoMJ24M
p/rCoRUiC/n2/UX5ABNvyYXoQwyVx/K99KramYoloLKb0sFD2W2ZBG+7ptULUTr/NOsSxBc/IP+M
BlffAFqrOUygwVTVeakITdT6mbjYYFflMsq9iqmAyLvb8QF1z36XVbiYMOKrlfwywxpupYd04lcd
AC8GQAydLto6gwWHLxKRStsf/pIUY91yzC0kSZcVOMzWaYNvzlTHNFd3rd2/E5GzcZRj1IJSqGwm
WXvYS088i5lqPpEGv5vi95N9EqCAEz2U/qXnKW8SDz1LEbe04rXzrc3VWf55gN2bC+CVZkCAEERe
NeBkMvQpKxtBZhjQ+OoKwpYDwekwxWxaSYUygqyduZkdCAMS2ec+TrtQygTETXQ1+rZ7+ons9tgG
4PVVMi9er2bJ+KKxlabXPqrQ/+SycHUY8PnDW7Ge4UIJImbp8GRTzeH4+4yHuUiVfaBKA3+5Ug24
Sb2E1wR0C+K0Y5GX6hKD0P/357W63QH4iuzW16wqQMDg2dmIvn3IUVG8X3gObRcD/kzDvl4OmpZf
TEofhPMOB56r3/vUPDfP6ENMGBxfS7nwwwzw0NZzzck/erYJ3Z9J7I2BsIpyCVsy/nTjEai9gaRG
0bumPiS/ksHd0fKxBJsfSAq1T+lZoPIXy97ToSQZkpZOdJfVlq3nmlk60Yd6Tzb4su2ceaoqWg3n
DXQNKBE46O0kIpQs/bZZsteY5WSG0CKM86WXG+FCNfWyKXbLR8dlZxBRsgOYILO3gBFJnOP07K0D
UmZzVlXfHrxTX5aJ/R0D2o2pAPrhrUdPyU7crMi+ulTlkWsDPKaue+vsuQGFaOK4QB2SUTrTRxta
O6Ks7KHh66wDdQ7XsmsKVRYJ5pa7h6RLn4bV5h4dbsIW0RgiwftIrUzv3YnKjGr26lBiRfvt2Xrz
X5Am0wDKOGnX4W9SPg1jhvoJ9A/5HvTWRbOsQ8ApsJdgICipx9xWrUTn1dJZqN/J4P/3rqOGdw6c
44uhA7w/CErIQYHLNkQWY4O7mpzsEcW97iYL16AF1bPQ8grO1Dh8VsNUZkL1YAx33f9Z6+EN0700
aNIp+MPqlr9dFBIXHDD+v5iYro4XCZApnQ5jhwd1IABqkjIrpN7E+J5HDk/uiYZHvHe7JhyDxE0B
VdYUm9wTTX2rZj+KCwBwOOSGawCwoRiG7sp2yS11igu6sfwfjmumPKIy1b2gahj/PLqDksXNM7lU
RJqweVHzEw5JNMgi3CPaJQ8nmGa11TNFfmU4lPkZxdJ0EO/bS+ufNGlZkWbUCTyO6X3whmI+nslH
VjYl3MCDyQhfWQ2Wl3WcH3Tymtkj91P8vISAMkmCOySmssjnuO12AuNvGcExVgajGU9MiSbGoesy
FXiEipVf518idjUUAw/EXrC3gKRiU6CeARab34+GSw18huU3a/xbOooSvoQPYecXRai8ZZ+cW6DR
mgOu6Q8SlCf86cVyWNLGfKfmb/JRBEazHeKtf/HvZ3ircXR2/ScOzHXyBna7RR+2vDIK31r7KLEe
/fSfUtx25NChhCShYb6ylNUZMKetYw+PAgr1FrujjM9d9tJ216JwETsii/rfcZcv3WDRe4H90Sro
67tz59CkSgfdM1dP0kX9pyBnlyRtJPhzmy+Vvd4gx5LAv6Y+eNDzWk15hQBKqybvRWPXj2yOtFAG
zOozYBafulaZhvDI8G4UGQWRjUty0YW6Xc19gsh4ifv/f7/YXzm/bAvaXYNKZe1gAR5t+AmQtWoK
XLckPHUrqDIS06lsrvf0EUh7AoKc6FmmIGPHyLrwPQBbUMXx/nnJTmTywgibVvECYd44M/+HOhEe
FrADzcQNQlPQ4IsGXd2unSgtk7FfHvo/UwYeDziqja8haL6eFbyCnfiRNCL1JK44uPVLNbtdZdZ0
A+f4xD7YaD5eMpXI20b9IR+Lb6CrA+RcnebyT+KUGCOnYNFPSwANdCIidAMXXtA1HdNTkEgxP517
ijfEzqU9s7TsEHPRvMhvj7sA4cm7rdn14iTJn3Sn3Y1fYvxac+oNxW/8M6KMcJqe63xncm2qPbYH
zGU89gZq7YXBylSsiioVoxokJVD0a0OExXo37e4EhGFJVewS3tecoT5bKev+10Vz399olGThkLXd
wPPO5kHSP4qn69+IhsmQ3rXFN8zSzE6Z/7f9RU1wcwkUyPGaCRvfmAqA5gkMHBP9mEbRgMbSYa3i
v6BMyYMb7yw97LDUKe6ZaZB83x5vvnrtI80EYkXPfDuSIthXoCj/lhSatBxXDtbx/PqNrnRr0heL
+Nnk2Zg9yiK+tYNm5lbUOEnXvIyfx9hp/uoJTPbswv1WzCx8QdalA2tMb/1RdYhIRQyi/zlDlWOj
QlOFXW0tk7JxzHLMHHhbLsaSEhJ7vz+T1h7v5eqvpbm1NTbS1PfPA0mxcmEYwq0iNsT40vOCu6Nm
vrj+K8ODm1HlN6XDceUvulR3DWRHRDsscHt/5qrlPIveO1yYSS8jJ+tsuKPDtbBCWwg7crS/RBK1
lVXxAMxAcycliI9JnpFsscKvxSP0efM2iJBFDfxJCIsAeW9ccp/xnPHQ09ld0cFLlseN1Bqjqfzx
nHz2Q/OatMKNl1Dd9FGGkT8pGN2Zag/nOej/sLDQioZAzmcXJjut4rC33vy4wn2JtUHp7q41tLPN
euLQBp2cxF6XIKUcwRf8ZPKoFGwEp8H61XO8/UNIZg8ykn+iVAEbUJlwud2gzUH65DvkHonHJDl7
bzIi+iKuzi1oNg4fsKFBPvdY4JN2Qtv9yQ9E0N/0ix361dWPD82xiWot+5h9j/HUg6XHMF5++qbB
Xhk9Ym79/Kk6hcE1ArL+etcyH9ToytpDAZS0Hgj3wa5vtJZZAqHb32Mtas42qt6T7P45NFv5nimM
+XdPcyo6LRr8bwi46JleuSBcD8NqeDT5lhoIhvKi6fkMIc6njU+5spBmeKqArXqvovKN/Bm/e435
nqbQDXSodwtg/cDG8al8fU7c77L5Me2hZl965xMZNgAzLSlkLXTIyKsgIjBJCixzSshDF7kqwBIZ
V3a/sfr95Xmw5sBm4C30rBFasnUsEOtvdAcJj0lQocbnbol2QmZqr/S4cczbrEnhnos+ePGnxCNQ
ZTMjsHJ+ZAiXiUlh0kBMMvVRs5pwdqRO42ZeRfhk9dCBaFWjDLK4mKjQYMafl17pvnacRpoM5QRZ
0F52iG0qJlC/6nqzny6UOZVwOqqzwlVhQcmS83XZ46VmniDbtrgRAhgdHE8B81W68TbVH8Xv+T1e
rTDTTeIqP+B8scbxoS+8AGAAWpQkGRbf1wN4m6Lt9Pcyq8gGrjYoIOcjDmI5dZg5d3JVsKty/995
zP+iA+o+vZsjTHr5eNgX1dtu8458xVfUM0WJKViH/ObTStDzZbpa+LnuPh7vevqaPJDtAttPKUUc
R5HZ5v0PDUxHxLKz3zOwbGRkCiwDRL9rEf9K1du9cOE5Ac+8/MvjZhJtQuWStohGJVtqwA9rddVr
g0eQBkE9qLQT3X/ZXka3tp/rwO3ZjyZT7meUreFJFFRKwDZTwX/pe4scc/oj73Qv0fWoi3Ei9diF
seBPe2R6rVQd0EmQr0euVdM4BUnMY5IysJacvwHZAAprdR0KTgnMCY1PAisrprtZEEdNF27F0e/T
BMC4cZmE6GWPhSueltsUTCSUsKqDQguE4/Np3POnaSgDL6Zy2/umem1CDz1B9Ss15w6XH5zqaoIQ
MjuCnDjqf4EXj5qF9oHlRTr1Ak8mCDQTrDh9qgZ2hRvCAjtjasagrFVYfeafMXGfhg3TNgm4uoyW
RpU1+ZFINZWfxY4IRqqCEe63CLGHonU9gvPdKs53jf/n0jCH24TH9ciGI9Yh/ogfYU8lJmiY/RGE
31B2+2rF7b+CPZ41ly2G1n1FRXrTK61hdOMGk3pBWq0OTmJ7wafc3HWSiEP6Ox86NsVa8EZ76Fx5
SwJ1BbrxIixyspIPcD11xG8cyuVPaRg5bahV1kYk1+bVNx0+4GVzkIovzXHSj2dCOCxSoZQ4q2Ks
e2HCXG/uRZQgShX8A6jSW6Hs/1/48U+OD3QFhqddVvL79DpTSWYESmj9xGsvCEXCOi0uMfKlCg8F
QmjjdkcN1CjyzKodPdwKaM4JYlT72o7hva9mm5NBQdvZk+tPW15lYPaPnban56XPDr/XAXYcDhGb
tbcn9DJmrnZRD7vaIPve8yufuUgQgcUvoLgIfWz4rwwWis1m3tx56NF1wl3jzbbqR2b+ZUXA1Ne9
weR0J3d1BQ3fdYbWGihNxCttG/y47uoYPfZzA/VDNf8vO0Y7OzpyrG4CFyWinyyv6LgWmuhksg4V
Pdyk6z0HaiVOjZ60WhbEt7odQKzdp2WGkK9DgJlVhIRySrMwCZXxmI0IifavmzlRfKqsBbV/7Lzp
anlg3CKeyx77hoFPsWm73WwQQZgzocc1Zp+wbOGXExw76N08EofcrUeRivUjRnaH08DgwbiHyoH8
l8dQ0aTZBYmCquGP5viAP0UQn1Y+2gizbBz9oDCaDzMwb17yA5Rl6RlvqLFN/m4fLfWH1JaGe6Kf
NGraG1fEuYAog7IudFdSM6e29dEmjVUGTv38CJsHMsQsjsg5ufbrLGGiAeTSvq3XpFUEFtl6Uvsc
G5V0GbfiQVqo6YLIqyY8zGe6N16iJ76ptKzs5kFKRXRSodr7edy+NviDlcz6ODFazJgx5ezwUI4h
D5zc49x+ERQS9WsYAHkwhydnb2CnthG/mHhvw06ZJGL9kjYUKQKQ4+jbvNGz1P8/eNWUibYgHNDZ
Yp6F0AsfOcF5oe7SPYwvKRfZL0PKwZCP3rDkXPJ4+X56aGoe9PBslyC1Vim+udOSw2IbKz9bai3a
crYITLcLAlp1zpmnm2XN6CvXoxVn5kqrqECq++UTc5ss3Bnx2n0CX+NY2gu04A46ETy+DxdbIM3B
tm5pt2Mp3fot9qZjXVuA6WeGjEWhha1XGNf5KXUm6ZF5R5mrGMG7r+nUwz+sgm/eDhzXXXqLSr+k
FSMbTZyFHKPZcLGE97SEMdS0lFS9lbepHzzZ6fLokicpw7MNDpfEJWbs3FX+9TbR4V90q+R7lOR1
Tq4PEnw/2G7not8Rha82MAKKSOV2q34dTpOVv25SDx9YmlLmqW/vhFvn+dY/86bFzT3PCjsIl1zt
w83VUUBP+fKebch+JhqKh9/yZIXs7V06zO38sIzZvphLeqLJzplvJ7Aks+ZUxzSi/zT0SSxpYrvZ
jn6vZ9pWYasP6vHuOBezAeJjtqo/H31CDsnTcgOy2sQcOFKdsd7c17setkeqoUq45LfQlU+gPp1I
UPBsgchu0Hz+JzwUQWhuzYqieCnQ55/fopuu0WC3h65KY60v3sMCut8IrcTbcu/bOAON5R9Zo5Ox
uXRHTqvzDr7+6/ig0L/ouJ/V/ypnr11TlKFj4Jl2pYBr53ntZ+OyeVxEl1N20nJ2q4HXi0N4WDJ4
sdYChG0lJwXA7fELsichvBkpLYpcnDk8oUvicALQdeE6yJfyQ5vCn2z1Y3CczPDzCo1kegPow4oa
L4s02Rwk9leaOxOFYgV0tt4gzO3jAsQugeGn5koHYK2Fv7b7rMlQBReDdKwcMgZjDkPGcreZsR2W
jIzrcMa3tABFH44aInwoJWZHjtRDsUXBL6j6ZHrXZFjjqQz971zd01Wtf1IRcjul7/exfjAeaY/c
jWLAOUB9CpMWEY6ijLe6VGo6dcjo1qmcy66fALXEITWW50n2uj76cups7zXTcNvzRHqIwDgk2MhE
MqvwidTHNa5cZ6Lc5QoEyx2ZHXYFTZEodnXPhPCKGdEFig713cIGhEIRy6tiZsh+qZE2YaxYXqnu
3k3hOoWAMZLBCgfIwws7MQftAfl2V+ZSkc81R7Mvgeg6q3kwFE0bXaybpaFEkYB4HcV/m1O1IXXn
yXvg2cwayCNUVxKNI8pcmovXkYqDRyogiHQOKbgY/5waZykGwSqYGMUbVMBFUKWOFePkK6AgHfpw
Kd4/3diEWtub3VOyQAgBDuzhfqp6rg+A8HhLzH+MI51u2zpgsvecfok6rPEFIqbKE5KP1pnUoedX
nRnvDKL1oT5TY8kohR2odOVW2z3Pt/7HzlFLwO2KVDXtPVw4ZKuTOB+z7RHZkJHQy+fXZ9BedGTM
fXaZoYO9CDw85AL1o4f/0MbA/1DpwguaT3xyaXkamVxQRjC06mm2JjCN9lR/8ep3OC+8Kxw+YSv1
B3y8+vxdjgyFymqZsP4BNKDPAvp/47Df0Kox9pOnj+rVVgqakovC3de14fIwMrPlGp61Yi8gDOKd
J0ncf2lB3H1lWqWJ9Yub21SL3O/GxomiaHer2wfsXL2BcLW6ghRei0BXmy8ul71IZtRoKQKeoKLS
DS0Scnj1uBEECSyY7v6u9TvNRRIc7UkazIcd0Gv5Pw+1q8GGtB5OxEuJPEv1W21zp4qOjfH4YuT2
ke7bfuZF3nMiBjJ5X4HPgKA2WwZXy93z0+HpChxriNtdRKZtk642H0Kc1/PpvlLa4+2sPeWNcxzx
6ILaoynajuI1u9nhv+UFjwYrLyO3k8+8jWGHq5eeYNFw5s22kHUWx9+YGV8zi6yeY4Cgd88GTqF8
RQkY3ewERbqzrviHCeToXL93glQh8MYVvKQnA2CqlnARzBNMxpLGRWTR34rv/dqjIKvw+4hQ5GpV
y6Zk/lab+Gm7H7kx+YDBP0yZhXiG/AdqA/8Z8oV3g0lF1dhbMbb2Vd4drVZnReFzOCiTQrMj0c1T
6si9UO12G4qrCeMez86rDfT8BrWuxI08AewAuSfttfM3GjfTelaD/DoZ4cOyGOrVAm4LG8S2bfhh
bkM5WXVw8gTjtuecXiqVTBeScyPtBhnaYRjVq4nctfkUzwe8jd3579ZtOJCk4+Bl1MOHGZl9x4bL
xMp0x3uoTLn5qdxBxtWgBCjfe9f88X7YinY09kalNlYkNfv9RE+4aIAS8gyVWRjN439gHKSmlCpq
rQcztTNlaU0XyDO1CoMw50Ko2ZoeZHHA5Oq9ZGN1LumotcamWi6vGRdHc5ygjqvx8t63MO33HA0h
Q4M+jWPmCHvBiyTkA7j/msljgdkNVXdYIWgBVzohCAn/nGhzvyDolgwaeHhSCn9Rz0Cyg9N6qSra
zgnfS6jiknVoK20v0Hyuk8hpa/kSzoLaqNrpuTrmwfYd6BjfEeHQNVrPhgtXma95xN+J9JG/jjrF
N4/68/IwacKq4Hf8gNZfiQbH0UM6HFEkSgkhjQuJMefnASA22MLWgyT4sqHtQBirY8mUh4j0YJmm
ZySqH5ERdxi6grGEfz3gCLf/kGoaPNknXmfAnjcS17N4s7Hd3r6elE2eX5R6CMqL2uFpFtpTpmbM
XR9HakEOozeVH+OT4fjNCge2Xq9R6hTi0Lc+ingzfUcS0WVZCNKO2ZMiWO9a08b2L66wqzBcC/EG
ByEzEu1aOW1womqLvPH6sHGquA6P1GVRKul4qGB6C/dAuJ1/UPoNoGIrbnUornB67/+B8bGLWpXr
xdDUUCH100SHy3ZUmJE8d2PYGOC9+d74gWdEOVJ6/hepgiWqfpkXkSHTyezpNjLdio9oox7EcAfZ
EHpEzHUw2EteJjWGkAK+MOesx8lWlCFBZzxrraMuWkSf4sId4Z+TIh0sbro1xb/+W8keyz0+GYYB
u5ogs2fGjIE93moCoifxQJ9nWjc0ur4CgJ5GvWE8kurtyILq6/r8LyC7RThmXt5obfbCj9vuiNEr
kjLoDsbHngeDTLjwb+w27P3BiHhkyKL3KSJdU1oEm2IjWbgJYmbqekxjS5EPL+XNGxSzop2XVtTq
/0W9Fg5CaZ+1BVqpJLa7a/jqow1Eobww3wszwLyon/gpdwpM/llOe7vQvJy9fgCovHztsBITVSne
KU4H46mYa+RbOBtkNW73zqZOdCbvGfnGMxtOYVvA2U7iTLs20Z0p7hsSFLpr6anOg2E5yGhv9v9/
v2LEbIU28AY+yRbh4pTHWk/Oc/tQbKoY6jXkziHWnuChfi+goyc3dR1jrM3gI4oedi1d3uL3fw1v
chdR3ETpuRlkyaNLCMAcJ0rl4C3BbUaUyZXrcEEq7F7TcKWDfTFvzUb6NlanJuqdJA/v48s6rYkA
NHSTqCiqrbiBljRHEfXgtQ7oiIDSAg6U2/Q87RSChBDnzUSDG3QuXPz5XHfy7+0kssdErs4wSYdx
20CuhuMZtU4Vr2UYKPtuK7A/1saSv1qOpIAtAW7JBixQ9UVfjPGOD13bS01mtTgvOrBSP8JbCJye
6h1K3KmfWC3+5TRaShPJUbaORxBWJMpzDFm/RWGavTxhojQtACp/rVZuSCNq1cKnsOr0GLbHzJkF
qOmETx/0I1nAsqgWQT13VkhazjI/8o1b7d2+v2eKeU5FnlcyAPDx3scq0YsktclCLRXDZWof8/7q
pp5CUoUh88W5VZt4W2ECnoMC5OWd5iOMeP624iqHj60uTh3cCyX0YZxdgOqqBhYvyCrUElovQ69S
wdW1J7h6yhE6MDMjo/aVB6658kddwyviYELr7TH3FcR4YIc0C6MuLYwMIaJxT8kFitFnsDbrKeLA
CRv3densXptuSVbPClM9Sn9sZZR8QI8ojYaOHd6/smOEGeQTwkmJTIfXQHIlA+DMNOtzCRUIHPoi
DWydAuMbPZbSltLxGTwm9+aXCenDxvPfLJjSCVLdtxKK0n6u2zojskjdAaWAn/qqYQHicbeWAmhO
ktq7YqtWyyVsn+KTPryCC4/SpGOPydgAnLQo7g3G7Ez0DtXIfBLhbIOW8WVYVkUC0S5mvo3C2vxm
bx5poVo3OLNhuk2H5F2eYLhbW9IQz0IPdEhTeHzOARrXMx8PlhBiCS0WwkhjECHh3/xoYbfH+cZr
+d9HmHEhiK/2sw9pzj62nILA11uPNITpd9QFG4ai/6pD/t2Uw7r69IRicX7+GoPy7yH95NnM1PRs
9dWPwb89gav4Z7aQWkua9zGnOiaecJF7VQt05N3qC8zzUJ8Wp/2Iwlzl/x4kW2qoNipQUA6DL4EI
IGQkunMpBEcNxPgRSPkbdjOM+Ynn/7XqWHfOxrtKo6IPYtBK/4KsPgunGEVqP794CJkJDBv0y/g7
JSvgTm7QjI/D29oEBz9/U/ms154N78BehrXT06gPSvxiciyvgCPf+jdHNwsAgJb27aPvAopzS0fx
OD0ASFCBvkBxjCLyDFiy0125cddeeHDPTJId1HKlDecIW8ZMYnaD8Z2tmpSqpxq3R2gPet+Qf94+
5K6ZjnaG7cNFsgng5NMamKQDZywbsCpXDzJKlGq/bpey2+G7+xrMnqM92SsdtLURwEpuvTaWv/vD
DpiLOcq3YD30ipy/aY60ucOSK1nPHLLQiPuhhJkr4KIqX9VJ07plIGyrCheqeQ/CmgugUTReHrm6
chkc9Q11H/vsHkPkCcuHDzNb1p6Ac+heQIGhBLwoPfbkbA9BW0ej+D0WNRXeQUqzR03FNSbvtcI/
T3BRrGGA90HHw9SQZQ119hm74qhfUrjIBDQrJRvb563L2qVxXQhhl5dX8zGiWaRPchgXlMY0McTh
cpZw0lyl3RyftfJy19M8yxZEq76lAJVoFh9kA5aEhXdYoytEu1sBGAP5foDN6M8CmbE0qc9kzq1C
UztTm6hUROc9HTChDZ68gVCrwTA7jgxPk5sM8qiAZkcd/u1/v20zcCDpP1s7LFVJPpb8kJ0SOSwe
oVgqlL6VkAlms/ymmXG4ppnHpftxdKQabSq/+QhQ8fsu7pPnJOQNzoE4An9C1UgWrBy9OUoLUs8F
IKP3NUqui38iX3r9l7aIJysgFwovaEJjmV/UFRGVUUg62iZfVekO5EWtRW0DP77aP188bKvc3A8V
hnTa2zf5+Wr+CHkNcgV2GclccTlgp3M4PnDH0VnNRk/meYmmUuBXhwza200F/Zg1GD15C5J4pyNE
tGLV7J1MjCtnzGOSmfzkdX8XbbgFOYURYwLTCPhouV2bHLW3flaFoNeMymz3dHIJkuNDruUEj89W
9Ou2e7ze/ZGKYoRw8hicwNa5MrS6GtCrMiR7/Fe3Lod4AyWwM4KGOGvuIvEXM+7lIq/ZIaGZa06S
J8d1kpln8E+ZTEvyYvgKkqG/owXhCeRt3oO7bBmjHYb84EtdWq5mU2qJt4l6qD1yAv3IUMSdjv2a
CN4tG9/HPVCUYjqUL5P4tc8lo1dPGY5YqOTA+b9FM4731W15lQcx1QUqu2iH+xd6+X2/Jp2AaoSm
ZQtd9q9C4qEAkNpLhMEMibsIxOrzZLdBAz1ve2VXUCctE6YnhGECEbNN6Pj1jTK6Wa/W6qwoquMR
rOyYhY01GDPv3czX1e0rvNWo4lT+Lk6cY2kybqfh6RTfEmgIPFeNi/RY7EKzx9MVoftR8uvco2fB
iRSHF08jBiXzHJLND0Dvxf+MCz/5VqpkYTtt2lYxOLCBrCjcvSKkDvi4CcTW7BfsMZV/f99uihjN
sXmEg9t4HsjXFezF5DhQcWyQ/+zpmqAEW/UIDnbezBIYYL3gmlnS0YzpsiUrSynUr/LT2vP2PE/r
JBgmUBnUemIzrsQXWeOtLhlSVeopZFk5Xb+xom3MNZDLMPQF6Y8zNHOeGumreEMF0OErNmIiCjm2
AKIVWH4NqNk+JHLdSgs4EdDsz9Rp9YcstXm+shGqu7USstN7DZYS+r4AE5fvipupWeqakFOMrI2V
L6bUsJKAN7tl9giZIDgv8nWlQgex62lC8FGxDUSTaaKJc9nDIT4kpYmrXorysTnSdQz63Xi25Rq3
Mk8h30kCM1TWJNlqLE0VwL6wg369YLhmVIOE6I18fAMhutqHCtd5Vtfy2SLrh7swoGnUPFL8W1HO
MSytyEJbXEcz3+ViPdEYRwzTzj73tW4YLUdhJ8yMtjxgfzIZOh32+ft8EZjOWy4rSHwfQH1D788F
mCIGEtuZoWHVWrd0A5J7jl2CvLyDGNAVgUjjCMHvH1EsMCOX2XWCFwjoVjsgyOPOSIu/XQSf16qt
zOYdB3xMKu4r48SednIgD3bk5uTmuXxuI57E+qGbqYJv4eodcyE36enxOiH7KREXKrRZegA/fhUc
9BH8ZLMh2fZKiB8Zp66jUkZ5GSC8HUPxxnt8I/eb6I8Yp1KrOJa8AFQbZSqDDckKXQhoqMi7zvHm
dfOMBRWrs1ssuYtGoSaJBkuJMBRllxar4NtV4k/brMOZRGG3MzTGTAXsUgO19W43fOQTEIbL1mvn
jie6QCZY20QVW9zt9zIJs2nDsFnXhyTdkENz+KkTFgrvcUraymXqwTn1eE/6Gz0c0zbOWL+vVivk
LN4rgtjaG9TwF5LwlTuxVN0sI8tOZBEk7qJUv2H0M2DVWovnyWv9LRqJSuL19lYPrXdsRW2F1OA4
RvYIPbwMQoQlnd230dDVjMOUlXT3KZohTTkQtFlRg4Gs3e/HauCITZfXnd6okQY3IDc8EOaNmrU7
z5TT1fhdK3qmeT3iZNO4B1ub89ustvFFRrcOb50JQ/fyAJ4xy18oVUZZsZbN3Ydli2HxC4XD37EH
8XsOZVEfy7gB11YDhLg2IyyjXTOT/FUo5f8qqg9rtWM7kp+sA+Dzp+k0SVrPkcl+RcfY8fa/DpRT
GjpJzK7nrDd69BXYuLHjn9sJAo/afBu8CDDyGgQT0QnnwutLbDT/vukVwlorSaIChL3K2FJhL7UU
78bOZHIEq6qcAzbQXX/bdKFpZD7oyRiUa/eAnvQCLBz0ciMQGmuj0qqXMnRlXp2liug//PsV/qxv
MraxTL9B44DFtz6GwWSmNnmcV8YufDMe98Non4jpUO4rgZ+7buLejzYd2bgLOlwdipmV8owO55/F
+DoxnWP9OZs/92IdMB3E/o74PyBh7SMh5U78Hir7huFPm1Ovrdl5lrTM4uTOEy7qIW5aJuU7gP5p
zpfYSCoHZf8t+qGcwijhwegK8gGT34BsqcHBvcEvlm8rcOqpuuxbWrzrvOp1isEQ0TfMMEhfnXqR
dWu1Lh+7Y8F3pqsZUaPzbViWpdgi+LRWsplVEec3oBuO+Z0iKQk9OnLYxEk/c1U+pglD0mXFK3NV
K+b8/3+q45gWShC7bFvJbFFNQf6F0Wrm9lV0Oy6Aq997fQR6Go/fK8ujWtPlYkbi0/1mdYix+BAx
xFOiHONekwZNNAs0OI6/9cQyiRg3HKIuSP7FF7y309qlif/Z9YNiaPSz4M5doDZxVwL7Qzl7vI2e
0lPY1HdPlFHcI1i34TF1GjDJgNiMDmwOIKq4Eudbz5QpdlM7zr6+Xxyc9PO3RzoOtosv9ez8Y+mT
kU44U7+NmhR0e28AOi4nFgOeJhEI0I2+A85O8whP0WBruoaXYjQGImVmK8nCQmVUrNlfcdzgoHiV
mouxbOMm1Lj+QbgOVOyaww7sKhJWKhg01kAqJX3C6er/9cRllcqt6s+aBJLf60t5kvw6WiKsmbDN
MXzrYmV2R13hjCDgpHxlK98keQQDIsxFzGqndmlddvgJQpqaVVi+5Z6yTMBCZBUGBgx0TWP77iHl
MD7qywVH88HQJAgzF81DANlJFf/RDKkp1OZUn22VVWSPd2yJ7UrC3BpboHzOIApMZv3slClMlvg8
V12PlDdp+pcfI001X9mnSozJIS+chPcmg802ibFjwE9mLRM6jPyzQQFtdSeF1fd1lAO1NxF+5bCM
stTFi9lwyjDj+2g3fwWFaGJA7SXTNhyVP6mVdSEq+r7OU6u5xuPlVOr679uUwbZbDa439KLrTq6r
4+e7MVWY1YCuE3a0H7y8vByydmiVUkrC6qlSO7gh1zFL2kJJLT7UwbQOkGMys7Ye2AipHsIt515G
is4yPUpj+z2aeKt9hnQKs2KSNJrXb8w3+zVo1wLrmRNDvYAMmmUG6TwldxorQfVZJwO8ADRuo07M
ozzaM76GHW28Y795PUJEk8SxUFdoDeKG3LhgfO1Uh9xlIHisS3xjQmhPj+2tRzz7ehTHuAlQGPds
hcagHA+Ww+UncePDSave89AbjAHUQ1J/JxQrny47c0ktyW2vcUV9fD7IcW6Yp+5qjn2H+sANUSH7
MmYDkuL9jmYo+3yeMliEXrgOITm4AmPZ59cY0auOoB6d0csNiy+eE+BlcWtZZN5+WzYE39PaBGpb
u0MmE7fDA+6yWdGa7GNjL8dMGICpxDAdhWbcaa7EfIKsuyaNXsBpOZlLu3UsX8XvbtdE0gpqdBW3
bDIBsRd/MiIU1K9yBsdPXXaG/OVa+Kog1kVnvs+XrqPscMX7LhqdVozEedU6mU/2nKSeF7N/wH8G
o5GM6yARLkQdIFlnb6AwN4McTrxSeEY4j3V5StIMoMimc74hPrZefzvj/UGIiYdj7APH5XEP/RUN
h1BK8pE+JSmmXt7UrvQ8BRi04Pfq3DrBccUvgFOsi6Ck9ntJ10Be29OvPi/opO7HMDG1IXIbmGtt
6o3KmV9wvFB73U7rHQDtU5akkhuISkMRdS7kwnx9hKpQfL/++tkHHTcEEeIhYhVfE7RNliH0dG+M
q4DCzYceS19xHudCOMCpF4G7PyczNRgx3q6IdieWEd1VbfirP1xHUskClWjfxzeHvpQnaO0h+KGh
6b58/83bNwMm3chuAq1zNHzUB6BZtFBln8hcZM9IrdwxDF+02LPIqO+pya1oc2AJa2zpjmpTn8my
w3Sqb1Io2XUNpW15ChgXX6VzL4a66fuQEUThcYmOl1HBHfjBP4YdGhEOtQNV5bI7jOnmq6udoi4V
xdQ09Q00+gwYs+nGiKaiZlOgTBC23CkKIPG+qTG6suoa6oy0ZaTCkd0ILFcjVoI+ZXbMd2CpY2Zi
yDgTI/BEizesIMa7bvrnQXqv1V6WH8ivc7TqVAGgBKtnYbzwK1nlJ4Vpk6H7PFO+zcFQYGVMQfCs
fRwR3YZheh84cWQ7J1p0RDroX4RkGWeD5ablF+lgqze7RRkVDxjukPXbpneVofABP+K73AQCnGIT
rn0ufKQdkDMAZhQ8g6WlyWEuTqCjIlibwdLOG1GTYk6HgVWE30hgQ007C/MwHDV9gFV0w0UqFOlX
HlCoo9Oy9EhHkr4zLBj4XZtpdtTabLRKcd/6FDyPq8i7TnIJD870zHmc7w0k9ZhD7DnduT1TuKDh
DeHh0YVIjEh4fEFqipNMolEorvQXCrduFBSZXJPS2rfVRWXXVrBPHirH84+Jey3U5NilXNoKPh9a
XV6RxL3dIgB6GS9NVoQGd92jg+TsQXdRs7ky9LDj6DotlM4KEJNHGfMgHYGEysPB2UggLeDAC0AZ
RcBm7s7qC2Kxr4+zxZtfV9Qg/D8oylQchyLCqEKQGAqyN4tUqocEJ4fghJ4hVhikmiATQpAYWOEM
vmNw/7pP1MElyJdCW6algUA83mMIFBBfcoLzNQUW+yP8mLs+dz2WNLAd2UmM1fPuiHqiFL/rEOSd
TlgBai0RTafySvCBWB3AENYulbh7ZU1gji3Cp/SBfn95UzfUv/harXXqIENTglO+VdF5tNF+wX6A
/pqGvAbLauatXu+ZQYhxlN0C3WNcustBB37N50ATpS4euzpK1LyK/9Bz5oUYKnMQUJJapAVTj4wB
84TEs7bFP9dPczU9luWWAcco42YlIoY7pdWKG5mOpuyzSe9jkb9XHvGa/WivYcYVbqjmN+yIw9le
0gvcZOs8x6/egitAG50ZMavp1uDXaBM2OWK3hJYobzgn9M7SKOX7YKM4c7oTGse400TaEDtYOek2
c5TmlRkwcW5J3rbinZ/DCY2Q1PywZ2AYXCOgy89AQLQjzR2DXVj11i39AB0uAeLLS0eQaNs97f7D
4aTkJAGkQRuGJi/EoFh4/btd8EFRzdxyC67J50FAy0ypgOVqMDM1vFDXZwHWiQhDA2QvoW8u1EYI
Uo9YyjqbtVurzPS2yLWthYgO7gTQCTKLejizuyk1Ea+0Y5FY+Dlr6jb0x7luedDfbvXiM+QIOWK8
uEwT3995i0yRp4sdXKlWFaLuXt8LYyq4352tcOUNErMSGiUzoqMAlQCsYp5p7nUJGZ92T+dg5n2g
ua+PG/sXJcY6dxvRq2+tbXDko6DvHidu6Bkw8oEeO60Xbso7RhO2CDPikmhjWxjM73Ar1gIX9BUc
+0TjNohE4etJROB+f1RKCBQpxI0vABMq66SK+Q6KSsgRpUQPTuLaH79uWHYk6TtHoKvqw8L6IGHY
KGP3lV34O0mslHCJV6WfBlr1ntxjYsQVW4ZaN5RpmDbCazfkLO9TKRZPL1PHPJiseXCXVgPBJzyN
40UJZrBLmFe11NunWmzt04aCd2TYoGdL4ASNWrhaHvzkV/EdHTFvJQfNZSaAVXc6DSHVjb7F9GIZ
IAzsCBIEpF1wyczJF0JFOyzfhqZWoC/Rc4GeunjBYjK156/IMGAZhQREYIbt1sKHrPLBPgjwIjpM
TivWlqHlCXKN+pI1K0sELe1KsF/M48+4dRqNZrZoKPX4UtkGUEmnmyFakqbKvKT1IGEnR+hVxC+m
3bLjhCh4BIo8w6v56vDsXpoibGSUNycc8fUXjHFWW1pI8K+zfcY3HcfFrlxJYBYictUIG+mmFw4X
YG/wJli3xgqeNiJDK/ztZ6n84eLffjx3JGR8vPauaHQf91xbPJoyVe7NqIhJLvL8Gm3Vu5z/fGdW
vkYgq97B5PeZuQd2F7pHlxyKxdGWE9G6n4PNShkl0YaGoQIYttxQ5rviXVs7R29OcYLU8/iDsYXf
UzSMFY8ZkrZwawaqfRFboH4uemK/6GdATLuEt5P9mtABBpGgR0HAlN5j+FjFPK0HzOERCJlcnTXQ
H4bWruVbeLR72Dng4W8y1Cd4KbQQoganOIZ64mgHTIfccQAfFc4rrrXNr6hrH2S+g9oUs5kQDS93
Ft081/rtLYJk288K+Elu5uXnawVBOKQh7NhtPv9dpZpzkHlMjRJiPGflnSessLVbEoz0GlJNoKYj
C3BaDu8JDHXJ45YLPAl5aer4eRRDw/Y7FCA5LRjMt/kHOqjuS6CqGNP7kFBRTmDyAPwS2ZMFJSbR
Wnpgs7qUWNbC1nXrXRjXC/+bj6GmsWtsrEt8ZlwXpi7mbchHl1kIp/DkZUiMyQt9trzdTpQD3/ju
X/KkE7pIFR2IdGZDWwErEZ2dtnZvSCoya/BjhpSGGTBfThwblW/bg6Bq/lXYgq2eht0+IJMyU3CE
IBhB9LANOozPsuLvzR0ePY+kElvfL8pcB24vgT4BksdBTrlDtgKMvT68vKw6YlscTccvEZSwQR1c
uMc9Mzl7yKUwP6fVPdb/+EAiZqQpFlUfFWKXQdRinz8Z5ctGIWgrSwwFeLCiidTdY0BLOnq6tcWW
3qeSut0aZtBI3N4uXGbSGiwj5hGchrnYNRdmOxHr7eWVgdWdDU134038bemSEr1Maysvn+08oE+8
nGt2zFZfxAP5a502vhnUmzni/K4rQr2PUL3S6JawdsI6mGY8D/LlGHdeppSoDC/Hw6D3ZcOucYNf
uDStAKh74XuJ1FsRteuHCyd6GttX/9P6NH8FLoASqUU2NRk+J/em43Hl6HLgFWhvynneRjBB+3SF
mKO2+YqmIKXjYwGQEOBYEhZeF/6iSPG4VwTdI2TufVugvqV4SeOQzhpV6Ftptd+8Sc0zQRnBbSpa
PUDC1VKA35HBZLO9bDTjpGkztiGTBdpdrliHlAFiRRtu7Vf1Yh+Bque8fHuQrMQnQVi2USNWsxH/
hf0wTgP+fWVCi0QcjhrQuUCnnaeuKJwo/0ogsOVtbS8yk1EZAN3FyeJLrKv/uNbJghT+VlMi54sB
VyUirOiz89ggKqbBbGMDNVXaexFY9R8wKGJMQW1ZZWA2gsn4igwMedWg/uYjxzt8+NQk05OdAfLm
/r1KzkJsXxDNo1E7yoZmRO0+/tvCory3gUSh3pyg+Vz6GOFAG805CoNxXXQG0OQJzpqOnibBIKAv
I+EVxx1bGwh5TSz8yNl4x8D/PcoQKCtYlLcGEhzfXTs4DmoIdrT0a+gkaSy77AsOf1ZeNsjyclFi
dEJV8kPtUWSo1asm5iBSgakyN9rXD+bwULLp6zMo/pDxzvZ6rsBd+5ZyyAdckD/zWze886yqO+Hy
WvB6KtsHC6017e1rcU6XNit8jw/t288osVPBsEDKvs1kCoSFzPaYEzoGwA0eTDIN8CUcEDpvLbxS
7P6fEI+ahcF5q6COtMg70epOaIFGp4IiGLxcHbqTPCJ5RWXn6zmD7fUxsNqeFEuC5Hbkl3HjeUst
E9pIy92chL3enwI+yAPiC+ae/GcZOPGMrrfLUUAAiH0uTw5RiQKG1eHlmIzDKKlc4C7DFLXYFrjW
LR/edLIn1kW8m6+VndixI37e/JfU4wwcgOYok+h9EIDYP1qbl8Maor7lmVacRyVYb+RIl7iNV8Qd
do5x4uc2WhiNBg0YjEYo6MKFe9UlxvlGsFYhHMXPh4Qe6Q+AIL1M6/aDTiNtEsZYFaJ7QiV1BliR
NOmtPz0uKFXjnGPeFhC2aIikq5FWScf7aGiCV4+6MCsBuegczSG3ZcOi2pFJKAEh2GG1+HuYEjRU
w3vOw725/jIUm9CrbAx02utzJz4EwlgjPXB1CiB1Fr6hv8mtaeC4KGfyQIt+IeB2L2GOOVpv/J/Z
JQQQ/dWvObt+argzQF4FEmdg8xgMypWUoSgx4p67bByRvUPpXPa9ksU8KkWi2fdkxO100kkz4cxy
RSRHN6reXVno5Miitvbvd6y6qni1f2J5djV1EGm/iDqf/cKQbl8pH/KNRtjrHX505hR6c1FGGUBB
n8hsbNuY+I9a9Y84P/nbfIL2SDcepzg57S5Roe0v2pFySS56EHDGOEn+KPf9V+JtIECTpTH+euO6
2/QKJFpz/JFQM1By54wJAUgNdgM3TNzyDZ3AqrOHm1MGbh0k6qYJo3rdfWBjhePABOucNqxY0WNs
Kj0AH+VB/9Zt9ksrSOCNIdF+yCoPf4udiK77CFraL4HeTTWRc5oXXReb3b15S62uOTPDNpLI3NFN
34zcb3LzAktYJ1BPVFIyS3G41qMAuDiDEk1IE0hL+LOte8u3DCCs8GlfR04usBZqpkJl6c4uJOCo
6DJEeqRxGDo3iPPJ8eau6UHpOjDyNwyW36BY28MggVI0lcKLx/E7/oJRX/t6cehy98cLgcmepskF
WNxfMSHc8jebbrSvW921geVz0u4y9wZjzmLgM0UktIeyKpq0jNPC4JxPorI+sBTsS0/Ton0tjLn8
Ztr3vv+2Rm7+L0+utGFkCkM9nC5h4MZKDuxq5WG0LI2wc2YXtjNNIFRudEPLtxlMZ81KUw9TOObK
hVqUltmtVbbH2+5+MEjUY+lUzIt8cBb2m2FTte/BdT+hdu+6wFRaqWuo7RgA/pVS9QTHNtDAgqU1
Q2bA4M5Yvfh3TLg0/C+a0DDtWmbHc6YYENQfAPXsXO0IdvQzOGPGyuVhFuP0/BK+wuV+I/2UbYr6
nf1Zq/l26dLNH9apZV8+D22Gf9/ztD13oXFSe4LghgeSx+2z1yGUj+EgFCJoIw3229HBaaN2e1VK
bYsk5nrQGrWZ4/ZxFX2BIPOnwFnyQ1F0l2hGyN41sHHZ1KJXsj5CoD3AimztIRQNmQuXk6dlY4hT
GIBpi7Njq75VShHIe1UwEzGznwK1X7prZP/nwJxna6dYbbj7gTdLpQTITdetS8CYSsSyhiDc1JOE
vafsN2MQ/VsVCwT2SwGlCvbYXpJeI6uSbkESR7Ol67NOqcQyHLWoHeBZg3gCErELz/ObzrpPUUaU
NK7QPINoFGBzH05KMX9h5oMCzKheLOGzyPGgln4MnIjEzZm/B1dMqdsIoXpssrZW7TAAt0cHNa10
2LIin67QcmngFp17AYhFyqaJOVN7td4EG4n2UoI++HJdhRV22uXYvGmI5PyOKbnQqO742srqAPJo
UeTuFINfGuYtpA+9av/87f9hjQZLkOX2oSQU8R91nzaGOlcn0wW8n4QQGkaQYWORT/kpn3C9yvis
RwBq0ivRjg2G0/jjNLIuCL5xIkcQZ33h86DdUFsrA8WvrymTOoq385ogKWM2yXRQnty+dGrdI8rV
6pTqaW5dJ5oFtE/soV1gOqforqZScm1dqw0vFE21l7S/R8/96DTTav1Gu4adfwLyC8GN61KpQpkS
iwe9XJ4z+hx3Pe14aRHHpd7pi642dMb0PUdHC0CBUX1FBsyz+B1FlERUUa1eHWOFH2dfE48VTPX5
y/5mFEvv2g7U4fRjRDzgQSGFewg4dBA/LvOsGSaKXlCsMcKXmPTHVtFqBfRttSBpcAD9HBN308V0
uK4evc+osEhrRfbdCqGThwHhibtkYl2ee6bapz/3EsKkQ2QK9njH2bYFme02Q015pre2FiMgYnxj
OViZRVhiytWE2FX16N78GAAWM9EAgbXItLrk+HOFyLZ2YVHrEWhSJxAC94ZPQCIGNywWlBgdou+v
/rLTj29SmUrWRy1Y3MGFxowoYlihRwcZ2y8HQTQpnA8YE7PnhdW/0yxVZnxV2RFbJr6aXZSq0Fji
DzzEt/w9P8Qqvu0IdyCbNedhx+9comwAdlkzPkTGswB3N9EjBHUlKFPROU5NuekvZ2Bj8HjWy2Ih
EZdUdUx6RlJ4+pejH7IFlvvGowA5kZf3myT5tqbmm20rfDn0MZ13Jos3Z6aW1yLhIuA7lEpN9Ubn
JxeYqxRHIICIrX4Zu98XfEVz8H6hOY9btSMsU5sPUZu+qhrLHfzRHeX+xqlsYNIEAFMprjA0B3Cu
e/C0wYPigMnJ4oL4Jlo3Ww5Gc8LsNbQqqAGbW9QED283N4huvjGINzm5EX4SJe2G/hkpoEdsOPgr
Dnd3R92/dpmez/iDkEB+CPj8eEmVDxkT+gpAZubfvvypY7QTKZ/okXOHiTIDkAN/5zPW6Awqwqjp
+VAqiC4ZbRWPoLZPecSF93BRTh2644ItqKnwpNvpxKzLoc38aFVcFSH2h4UWdnxVP/FPjFCyqy2f
nHM/19nDVPpzgGrh5HAmLr8ufrTuR1lWMUEbcjL2TH04JO2USrwZe9kGCIZuz15G7U5Lw/yo8iCp
2RsYyNnUse4xM3GYo8dJ//0w2GTJ2Zh7cPQ3Rpx12K7rXlZDu+nYPNBIqWHCw2x8s4lyNj1qCN5n
dJ6hXm9WV8+/HHLldKIB353lh1mBmHbp2lI/SeacrJT28sG2pJxq1VPL9dOgIXT1iTOxd0AVul8f
1F9w+H1YGIKvYGMSYkqT8OgIUOwDprg5W76MdLt9zWBrURYte2J3+bKrA+YOaqkFou2NK2wDThaB
vLRXnJv+JmFzTp8BB+PhDCDqjM3YCaUViMaWdmHDSk2OmHDUQIp17SC9UevY+BjbW5+yOIJEV2wM
1+bxlKxW7q4IjK1CMt4+B3t8ldcW1+xggM9dW8nqCPnAQXJC0OtSCx3GZXWXVq+9t7rlUVpavjZ8
RLA3iX8mOPQayn8dbPGvmNjak7OQDhMoj3QPhoseIlpJind9GxXEjtY43vCiTS5WxxrgQMP5j1WL
y93+4SCYBcYDnDh2OdY0Jgg4992HjckLgLblvOnb3BHKJhD0nh6i0/bV5hIKo0UWzoBZYzJGpa2b
vlOPl7TRsH2fVaDSyyeV51pBNe0EwM4pPVdBIfMQg2PRRj8weTN859A4PcfHha2uymTTheM9xBfa
CcPjy/EttKs86RFXKJTLwHkXBlPf+7UXsVTEWtgxeNz+WjWgu5XKcxsYE/jEEI7bu1ra/axENxBF
H+abvUqjxfjkDDxebGBIqdNhYTqR1xl7pj/Jwy/VCJUmT652YEcrsKO+mvuPVZErwKMdzZPxJWQR
0lV9BcHkAsg3HFpHfHmmLApV7oU1KxNCDHhfSz7Q0dreU+qQNFbdaFVROpQQFB93wURfIJiM0ppp
zuwkGmcOhnLaRi2kKN4MSS7iIywFyMFhN6eHf9igiYO2k22uS7feK9cAwr8R29o++owwj0CuK6H2
Vli68ObQTR/rD2A71jysts3tQ/YWxf6LwGer/Ku4pKbWrq2TvKUUBreqUnMKx50JQdlIbET/DZoh
+O3vZNJeMGHsdylrxdcD2Jn3eqDvX4QxYHmDAH5OK/g2BDnuoKt8iaPYQs/EHYA+yeaBUBgXu6mV
UC0q+4o9PjUIff2fN2ebu57YYwC2e2vhztynXwiLBKCmLZSJ1fj4l9TJx8fFrJBqSldMI7oMoPZO
CCPibWd7sCZKfeqoiQaY8roBYyK69Tec9VbOyiAVatLCFPzS0yPMNd3hx7G7pwJuHWyyASBrx/4Q
Q/WZu5qmTK1MNH/bAoS3G39XUebwo918q/qYey1bSC17WmsNO09m96/pDtoBHWbAR8I8fAWpNYWC
U9Ach+v34vnH0nqaoUK1F6kDA/Yn2i3re4g/wAjHks0OJ1bVY5w5BZcKd3W07a7ref1YKrnkmWyz
+JkODIph3CiFn50J203MJ8M6cqfcuJYPVizdzhwBF8yABnETxmjhqFwF/Wvb1W9gZOC9r/DQvpnO
HfWjmqyehX9Wjr/wJUI7M38WSCtecZGqoytNqrMy7Uc98IJbZjy1gd9olc+MaR5BZAGI+CsxxMJU
FOoNRhMYlmrhQ0treom7R9qc9uK8P6EJwQ7S8n8WWBPp43sY83zaq/b1gqQxTSRhiVrv5xR0Bmed
LcIvMHAdXpcMeyTClKROlmgRxJnAkHWd6j6I1Ey+lxbx+A7pgrrOdYKCX+bhalp/RihAYjf8drNw
euhLtLVcLFvqQ262e3uE290ZWig21EWmaPIJXMSPJdA+PzrKNtshgz9MjdLoTUlerLsIBn7099JY
jZMwbDneQ1vNQtZvaByf+S6DJadobP5YAXkRjgi95eQQPYozsOFVFiaBObPloZkYFBlb8fmfsKdO
k+OP109pEWEMQUJODuQeKSN32OfyIj/TR50uDRrmgEZEe0b2K/XiMZElw9dRK8uWsZ7QFBiteIx9
nsrSTqT6VKv9GOkDeVCK5nlHWfI6gxIae/RKI4TLfSr87xmxoUl4xsLokaWdVVVcPD9SKM4l3fqd
QaoYbn++3kmkwgUfyf1JtqiJsjfZ+FgM50tzkkcw9u770BXvhHxPDdEKLIkA+FL8kqluN2zodJWB
e2pjWbxg/1Q4b36n1ErdLE5B3T2CUalkEKx7OIW6/dCliZPUrIJi+t9R4EE2DW50R6bEajsI5VqP
QLvki9XV5tNkioTxR4WYkBj0VDy0tHCx+NlW/+WwZoh2UbkOcj1qwKUpaRVcfRyoimgmg0CeoNNK
3YcImAG41cxAtUYlkVm504uGC8w986jZiBWLWANaO8edZmq0SFRcH+wN5jwlZnqmdizTEdwGERrN
Bu33Y76MtbOQ/4CZVY1q3LxNijUsAmxjl4X86nUZDOG6e54ZcIJqGvVaXHF6OZjcACFVhPL8s2CE
jjTG4rgHl+ov9/ce47XJGiFRny4g1BdBwh+DX0Y9mOGbJBXrl5sV5Th+6euPP/pW7djyCNA8dcT/
o18Zp9DwTvgwi2RlbetkCFDgUb8zd1Z9uz/4r4wBn5LjjogAMUqu4BsK/5Nk+I4L502FMJDsfLwS
gZgOJlYkhcaOVbVnHwTzV4/fhgGNCk87lLTAMQQBvhxM5MzXTpwXkILgx1nEL7r3fdxJ7jG6zPUU
HbbBJvHmq3hf5MY2fY7pUDOQecJV5PB9oS5LsuJCy5dh6pEtfiR0ahXLKb5izcYR3wBfFd+rnOth
fF9YAiepsZVK6JpZaZ8MyEvbsZQzDIxc8c3it/ru0/2JGyjGHWlpHHqYpYKtlnDZNiQcXhbDY0Co
Rs7fdUzYw7sggZbuu9yuoHwuZgcQ6Pihs+V7Z3upTu/nWrEhif9T3S+YoBppUfHhDFOPMHiqeX5X
vFp80ftUNNd/d7pgw+Ln6uFxAT7ZIvpYRBsK/K9A33MrZ/PWYCYjoyehgIuNcCYH/kkP7YYSl10J
aCgKceGyN2W+hZH+w2SdsszkS1qGruJ8H9lI1P3jcCS6KG9QNZ9MqRfX5WtOneFGaPhWJJJfmObR
F6Y2gHjXj9k6xKXS7mLXCCAr5n7Fq2/U67UYwDgcMOA//y2fwQ6+h6cas7zFfnnBkTOOd825SJ/e
e0zrBf+CKPbp87WV6XLTSg4nrvxAEzdbF4zKRSJ9StHCumaSiHF2ZEFOnmzjlu+It8ak8LCcQ43l
br440Aap9b5joOg9aaUDlD/luQhqn9WHtPusSl8pYBOKQU0wViFTdkm2WXltMjc3q0UCPEpD1xbe
tQdnRPStU+fMJCB7J8hYFNti064TkUbWnp14ikHNPgl2N5pMI0g4XY5e82nkMiQ4cN6I+FgooEHd
rv2bm7sEpxMezq8rLszon0f89r6gdQLK9KmRn1uYvPWnzMzfcIKKi2K7Gd+2+kva9FFGfRuOOBL3
0fRLLR4ZYepNjFT7/juTgIZqsfx4wQuOQWCd0/BFPgkRAeyimurqKstkp537s3aNJ0xdJBuDbH/U
RjzeHdrwewMa7ljh6ohq8mhwdLCYVlEvvuLtu5vtV+hDKgTgP9p4XtD6uou/Shq4HNYdGzKi/HGI
twpSjoswjmWr6cWW/SUUs3XIkBvmmZhI8UFsy7VFCmx1fUQVu/xFwfNODEJwWpmNfuRr5IVSaeO7
cHJBhJOcof2rb25okFqyUegaBFhMCdKiGHlsZawYXIX9dGwDqTDlnYoDfrYcm5/uufX9rP2WxO7q
/HaqG4qmVFDXSFCJFkAV90ovVX8idqyD9ifWzRrWJIB0GhvRvMiR/ypOtbnElWI5gg+OJrKa3BPT
VDYTqN5Pz0ii0lJfnkenkAJdLKJeEmi9bpgANg5DLfDuHwf2WIUVsJ6Wa8eXX2I7glM7rhC6xPts
uYylPRgD1++N3sNv8SzPDdDqgGYfpb9FuhbRcCfvGZo9kMLJDAJj/VML98jKb6RfDsGSZtCKoR78
XSDoU6gKixt8Mk+buvuZJ4EOADY6GgrvEwTviKo0TJ8Ys8RasaMIXu60WZ9Ji3StY01j3A0XKBHY
KbcIKbUAGW0T8y0fF2/Z+AoNZ4PBl16TPttDzIvFtdvfyviAOZ20hHi2c5NcwOjMCNQ5YRsYQVe3
6xoO7YS8JpqvLzqzR2T1D8HBcHz5W7LZNtwb1Si1XjR6VL7bs7TezGXj6oMEyHcdB/yinsa0SBUT
QHsJMqfhkwFKNDveGp9EkWMFGMteCEtvSzqnnzSaQPLOJa6lkEDa8SxqC84JBW1bDoqFOwrUOK0J
6uWlySFlM7+heYU9ixidoGASlHcDjJLXLTTca8OKL3bX6YyJKXDup+JSjjBnA5oOo4E4NLOyvdPp
rP6owx/6sBxfN2fRMqqz7sA/l34R/3IsnKB65EPcXjPDBzdpEHlHKHQ9s6ohPd+zangkmK3u/a0u
boubLmd5ilRn8O524wMumdBDsBQL3FNDqAwM2Yc1lDRbb21oQg+5CuwP/ENF/GXDYsQoVG254ngW
z/jSAIdZbeGeI3xRTADUaC6Vb/a8QraNmsasDyPEnKtPJfdScdxxk6Uki/ImiSytzsXDiiWcf5rW
Cgd7UtMJjJIkSq1yva7sG7Yvtm1LyXfQBd8CT3hDFZLzBpPtiZowPBt43RxotE54MWbce/6WdLvA
i0rK1Ve21E5SIZF+OWSeY+9pp/pfiXIHqzdht7ZeQcRlFN55zk/q6YAPeRWMSrfwrh6YvuOWZrT5
DeVahbvMmI2tL/8/++QhuL3e/QRQOHEGoqx8WhQGzAnGMWAKCcAKmWqNijJZqFyyLyMeW6wkw168
8whn+0KOzQFfeQthJaafvC7UlQAQoIIzGBgOfswBQlGw9e20J5ZzF8bKKwdO8Wwks44dwJjncfO7
f2oCEjT2xgia9iqypsU4j5v0eSaaSosJBD3OGQp/fVolZoLxk67Slf/OgTyPvKCKG3tMMyjRVkbY
uaYi/7fMvyI+iiqKf+yRh2FWFfj94y3edlWfQbZ9w9ywy9ZQUvhf5IKgVSf+TeJmf9eYyYlh5/Gb
kOfRb3QK0iZXaTeMKOJjv1OAy2FNiOSc4sD6inWF6lSVOIbc7/uN0co80DV9PLjobSHjJ7PUEh6v
KBDpOFDHWHTn8uHVIPcf2ZNjmboKPLcLsyfOFFvXEOuyGeibWNa0xi/w7Rsb846gV9HnpgIpwTjH
O1CMjC7oFreqjiZE3MfHyCnCnvIk2PseboYOizX6yHqlXLmGzFNkJqSvEZWTKM95ykW+7ObbTJLe
fEFXCJ2oNd/soQrcstRHjrI/J5s0bmfUN69Kh/YqC/2Lsks0oInz7fr3hKme2N/HYNqviLPdPA2b
tP3oHu5gNMCE9AAhzc0uvYNY7pcPdf81hrhgfADDHMSnQmxOjARztdkAMubYlymxx4kXVNb4Cdy/
0B1L/n+xxPCE1cdVgc6J1zsCatwcwcSFkATpDwHXvy8oupBwQppZVC+07a3C7UyWAzJJZnReusGi
iDsKW2yc3Amh6MWMhTEpgx9FYPzBkQQAP3qI/NhxMWvUA1j7Az3vc+ss4jnjw7Ztj7qFnPSTuhVg
UYQYfgAfufKa4L1GNGotNMxz2YVV1lLRVY/c6Z4l0WihA4QJlS+KYXDZfA6djDfnBl7fXHWGwcSg
9RAFxhUEl5xQ04TyX+VICISBrH+czjAprxjEhFackiSuHZLiVUaXyO798mzfOdcFncqtJyrPsMbN
IVEtZqV3ji/tm9ic/HPJ1vmLHKJmEi2DfJukGhhPl8Oek4HTUWYhKQA+an00B5Ym3ytPj1AYwr65
GcqmLMnGre0QKJgNucRCbDXdaiXoSEJ61bVqYYlIMwCwOh+b/PzZXcUK+SNIJF2KHD/ysPFtFsZ+
PGbenI+0Diz7I+13Nvqh9uDzO8BJoCtqdVX4IzzqQNQS0CYI8TNzw8g0a/9sR+BZ8fRHOhLBcUpb
CMtihxTscG2D4pWYArv+LHkTxAa+0cIoqMKoy8msBea+Y6GpxqdFwdTtG1irpZF8/pSlacKCY2pI
my1qWeamxS0wB9m3uQubKNsQ/tR+4GViym2fMWN/tuhTr+j7F6IdvVzLyUEsmQfEijGWtfyl/Ih0
STd7Ka0qSTivQgVGHu6PZVXbhYBVJCzMPKvn67U5Cyv6dDPpPf9NeuJnPQ0btd5hlSr0dXtrRIr3
Ig5lNF09cfrKGisnJzD/2JihA0j73uwQTpPAJGexkglv+aWgy2HbPSe5GA3/Fw4CovTRvSbO0+MK
Tq/7e2vZED39j8HwEp/A6IvEjrExeBw/4+lFJee71WC7fxKpOcR0Jo2lOaDyptVscE9hNzs/glxY
xtlce9TObBVJBDe3zROa3Tfqe2hsC0SIbwWg3kL7SGbD3UMPpf930FFmzijhOlgpjVmBPC6rY/pT
lJBtqfpb51+WeKeD3AOeQw/qCeOwsuhgqiGDtIaYAdH858g7uHzXHkFwk/SWsL+1hLIdbB36Tuyr
Z1JLbDLKeYf+VVXsT3cO+6XBHq+G419OlRUVS4fcPE1rWCz2RyQ/7KbdGC9J9W43sg3fsDfiUpJD
7MS78QjpUSR9zTulrs7rIrW+MbFxWm40py1WD50z/DrjtGgvv8cTrafMr7YrzW5h9EbwGA9ZpdXc
tD6E66OKePkEwFdn4ofagtUtFtI3ZGyGraQ3Od33PR+m1s+a54gf+bDyFKefEvs4vZ4P+117SJZJ
q+KaDRRJoV8fzCtY7jlmt1Pz3JJUacfHjZnxamtobpL56Uj1IyQgrstwqNNH1t209h1IK7OgIQ6p
ilB/hPEmhNy2YQXXtAwmJUqsVleuvWoYg70tR7CelcSzQ+Jgamtqi4YC/TT1c6twfxNwppwFidhm
h7ydZ03DqJjTfb/q5kDCIuEuU2Dpi+xULufiEq/dah4rZDYwnf7vb53Pi0JZ95OjHr+lsSFwN8NV
PnAAb+JMKhcPBVQ1q5QrlFRNnFWxGCWHEcBBfbsw9MoOA1e4ntiCP0QTeSMcCd4cxCaXFJUUNzdI
CoFDEAfezKn8YD33MM2CBiWuY8hQof2+jP2l/pQHE8HPZcY0xZIEQ+1+gbesy8iqCXYMxezJj0po
afa6GyFHmHJmUc0SHXyR4hKi1vAjYliIunEBaedKO541mnHjpBcCczEBwjpgbragxV6iKJTEZja7
S82mcZvEW3DNm4JXU7cSmJ4qJ0bFxNZ8vgXDi6UDz9522XhUsCW8hdbE+vyjQI8AcL2wfOC8mBIU
jhhqaJ0rNdYfUceSTSvbROznk78R+5+qrgYduYIm43Bsv8GW6smeF6Ih4AqMerAmFIgohcOoZbDN
kKp3T+9WWxg4JOts+/+oB2LPOaJCCA70ZWWJtY2Y8h5dozXu6K7Cvw1Q2/g6BpSrv/srJdwH5N3l
CKx10poCZNz00t2DUOU+UeZ1ImucYOuq0Upi6c3dYhI4yGm97mHgtJ7RFL40d4eWas2IXvzRsi80
F9nTr4Lcf8oN7Q3sEO3XxEqkW7uCP+rq/22eYfNCTwEFyI5CAPMKo6B+6pqhpXZWn7h5shmECxIX
71mnr1Nbw8PXyE8RJPtBAiappm37jWhdWmpg30f5zqzkq9Oh4B2DquqNGSSy3cBmm3EiNacM2xpO
fIV4ht6vI/dXrtRycL0Eu2suKcji8nDc7EtMIq7Jo+BmJgYPvlBsSeLwpL3g4vJ5Cz7tV09f008B
fcriM3CUqnT/LK9gZmwXTkpXJ6nl2UAwf+0lwHcH0c3VUeLNIFd5Lj1i9gPrSWvRh8UPupCkYn3F
it5MWFy55vR0HfZrS201zB3VyCEehNOVfTyh1s4V3utVIT5Yo7s6SI6tk8ClDqHKJRfld9s+O3VZ
Ag+CixCRgwdMBH1JxlsMg3J7Z9bi0lBjIOAJ/m74Kl+wvmR+zKtebuKUmsfazET1kWmUcuL86J2N
ck90mVsMtalD+rR4SvCTKbsYRclXEVTyiVgsF7Yfm5jifQcLwuaI5dU+zm++3sc9b5BSF+5oGvHh
uebdhBoVbTgPWbyo4EEO+xF2FHWP3GYurn657bKLH95ldS589ysfGigd4G0XSr7A1NwcRjPZbiUt
a0IKdZcjd89HbFXiLVOMHPrKHactlIg3JQKYMIYp3LsVRo0rL0CcJ2o6nlh5TzkVNJ0oWUxYu6xI
WaDRMvEvdH/ksuLl+0hyStXyuOUkw5xN7qlGerPOSWQGzLIv9Dk1FhTFbKAdiKgVjU47q2FA22C3
azwl1l273bmYXHWVmzrpZ5hl15UonQD6K65rX7QV82hjYdnocQHfMFNYaur/t852Qs9kytOZW0zP
gl6aM3kXyIwa14Wp0gkUaMsC0nOdQdztgCr3vbcDIMD8u647GXtKQ3VHK2DVgbcvpBYMiedK4sYU
7/Ylqx0krkIxQXieip2DUBQpqsGmuB4ZCRKQ2mqAXQ/XSG7+jGEzXcfrkKoXPprzcOqQUMpH71t3
vSreUxZ3UmrQkChgj2xJ9epYMr43UBiOto3A3iHexgE9BsEapuuud0TlEPmwbPaqDwXsXZBOfipY
atHcIyXL3deAen/K2aYcEZvADkrGJqNjr8A8q+sLwtz5RPv8e3XiiGSSi57SBEgcjCiEmcaVMYRD
zw2rCzoomGQh4FEtNQieMbGQ39kDLGdSsntID+1oFWRh0Cxx5kI2UhHf5gv9IN7+GKATsKUudfgD
lrHE15h8AoIpz38G5uq9YHqi/J8jRrU8vEHNGIEqmxVX9LPtVs9MwHYiYRRZewQRUCiJaSqp5RBE
Tkv/BlPuIjId6f8ZRol38ZQboWXWoGAoBrmBHJPH2Mt7Xt14HU43Fh0BQqvAFRsQadvWnUFYDXsL
YeF6Vrx8z2eNL4zG1t7Mw7lz8mgR7lECRKbT4l+3M5NzNylE1bgg7h//G+GoNHuKCMCFEEuRROzf
xBN5E1LgXf+SSwR7FsICfcsrSQLw2R2Spvme0HQv3/0zPqmoNI3k2A5vkkL93D7wwdhNqu2GzCOK
18/lSL2LnU+yMzyOr780oNrSnNLNURq0MznzLqEWdmE5F7fh4Zch1li1fE8aVMdNmWzoFsNB9hKA
qhAJuSKNldMwUBpEYbOuhwl1QK4gWLxxM0zFwdVj5ezyboiYQ+0eOlgglI12+ThV3W+uLSm5o0f2
NSHzs9ON8g2qfHieQ08Tnjtga70LlrInXECgR/yHbJLeZU9/4A0w73/GIJBbtS3qLLk6CtsX9fcw
N9cHZd3EdLmnLJw9SwITMd1k1c3Yx6YRldxXaGNprKaeh03O9whvkfd/sU3j2nUmEz+Kh72k+uKz
Fd4VIrewWtsGMVdqURQ0qUP6eMQVDgahGyrnGS1fl7aL3ur7xpRafj/HXp2F+hXqpxPk5+w3YWLS
+paB9bVq0BGovnKnHattVCOpZ7zi3oaSWpz31Q5FTn+zH1ltmxERmydXrgjbJ9S7NdBqecgluJ3M
a+HhuhWY4+/ut6OlOkU/xkNIF0A6Q2yTsnKPASr8aqccz0WBJco1CGNHBPRgi5G4ttOJsLyJNuU9
G2x2NohdQWzkmzgbvan3hJuTOkgMCUE47F0T8Ce3pDjW+U3LStiWgAdM1FYV3z79vysJLh5Oeo5w
Wc3T1Xe8KsS7Jp+vj4iPfdPPBORpBAAMYeu9Cmn0zamOybE5tFSQEL9osTCHAk+uHS5lTzQSMHsu
FSSjuy7vg9T6WBt8pRwyUbksrhqvHdHHzlmjfKYmd6exQ/NZkW4dR3BBNyRoo+1A8iCD9AHss3CT
6wyMW/30UE7z0/EpRWKknby6U5dEho2eWKhCIMtDyiyvpZpoPikFpw3SC3k31EX8FzaS316NjrkC
Re7wDZ7aQyReoiWqA7s9a7+SMTMSKZcmkpktQ81uJgMoaeYgp9G7E2s5IlKt9tycpG0WD+7ZJFTx
dz+QuTE3ADzDiJCuo0DwNQ7WXqRGm5jeYGzvfANT4YSroMLO1mcx893XzO3GGka8NCkSYxvL4siK
v1Evg0Hoj6wSHdgACSjWMLEUMkMxf4NmIpN291SVPt+I/MTwhJkCnjTgORp2d1T7lnO4LkWWBq8o
w4mmcdN/aSuPjt+qCOx1vtny9oAiZbjFhyD56+q03OgeCiuW455E3YKWPNWsTcIZnXSKFvBJUfQm
P0BpMdICSYEVR/jCY8AQF2QF/C2VlQbF7BF/LiVdPytRhOM1dVEoK/RRDgToYK3tOgfjkmscXaVz
BdiB0ySvqb+YsslD2T/ttv33twB0IX1LWEtiFlhZaTgC+vv60V7gGva1c7CKXdeDTgfb+7oLvr85
XIf7KT7IHjfQTE9wLOUiJk4sReTbJQmg4ACHoG/IL8+wO8/WVEF/Ob8cDebSvzjnXIcvAED6MSOH
Ro/CUka3955r2kblNXOvmnc+gST1DP35sd1Ktx3h+qemaYLHRC9g2qf0VkFvGp1ayqbEqbNTrda3
jAsazNUahUJf1t7tzhGUZWU2V8RhefTc08+yCZSYzcRlHXRGd+nPiR+FbFprWUEVxwpfBors/r3q
krrBbs6f7dG4RLKOlNy+Iy+QEurX0x8z+Xx2KKEog4iDFnF9DtH8fkFJQUVJ29y0qhyz8Xwlxn5u
LwjWzcWIrvYf+AH5LIWTcHZ2moPQ/b2+9qkuC0BT5Q3d5sVLkPT/w/UfT4WAqk0ru2razeLdFJ/c
59EG3Oy2YHdpJtwYIpYpWZ86sV/uwzf8RKMvNZPZ3BpumsoRCcs3012qK7fepp6JwD6nGcO9btZF
jRsFxmSH4BsoAv6GzXrHImcvi0XoipPwBPngrARliOtPxj4XS5mXxeRhf9l92hOw1AgSW4DQNYYb
UT/yU48kCIc92cUcek1Aa4QIp7RTppnCWSHaTE16EO0YXIWaID9/h0SS1G0W8arlHXeRCWStmBIL
K+ROsZ0KEzI2ZIL48SR6x2V0BwL9MkHNCEe5TDIuBZFqVMEQ2JpbnMLmwW5EpN6CAUgyXNfXUdxv
bwnJ5Kg9kIpJojWzXXQxQ2+NzJlcZvrFYvGv4beZWKbSQEYnVORMayenqt2jkvpYbCBjUak6sTeX
K0vJHM+oVI0U6Xz6rmyBdbv9jMXG8xGI7D83Vg/uFt2pfGT5ymYFpb1KVMNkBnq+d+fTHO12vpZ5
vYI2WxYZUGBV8p8IlGbEp8aJVrVhhX57wGS4HeeysVnGW1Za0qHDLYcwnicaxI+9Oab0yfuWY82B
y/6Tmn/f7c8KxsW/irQEybG6nffmPbTPgO4HInSCjj5NF0nwcBAUB01f4hN5OLQpRiYXb/nkN6iy
WNo9Ln9kYJyYxoEsGrVWOkw0gXLrkr0OLqX12scKolZQFFQ52L2M8mzRv5EFRHdZhfCa9v2RCriI
WsJlWP9G3IaidckwkIoIQSHx9abl1dWPAAqDYrfB8yRDcvKEZk94hORQCSkWig5Wv3WT8ev6z4z+
I2cMLbMAjpg4CgxZHA+A2vTceEpZPwi4kwBUyLeEsT6X+cuc9ua+EEFHh5+vteCaFUn9thNl4u/0
NQoctU9SWGPW9vMfKUWX4jrp0mCnR6n1TBuEkP2VDxKx2CX5VNlwpXuXTN13RYhD9mb0NXXfyfcs
EugSxCi/zYVxydoL7FuoYrfea5rwREeeLx33LGF0naKTxd6yhm0V4QvbY9FdCXg1el9AwdgOZhqG
QpJm19rTaQ1JNei0dgjivv+mbfQ/cXPATVkVDXw2vKukvwydJXZi3bA+0IvJ/3bqX2kP3TXwRwh6
z7PvFEkTez0hkpNvgGPNprfv6eTIQA5b6Io9Alllw0xmd9sSY58ncdZviDqXEYfHrKA+hwipGNGQ
YFgeXkwPeR806Hc0MplcY3X0CJXHvf8sWVDUJMOZmwQc8BKh5OLDdSnxVNL+18pTPcvOqiR0ySwW
oZS0d0JxHl5eWK9kT4p2vZdKFvTQr/OKYtRpYDkynoK+V98KLFQZPoAB01zAIjkYoGXUw0eJdHqd
vO9sGR6lw6T9nkO++hfhE6+oBJBQXf3zosQAV7VrRoRfLN9lDG+2iVODh6roiH15w/psloOGPY7K
F+peeZ5iUhxcJh/iuqr2XPDyzgmmpS4xKLGZoqlE5t8EC/sKGaOka7021RxRM+RMDggzLt5TGlS4
B+tCouLiwzQJjsfe91OKXI6SH7sp3ZqrsV/Cl3PfTbvk3ce81dIXdh8OUtc0vibEvck/cb7AeMIP
VEavPF9oEkQEWUJuurRCWOcb6UnBut32lmgymaYdQn525wFiGNp8pW82MJRdzJbPAa7s7Pnrtkql
TuTaI8Xh//k2s2Qk5wfuX8Wpyu4+ityNJwHuKgOspmNiPhNEEGNUBxuuyJUW7iqx0HhKLqT/cSvA
kHeKG8s6sZEcJgsHblUkzdBX1T5bRaTcnoW5izdMyV56HURwf7+XPi1rIy6fyIJPoW3luxvIhROu
kF88BBiik2fscQQKo68Bfr/st3Wa44X1Y+AlIxYuYWPkZ3H+GQ3enhcGsh87jrWYhn0Iah8RwWpB
tcGfjrC4WdEFYctJkIW2ClfPSvm7zSv8y9o5FZyR8afIzFpoE/WaNrXwIPJgd9DTsLACqjiF0RLY
ipBgXVSRsEY0L+rIefQYM16fhVttKmLjYi7SrKDqUs07DJvp+Edkw5mZwc3Qgzi1JnbwxRJxic1o
lzgIwOo0C8TixV+NM7dREHuMZPTI6sufe6YOJwcZX8gm2/deyhX8qs7F0t7PV0fsQHirJUgunmxR
THfUvtooL05Gkn8tGhNLOt47zmHvd+7vq90VLGwwHNVCtgLf+E9+sQ1FpXYzH3KNBYzoj7Gmqbdk
5xsVJubCaYM4xj2fRDovCzna771bRE6CVsWj2zgNMpQqV52IdxRAb72S3E6GzYpmyezEuJ3gqdLQ
YTtTqU9gAxlsUgnzwOPbGCMj+vg9EhE176ZOPN5ZsLwPoOZwg151LaaYHrW85J6RlbPPiyGIhVpO
tjlku5FXDVfiZ7ZrqQkCvg4jZwGZW6mIT2te0SRrCZzZcmS6JW7pTA32MXoFjEQw2sg/+A77fked
SINTsulOvoTYB4A9fUIk34K17cGj3hcxW0J7+4iXzTmwogSqP5gfCoA9PntmKf6/Oz2jli1VVQW7
zqduUdi3rZLH3GZBs1H3SL3jxORJR2GmNlfhUwaKhhtGc5oLQ4JRJ069Y5wiZfgDdj3NddJ6ufCl
pIbWYKQBr1EbT/FO06uG3UI3VrrrYtH7EmwMxm81/ezEnTi9BsgHadOHE1zVn1br09BYqhZWMOnp
io0wgJA2rifA4NQp2LmrtsFJkZtfNrV4u7yXEShLRNY8mCahUtcizyY9Wuk9B7FJFcJTCWqEfFfY
VQugXURjW1v6EcH2ivaUQlhEOz9ZtcWZZzQ62VKdKUYC2YkjZIdOpvXe1a0y5tiT+eY/kZz2X5jf
hK2Y5UDaDIRQUTahRQUrcuRGYnSDyiOIHDP7Wr0Y0D8QUaDhU1w8Te1VZ+nBrxkB1/ZqLf35lZaB
lU3VgjDvHbD679nIZ7mLxlSOPWI5yubYhnTUGf0ZjbO4eTVGBSUuR17NHqIiwVHmEzffH8/JSAl8
epnmR39J+26W49/O9kJkrjRo6JToqG7XaAEqPsrgjkByVlYd2MI3KR7ox5wt/KQBPyOuXMDvHXRM
b3cjRd0gFYraxFLKrS2dETtwlDYTIpt66w1sbkyf34fWTmgawx7rx4R0OVNsYBE4lx2LDVWpSvIg
cO0bydnVwEmzRZ0VDRphdnz1MXCdkJ+7gO5FDUiCA+qHkIfDYvKIKS8ONSGll2Iym/Rzm1gpwTPW
0J6tg12e0kSzYOyPt6TvU9wS9E2wV1PREqEB9PEMi/MgYAN98hVlb62EokBenghF+x9KSPdnMmuJ
hwv7VH3zul5FvQMCYntlRIda4XmIs680LPFRGd+eAhgBvGyHk5jgR9GePprVkr5xL07gA5xKIbfs
KPF8vz1OuMATlCvJ5OODEkZz0W5hQCBXveM+0RIJ6ONVz2b+DI6sh3b1teg2z/mbCzK3DtqK2PJz
Z1mWhxrWnC9Hh8wbHLzdfsas+SROfaj6hFlD322XIIlBSXds1gzCvUqztIMwh5SkTDQQjH4L/jla
Xu5WC9ckhXkPdAPIagI9bC+F8EHeB9tKviRWwW/dwyePC6Z3PLWf9fK5DOzOHPOI6jQ29X4Nt/be
vnzrlfXJ5KEGHFkHl/7PTvJkg/1u1UNlxRTTe9vddoyNDaj5o7UJXvvUGYJlNIMFdfjvsHpN4zMa
W4o98N3WMvVeLF7IZ/+n3yu+xYrptNxAsu4E8YoniBal+IGBXjiv6Kx5K3hOF0C+IAhKnKdcnJCF
V68bGwA5pMAE+qTgCrViIf5+FinZ6c2Xgby0iQmyN6cSZYBycWIse84I1hFDXeDsYxvk9jwqj00b
n8iqqGgpGM0brLv29u1YZS/CGSt31r1Z7SACs+mjFo2vovECpER257I698H180Vu4n73PxSMT3kM
YURxs+xndiYdVxo2PDLe+QfZIFhc6tMRxHmzAGdgNhzg7Xo6ZyqITnhc+O+9WVycBng4bc3sPGax
9ZaAym2+ucShZ52o6thb1jZ5LZY+I3NyTPFFueb46J150bSe/V1j16+/ncGR0dhSCwYyEMziPzXf
euCGA84x3WayYdnBd/aXa2v/toup3yj+tXM+T8Lr2dTUUYbSdOc6OZyo9OooGoVGMueUTaZexCy4
D8hSsODYpb0wCFYrNNJ5JeZurPrz/8EdbdwIFknaqoVAsSjQPmeASNx0wxA9bMBTG6+MTmP+QCf0
Rekg7OLXWxpAQrejToJ7In0lv35ohloJSiawDpG2QJ7Ux62vBKV4B2CppWoLf6OaSZy2/VopIDrp
Hx/+8IcuFN5kDR6vo9VlZjM/bpCOdoktuTagEv4Et7LB4RbzSSmFr04e8+jVC8JxpPoyAwgpxIIG
0wsACNlI2Qo/pOOxrSUL16IwZV9OGSl12ubMXIGkR2tfq9lygx6zBWRqxY40OQ30NmyzoiE0l9FR
8cSoltgg0Skerdknb+QVxBQknFdrNbuZxlpPNTlfAr1dS1IgnnOPmByVWT0U2nRu3bZyDcdmEEvo
kI1Xw01FSe1s4905Bgx4jQPbvtCcAlbPWAGNrsdxOGP4X7p3Xm9jdxhnjOJJp0gozwbrhvb3saHu
z5fCZ2kAaD7lnFwVEiYHI+BJovgJVE6YJI0ooq4lZspDx5bolFcu6+p+N367XeR/kUAsWVg63keW
NctjxfHfG2EwACOVRU+WHelN2STtvBnZgQtIVL0P8RxM7kTv2w7jUhBrbXNaI4LUMt5QsxmVdVfV
M6w9Drubn1xzWjwnieBtXau4Q0alyoEV4U20lYvypxYidtq6Sy1pgxK7A9NMeXTgi+Lmc9ZwNMp+
+li9GpNP1OOQCgtJLqOLgt9hqh8ohTk2rEeAdWiUccgEXMRXiLOz5+xHq7MZVorf56jCFPx8g18Y
ufzPW+P2PVuJTvlNCWKwnnS2U3pSnhwBuXPV3wwxNvNQNlnvetjaNG9+Y73/0afNftp2YS5DbZ6y
ZYLSBTi847sxIEuK2QWdtOMXVnufdhtrqpzyjNlZr03ZCn5P/jFiPsGa9x0Swtr0uap8/b29VnAT
Cwj/oDRwYCVo1tC/wVTelMeOuky2ahNs2d5LF9e+FEPeaWYs2IiR0ILq/VOTWnRo86H/KecAwqFc
pQ0U3cGyDYfUV3NSvagN1McN5QVk+bQRiDgyQcQXlGdtCLr6RAP/ZW9IAmptQn+OI53bn9uXg3CU
mkAcqqUKKGYY7ZFosoGZwZBDUdqwRQiy77owh/CxNu5IoTdEyXPB8s2zhk6wYuHttQXunhKnhYUR
iEJCw4KV0VSkbtrtb5P+kqE4TWKOVfSc8F43C/3ac5InyZgy3sNJwRclPTItTW1I5fHaH5PQiPqY
dEWbPZY/ZXtthGDrbP7vS/WLroCUqr2SzBhkestSTXula6wfz5Nl4H3AFz2n/qUqUMjTEjLVKrew
HzgrKPuAzv9U9mor3ATGLZ/Cm65Kq+AqjsL2GNQkisMglFjNpup1Nlh5kLivjNcCa1fzKs27g9Wh
xhLpKTIyC47phPbgNLmjwWI2tMQREf4BR+GySuzrvnr0BmgdMs2PxxJlO6MKeZXQ5obKIIC4+a2l
F/gBU5LCFFhPejb7fbypbjdR3PX+dZUwMkR2gc5zp5BQMiGSc2SXi8Vg/CkWCUNCyq8iw0JUbY6Y
gbq6HHyYFdxWLs2Wu5LHrMXk6MCPcgEodZyDcMXN6ht5I8SMGWmzEBOdXgmUHnqY/P1nWnZg1Utt
lmJLWAiBhngNEZLRwngeqIet4prg164nx5CSPUF2VjZNfYxxp4ip7ErgUi33elVtueVFghYtSUso
4v2I9FU+i2Ly6vqeF/ADuyRua/FRV280kk1az20gEBhP6W27Ran3eQiuBM6po4wgBtdx3oblPlui
Wc2qG6/SFi/sGArrQlQt5ok9LCoA6IGrL8XmJOSXMmSn2KEdqqAwd70Jt9lQJWFnFdFURktzLpm4
W9Etbys9FT0BKCxD74tx2o0iuZBH9kd68CLGficNFZ9opi0RL/P6xqMg22kn9IEOXn10DDXu8M8I
TRYoYB3C5wDijx5b/9ut5Byhz5AqPLDPW9HiowSf+dqRrZo08GXCQtkAi5ouYwd5gG/FQIVCDSqj
SH8GKbZWuSgTvVECh9rylneLxgyHd0jE4QHjDyAXIcT2NkhH27s7n+CPQrZNlmNP/d1JOSN1YNaM
UR03MXz8f7b7pa07xvGgg2JXi/XL1TjX51l/YySKSgs4g2EPM7CMIBQVrhSJh1lIq5RTEuErhihE
RnJliBEpBB0OCy7htPQYar+cm+MzuqIs374NloRFvC8vbe9rOIIGqMFqoPAu+mpRZ2w6wW+WnzNL
NAJorC7sMSoUhvqbJag6SvYqoHQ74M2lqTkrSkS/xPwu3FPZ7AW+5edjttn0DKyZsracyF5X3zur
j1wxEx0G+G0dHW5Dn8kL1dSiMPfvJawbeX61n3Tt/+kXjGpsIZgFakiH2sf80QBDNf308tIgGfpc
KaGp+MA3XvIT/bfKtH/qLpErnUuRBisUee+mJ3Qcs88hf78ksQfxI7jw99qlTjqlBc1trjGHP+8o
bvr7Ac/NxrZk9Oxjb4SeP+hNrJFFEh4Rc8cu2ihTXgw+cdMk7VN7e99KE7WPADBUPa/5Ep3xtiaH
So/Aeuju8z0P5TDOvsweWK7GGZEUbNGqJMYYER2ACoSx3PDH0Sd6WCvKdBH3kjrHQ4qRp3bL4Duy
eW7D5UbdN+xI34kbmVV/Vw4L8ezQ5vrnuDsHZzghlrAhGOkbReXgIsOuPkdAuY6O3dY3om/+McOy
v93ax6iXmjcP3h7QyFuIUr91EYsbiOWy5OQj/+RzGTRF7UkGg/LRKt1cGlUZxRKULqJds1eMuI7w
xLpkYMy/LQFns0IcZ9H8V28q3GSnYhnUrIsw1HAog0N3gtikNPwbg3/TI5WyxqUcWGxq6XdeuNBe
v/QIwhT9z/Vr6Y7kN1A2Q7oP/JLVtjQscGg3le92wJFeH+usoSaFfO85rWW8bd8IqraDSHBOuUhQ
j+/ts5GGtt8g1RWJWf5kOyI5nuqHLR1f/zv3uV1LiOyk29ixld8l6IiKGcLeQY9X7yyQiD1pHP4A
32vDHzIo7r1vl54gOfstidM3VGrGYxUqi8QwIz1Ht0ylenVJ2GaeViRRpNVBcE3Rbtzy78cfVRCp
+kDZHOq5hzc23ltbqX95dm4hvc3FFhHAKP3MTZhNjXQGv0sjRUm7GqQwZy6dEi7g9RScnBBZhBBj
MbqXHtvmddNWDT3R6NbyGJgrsTBrmHqlSiRCVy6l639welphFgxHKORn5r71dj6DhCl7820Dakty
DoT2iN5YBxEmwAZssSvyBqhuS+TKxiUqKziO/tuFxtsE192ag8op08AEn2mDFdXzNb/XuNa0Flbq
/genlV/xZmrvlbrOyh62hYX1PqI+MqK6dFv7ahAL2nhG+hRbmFqxCUdMdJ248/cfiAgXmKJSk5rp
bzQXnaisO+7GwTD716Klk/17+JhBopQcNWY6xHC0gSi7CnSzEmID0+jU5dWVqO2NDBoTYvn5kMrc
Gz92PxI4bWAxbiNZcQ2toC6XOoz6NKU3AqAGrsFzPhBJos+dBMohwurYEA5BXHq71XAr7KWid4Ou
A/u5igN8EgYCI0uLMrVoVfqzVmm6GXwnmgLtKnQE8IRI73o+ZoQBL332nZALdhmVZBqrpqfGzO4W
b2AgTOz4fLuqSQ1s6DwDLPUrbQBUnXNdx6dxXKg04ENFNtaDdi8mYXV8RmcPf7UghYvTVFsQ3/AT
ze0CQt7YLKo3saMUApWMNsGrkFGprnJKm/XpFTlOW9eaiOAFNHt6rgNdWDL4FB7djDNEAk3PqJaP
FrVDAvT6L2ZyVk9BeWKUgeEFvFAHra/0PtMNuxVPmwvgOu+z9JCq90hWpoLeZN9Ogvv8/aXvscnD
1atJCer/WJOPh7B7PerzWMEaZum6P6HuUhn2f0n7tGGTLQouRdCwfP/kZXlhZagNfy6/40f0zY6p
WiozDI6kKjKhE2iiCU6RPPx4IwaAt/dVqm9aa1KOY+NQ8GZLGgCGqy9f7/VRA72YHFkhT3UsFWX8
pIWPSvLD65J5bM56KU2POTI1XJT908+NvTp+dRG21d63WKrZOmQHKuiIq2LwHJYoC43IoCe+b1sI
7y3PJWuhDPxWmRfzhsWuu8mWDUxyVeWm9bdzVB6M7Bi0BApO5BxbfGckJT+YiJQLtdAChcNvwtsp
Ei02aTgTQO6gCUFWZIpbqAHBquuzI69PXt6tQlNH3lsEL8eKICzQFa61YmoZQTUMdY9PStaJD1d7
1sAfj9JqVOKyWgoAbbHi4apcRcRSBjbVCrVjbD2VTj2l8p9qFXtqgVxzeWyf9d1xkxs5JsJqY6hI
KtG35wQ6QLHBXBZd6Q1EmbH2KoCbnpXaywwp4mkZM+UhWx9YXuXuSnBW0CHod5hWp1sBDNtSHYqH
dkFL5InsWSCJSvB1VMtMl/3OOEbxoHvlAYsRR/blnspSSU8Ri0utCsCdkGu/5dfw7gfysQGzjOx/
eZiUUIl0eb0mQtKW1Y3NWahd9uGoYaxOWMm3HVTFAMkpP9yptjCGa/nc4JlJDf72Fd+h/XnORbNr
fkUviP/gVNeZLnO0uoQN4ZkApwggQja3lYKJZK9hII9MtkeENKs7AGpvuJBTIjCeB1xUr1D/0PoC
V9N0+Lo5T2WMu634/OsuPqyIBPTTSLmMPmQFV8ZT+iLeAw15kx3EmNFJWD13thOh86t492o00e9F
sUQ7wOuWMTFIWHxM59BvwZSa5181Ux4C+ziqym9S8LoIR99LJjKQVH4UakygjNqe+rlQV2e7KHyq
MEm+5E/jAHhvwm+taJcHFeL8H76XR3pqHX5clKUacBUOAIdB7RsYLLFGIwaBqqZE8rVpVSyI817i
PTIzrWg3VU+jAKBpwreckxAxehbxViBSg84OGwF/leVFk5t0jy6T0e/TgxRcb0qsrRAkAul7aE3j
6LZItTA1VBa9CF+EFiM8EU/MZAIC9Qj8kNsDzId32wQH9p1P4ujjBWz7RW7w7nNM5OMQbrJnbIy/
nq3v5N+u77VumXZSDY78qTGA7v3JeOVIhnXj4g6XddGcdvHfJ/lbUfKsCkQ/OKRkV0vVig70B0gE
gypJMgi8VKsL6Mx6gr3YT1pwOVf4ZGwrFDz0frmCiXvqVihlVYsq7DvWiw4Qs6f3bR4hNVyEO18N
PffG+sJ5SS4V830ZElq4uEQRHiDPRdFUJixZnM9EQNwrA/jWtd0kEIrnrtq0mf125mVpCwzKSrG3
/34gKq111HHjdP7S2oaN7pFdNcv/WLpgkXRZGIDscCYmuPxnqMSoosQud/aDzwTvttI1fPIY5rbl
q64NPXWMEJIn3XqZJfTg1hPnAeQkgeLuQ/gIZ+9XofusKT/JGG2SEPykyJInaccZEOt2STetsP0M
JmMYD5tn1D087UfDzIx2EMT3xsBOllecpwU4vq8OoHRGpWEj3ojOFataplrzaWMvbnznY8Z1aQ2G
itG9G2/lGLyHUV1z7rZxby/LJoaZxAInIIIuS+ggHSZhW9NvDIh5Moc4/JvljLZFAseV1dc15za/
lJ+49RRxCYGGrXuXIc5n+/v72RdY+wtYXTyqGwTXmSCYB8Mi8lvdcqNOhkBkbq7tUBQ5vBjuRIYc
JubQIl6Jy+cqDPDnZxaexZmpve40h+aHkzOK6qxzjZrsOQMrSj8MWTWJU3HUsxUyTRqaJIreH+Mk
4Eb79chdWgBo2XjacZI8LHkWmFz4GuTc4LDO/0CXWdXDYc991DshdSSlxmd1QV/T05HTA/EsIw1E
XaXVUR7Zo3u34e9/4Q4rtmF6BDVxW3tn1MflcAkOM6gpU3rxrmgewMsHUFTuBGNmBMSMVGRR87t4
IUXaXr3glZGOpBg71FsBqtoyseM+w4x+CI+z4rMwBBQf4OJXYy+SbD2lt61tDzxK+7lQTCM2Hz+p
2Veo6Jfx88G6Az9lkRW0EIT00ZLyyCsV7zkdBsgJVWnqBYvglwk6F7DOI/pQDZbu42h6WwhkHH9p
Qv9isr7r6s40QbOwmt7CaPtg4vMDcFWki0Oo7KBvwCS/AqDbFyI2MBJT8x2UoLhG3a3ZGy4s/8Dm
geEw71aj3DiQlPByCTTqB+5dnOoodZuF638eCjxK14uqOhPjxK2JLCryx/M8urvJLSW3fhi30k3G
LcpZpeVCB0kDKnHdujH7q96F4TbF0/uH4a5sSTXwfWsltH2l9ZDahfVnFLigjWM3pCy+0FcXZqh0
Z1eZyoZ3wOA+LBhKHTPECJvg4k0rsgea3tI/BlJDZe5C8OsgGdez+0KQAsKrvlwIUcZ7ztvDqy5Q
9pDnfkL1R5f5ipR2Bo2Ilp7eEA/1wAifFTIc18+8nAOH1K6k+mBjfeDPrH/VkhQZJxWZ5lhiicAy
OOZZqfUURuWBHdU+5jvmw4a1UG3/S7GK0kEYcp3YlrWdToXPxMrhrUevPqNmruelVKSyQknObBr1
ei7w2E8CJDCwKM5cE97wEUynuH93PJb2+Oo2OsIZ/KyhnXbKvjPMU1UBNBv0Xr15qtvvPPZXAbk2
gdWtCGBFAbMvMKxRSRjT6JVhlKWtoxfWQH4XkwDe4wUZFuJSSzNjINoHvCfDmLTENp3L4Eh98ikk
2KEpkd/Aoxvn8ta/7vtupCIqzd6VWK+PvjzZt5pgXCEAqGTF+vU0pl/KMGUNuB1qx4jKk/KDRudp
7eTh1wTJDXdsLVN2p8K1Mg7sa7Jp257t174tROYxDaIdDirnFfRWAoj1mMTpQARsXGWJlOXqd7Gp
iwnCMwAI9BjT6J1yPaCZVIDFE2nEISNmSvO8JouNI1FPZi8twF9UuCE89wZGwrwZ8GuxmkqLjvFG
zYt+5Ux/aMjkkPbxBgT51FmVraA+1xSFh6WrXfqv7Mlr0duxo+YuyCs333jTMuf2fbt1XlMPhwHV
WmsvURlnyeozfnT3XZ5AJATBE0Lsj6mIKAYPPCLEtWn1gLe179DUj09vedVM0MxkxHbmvW1kfTy6
ZbYl5dapsHG5yaCNwThwCfPiWOT28sjClGXB3z+VxoVJVyZhFwWao/05SE+NLSSRFJ+NnVt25FZm
/shU2VP4+ZutsItkLOxmjWhhOE8itP0uUPe8utyD6Zg+Z8B01GJISfWd/9bvty3dlOI4z5tvhoTI
67326lJM4wqynZ4fdkNCUTUlzYa2B1Ild/TFgVNQMYech5X/+SLpEMIqr5YDg4s4Oa7FYv6rIXss
sdob4WExKT6+ZvN3wMG1IgegBfFmLkpPENJXL7KPQy9HaTbTLo8Y86B9QRk8y7DYGvZNTLScpM0S
L6ftLGeWWdCFJLVwkig4+VgUgJRtzWDVU4dqqrsZ3qgqlkY+Bk/cZcc5rcHRqKYy7b70ZEgUQlDm
FR6sETRFf3iRSBcS3BYGOPU+NQrt+XtLze3eLZ7dC8eJ7is4bmux0So6AL12DjNUbNzPfXbaXJE5
iH3vLZfXwVc0jvN/CBEDmQZST5GNPiKWsPGzmmFzKQqn6R9gGKfe9gO6dxxBkVd8iX5qgXnyk/LI
qaVsPg2GlBVgoQ9KHQosW13IgZFbVOdQjFvCoOcu0T4MuSB/cKYNlgCSdZ07KW4XqqjiFUvACKUl
PIYBrP9WbNveUbPS5DXuZilcLB1fpcwfKO22tVJuZwxDnDJEiuvF3DWdMmtoqvDrO688i7XAxWR2
su3loy254R9lHeGRrWpwWM7qcKRQqTmw53KLbyTmbA7N6F5dx1PeA1wy8UhnNe59JdwRPeBa82k9
MWs5pmYKw/jRNXs94xWyih5nBQFufvFuY0OufwEicxtFfbrbdHrImwMScJnuPSxvCwVdWaV5UcEu
vhPK7dS2nITdyEwnd3iip/VCajZXjyW2RcjArSUeLWXuj3tznvazYxGvYpn/NBmVOsmaHM2CUTEE
7+X5ig3GjDPJWdOKJtwem3tnXI8ERbuQRiH1WJJJlTIAnx4iQ57ZubWp8619q+B6HfLylE/Cw0O6
jW2J5MgsD3c9OWtddBWdvYvAVlvaxHmEp71JxZDs0mfqawEhK0nzQ/JoB16buw4hwtDscw4/ZuKd
Jwgc9tvEukFXVY+LjIJ19JEwA1QLsGyXZlpKrtbFOHeywZQVHf/bcrUFZQMzkpeV5ONGTyvLhA8v
5o1Aqxo3LvRUM8DUKSX+4zq+Sgzj+C/6bYDthaZkORZtVyXvH3TxJBus1JHnmNAgioHFGZ5fhgLJ
9m2V3XfOYn86glFlVyOyOmSytRX4lLmhJP9p7AHot9GeatmEY8C1zX9d7paty+LV/BJv89sp3l4S
R6vh26cH24Up9BSsQ/XAkCanCsJgy62YksjFe9PGJLQddjrv7HSz5cvSSTG9xW78gp5KdjcSW6Iu
oGF6akOzFRQi7fEBE6fW6WTJVgzaRTHOuqqGyR6SUdKOo8rSCb0bqJiKQ/XoD34irNlqPwi+BwD5
tWtcbQBikre7rSQ+wmIWnbBXlYL5Mj2Goqc4BhjjapuBQAgkXeV383B1BegQIKvxWF+QC9nmw2kd
C4Xo2VogNSLqzvFEod7o4J7iP1ekWJ1PDVXC8kOUDIfMuZIJVq7RvbY62gBE0gCysdHREPwiJt3X
7fPpY2PexxFCx6ZmxiltH9TQi7FlyHBP3GLkcpn5sZ6Iay17v2C3fkwpxfsa/oKZ83ycMsJ3t8nJ
M00hN2OKn1OXADDaa2FiyL1dyYhFf3degJTpkcBTrwUxI8gWU85Z+OH5ay1yj0Xq594skmB4gSvK
1Oy0P78fHDrlOgLQgTqXkT2g6ohWeoLhEBZA8HxL6nfGXpZN9ZvSp/Sv/eM7YKHIivDPP7mb1PKe
tyF/YZkQ2iwJgMD4cVr2dSQO7x1y1awZTv9ScgSXhtU5xn0/s/OOe16Vo3i1Te3g5Z8B+GtKyGNB
ndobfB9XbEAZbxt1TeWA1lJ/j3Rh/Z4xz3NoVlWQ7NOXmhG/3HS8cVLf5SPPeN4p7a8PzfmWi4J7
CUZOjwi/epuidAE4LHkY1N7nZhzidxxXqrpY2oaRRK0o/F+dh8/xpyjLZLZcCYGJ1SFETbNyoDBr
veNL602NYAeiy2P/ukmSFk9v16Pw+1r3OhN04cOxeAO/EwQT40lNpAxoQ9J7STHQvda3NGfhuGPP
qqeFh2b16jusSGG1ysutVklMO7d651fFawU1ue6I9JbMBjLHe6y7mybb0cfh0xw0mwiDNNtZ8mp+
Rm3kI5jhxjB4A/gIyG4JfI4u8ZLLg69LYe5B5J1GkwyLhjfhSIlAvVIIiQYOlk0Ham8cZkBCDcXj
77afZdlBP1zriibMymE/CQ4wpqfigw6sV4c5NXrc7iAxued5tdUf+ZQiT+h18m7vw7w2dEqFvJ8V
S2nQ1fORsxfoyElbmNwZvOTA8ahY2Lc5liArtf6JRfjFooXPVOvzds+72+U/xN55cY9JGHv7YX2c
zmWUVyASQHRtfet/9y8SVDRLo6o6UqKtYPkswGxyo2FoEmNIx1m902wg/yuu0Hjs0u6B6uTW1yyo
qqMaRD/SpsO4c3cNYKablYxe5qKi2FbEKjjUlwGhrFEFcAGD/CCju834SKLu/WOpP5meZSUyvVf5
2Pf6McgJeCPR62S8ixFSf2rMpKS10Ifta7EE5Yg0mxJA1fRZamJ2ri/RYtgIU7IIGtZFO3PYBA+j
kvg6M5gnxfWkLBsA6KOzsvM5DLTAHLpz3FmLmdJNEgt9MMfYQWIuomn1tyg4HE/Tf7wJekQ8iwNs
Ij7igQRlbq/qeos9rq6epoulipUoagDXQqwmCkZ+y6Nyn1+cwaLAIJnSTkMpoGVun/khDtUOq+QX
i95mnwGoCVIL4BT8bXeH3wqKronTQDCOxLibq7WVD31Ueha+I93mWdn+MBlxupJ1RGgBrjF8G+5o
SShzUAkxl7DLoY20LMjaOfgKWQcireKnPC9GKrUebgxSmbPoizKw0kArH83Nzf4q5HcINuGYZ4KR
B8YcBd1nE+Wf43JO11GmhpxpYgomjLbddu2/7S7+gy2ByStoU0IzV7C3TlCxbvNXJdx5Mpj06f11
BcctxweiXSZjrGnuSrDJXf5j2+OPbmXCe0/MnEOHDuvsmV8DXzKpnmvjB67aukZ114RZLiKj9RyR
2FnJxrYPcHJCGc2hVeN11XQJH0fLOQlPkMvIRQRCc64GApR7usPbGCtMeQWfIKP0KpPRIt9g0Za9
V01un3D7zDA0wTlJUQRJoEw08yKlJOSTxW/vUf5DvNhRh+xWvuoMwygn2gspC60bLiEi7Dtc3uXn
y62EDXnst7p7b9zM5BmQyH2WwbEjMiyV5C1GL71aPgk04jlpIPdHKuhE7nAuqU3zpFwan8AkM4Ly
rEV0iwUU3MMVzUAvH5BmrwPnZJwDhcHZl0V2GbjhSWjVqi63VS53FoeEHBuHvDhoZRuXosHUuH1I
DRcp8K2ko3ohw1B9c7aYBj2Y21/0Nhf7rvGGBB2SiT0FQ+B1Jy1ZCRrvGyhPk/rZb/MmWwfs4RLX
rHMTmg7wn/UzOpnRqIhTUzIZxbAORycoOIVYA+j5rlPn5KqVZHgEN5dbWrf0kFX7NLm8fF4o3E9z
nuFQL6B0f2w4SSH5auHpq9AyjKJEBw+2qvxkfLDroB0VFigEXcqcaKA0oVXLcerALbiSlI3Eq5TM
2zl9wqebZFCEvqx0OXBV06SU2VZBD+5LDdHl01hyx9qDucZQ6bnizk8Aj18A9gdr3oCGnx282Ipl
/IvRX+NbQPhpqhtB5M51+tKAeNv9X2b1JBanAD3OjjTBPKs96H/tRs1u8k8xIdxYBCRZG43TOOn1
LKYGLv3XTReDpDeNINkMfDpkG8ceFLbaij9j0GiZqDl1VaRRrr4cwcSJnf0lwCTF74A1tGIzZAXN
Zy24EOWWHmq+1lFGnSpPXSM1mo7iUSe8fQH/HYhSRbRlLx3zC1YkXpRJCB2Id/rJBGPjbQXhNfb6
GJlwBmb93+rGFFu17jS4J7X+mZIrvmHY5Ko1uR8GZ0bLNHH05QdPUkd5lbqx0crNjGJsnVE4dRje
Tquz80F7SJQtoe9I+d7+V06JNPB2RelFIjL6Vy/CLlRNcUN/VFLKIKT4W3MLO6dj79sAvZ5gFS+b
z0DZcFg+qPKEYu/OjyiluqgYRLXJGX5+14fEDGs999nfoQEWSiNPIQ28aCCoHaeVWTvgjYc6hNRy
psC0kSy+OQEjWf14ObJDMdzN37aqYyk2dK1ezip6dv5IJBa9A/ephDSa2R05y6U5ftsDcbxMOt0J
r6KDexlnC1eRPrQxDJ6kAHySc2QVzJn+jHXsuvOvDgxs1PRJ0kXLdo1kyaPe9xsa4UV2nulSSikA
b8UVL6w4es4F581Y7HeV0vg30bLbX5u1U49zvjgCf7+2ZroA6keZW3HHcfwm0Ok5eLx1oLLyoEL1
Roffye9E/RAC6YrX9vZRfv5MrlPHjREd8GArADjgy3IB/yAN/rnFs/e4Gk0UuTs4X7CQ19fUcVt0
I8HXUTrl5GY2l4gOzYRVIp7ad2KeQo0btETVbzDcDr45Z/LagQ9Pe0ShBsCVvNq5eXTA1ocz+YSO
QnAe44h/esJOD1VWdGWld24+htdte4MIbv51G0Vo+O5jbmDwBgaNP2y+/y2qJiFvU8RRD0JpxLCX
mBf2duybZpHvmJmh6Dd1pZdfVclLWBDm1i4a5pi6ezOGUH5FlW1n9/9UxMWQTgO3inXn8AxoW4jI
TFoaM3/82BkfNv4xQTm3uAtn9tbinLCx/Q2h92gKqdbCV8lXo3nceHDvsTdiPXhGPgdgO6BwRY2/
hVI+Bp9xffSG0Z9YpqLMyw9uMgVN3gUrtAsIASg/QyM7t3QVsOf7cIo3zbj39ibdMXqKnZyDdTWQ
iApn0BnrIbQGWoBJ7jpoW1/yqvmxurKt8rRe3DGwZkbmUq1jhEc8c2D3fAkX21IbLMcOpsdMtPfA
nm0lPpsEK56gvrcEKWYLdmeQVi1cZ6NvQSvKXb0Ji+Njn7etHjwCZGvGpu6XbMsSzmelrX08n0br
iUNVVrzBjaDOtWHxUpSGiVSj4ia91D1WwEuNXyiBWa/a/m9ecFBzjfYLnSqzkYk5sfoYn3bGBZwY
VEawIgRla/diFpzx4lIvoY9dJ+G05AGDtfKXg66vW4OaYirdO/BEIS+wz/wf5ErDBNoQSr39Xd8X
+81AJ1rwDWeAxZ5ZmVislTkW1FygvmLD2mjtJleO4YWTaduTlVEXJz9518uqYo5VcBHWJvuZAc+2
krP/bo2Nh+tdg4v1/MOMAEEuR3F8x4Tee0asTfZHHhvc1bjK20CXa8R1g5vSeSQY73dA6R8yX/77
eu+wcZ2mh6b+6vKC8a7rTinFYd6m0VggwKOrk8YRY15NWnpKhZa2AKkwdo7bohOYsznJiRQvc3QX
migwLjq9igeOmtuwxTYLVSPnqQl+KSvH1w2DzQWww5/sxyTEwjk7lXaXw8x8EkdcjDs/rAGAvmXu
I8cwk4Qd0UQtxgvZ8XgiyevWLIvol8s8UMavrdTjdGWxBIPGjYl3+wYWvC17ES1b/Dpf8bIJ6JB7
jnseSff5ci51Q0mg/I2FrxJqOsCA0+hODHKaQaumxs/k/ICEXaa3mWggIbfvD+ZQqSpbonsifSPt
noVWTGiI7FB9jzsOoIrjA4crBt9A8NC+Ngo4QwA0RGh76yreDBw4jsIRgEcqPzUkdSnucZn/296T
0xlpxjpNahijjnfif2fnFXCKKJwsA59UIq6kGhJ5NhvzvdHScaQ+ulCgLHQ8IhgbdnkTH0S8g3o3
Bl6LQjpt4aKzz1vVYVel4nNjbT4Q3iHuXWZkOa6FihyYMskj9uUC+A3dtJJVniWBsVIdq60a12q7
1pxDqGiG6BRsSjFuNLd4nBwaPOVVefZ2cn+9wNZth24GiS1AG/pkqEeyBNUjtxAuUUb2ankCS3xb
hJ8NwpBvrfsqBdQf3Oa8wQy1zDDH/KjlcacZD1xmEJtbFotuxIv/jXlyVkDbsdmg5lVfkJnwOZ6W
5xMeJjUTBXrsmfKMA99bR/LV/R/KyeU2rOJydnchKisZCUAW5NS6Dysmm15wn+4UqAmnjLQCFB8p
CGj4OGIqkunKaaw2+wvzmo/jWGlnDIRrPe6xe4eG64dJOoDLQ5qYktQGGsgC38I5PV4izj8GDeQG
Phk9u9RNzp1Qw87f+rbMKxpaSo7UJ1x/JNvdhF+eYP3a6LMk9MYRw1xbYuczeOThNaIQ2P2JEurG
MjU8hV4lR26DWNF6z1Svrq6LoGggGS9aAvaDpxMzN5tXCsF1PritDwsWr0tUpwsVENDS9jc5RXXm
KTuKOKpkTwkeCcSA1LEWqvq8tpiQwOINMhFZ7yxs38c+HtTCUhZ3mx7jLWxfbsx5UhJ6JJxlzh6i
2T9ZqpwPSTTIz1LzYjAaLXjg8/qjoF/N07lxHvI7GErcHoxYCkx3klHYLk42gyFfKvIVh3zBVfDX
y7uWcBgcBtWyQ0oPabEXzqecxcMFES0X+stxZQY2BTB+b3O8tHKOutrwnuJkZ5JPMNi2c1S8gRur
O5NYgcGWUQYVGrW2AEDWr2cmwRymHg+v6hi120NZwcWmgzkgi6C1RpfmNwSfgvQ3FkwKnc2DKQAG
ipymDfzTQ16AQXJYTLHs0dMnMCpPvFISvdj9OHSwsU9yExCldPAhxPDA4UsFDWAqOmGqSqwY+/1o
w6fxHwKNVN0CDpx3F4vTi6RTZxEtb0pAn3yiiFxqYjRwOOMEbsCpJaZeJACi2QuR0ZPbmOS/zcZs
CLqfVUKxOH97biMXPGm+abuI7fbo+6vc29ZKbtGhxG8EyHgf7muKy28LMCzExSV/SHQpGfzu5Mzv
1sUwk/HQ6idQWPPIjHeS5THLU2AKMj1UA7rVFi1YwVfPZsi2fFcq0x6Qr78YsKjVutZt3OQm6guv
u8zI8gf5ZfpHYvq8jEnvgJBLWYpdWvKTi4spbhuwqYOeJ5MYKBf5A5Ih3lwXnnD5Wvo1c+15I93O
hiJDry4NFE9lsBLoGAdDOIXRsH4Pb7OjHNnj2clsAZiDceFzbh6lYrSz3E7kW5LyosqPaZS0EJCV
ggKKlV5fKIzsQvcADzxQIuhhg+21VUu8kVzVBl0JxHN9+PIvWSQfOobH9Oi1x+d9qENO80WtGg0D
W3u/WPUJIAlL4in7GpnAL6nBqSXoYqlhbdZTLHN39vNckgEsRhXnzzE3FDRmw9U/pTBEWowdluGP
unVeKFtCIXywgsPHTFa2wzj21QO8b6J9vkWpL2Km89WoBY/YMfrDNOXBbr4g7HrBsFfAwllXTFhI
tebWIcx1bW9hraM8lzPJzbbOBxpmuRUqxn8poZRBvk884fhvhcAP57kRRVIw94M05GcVWtr/pVNK
O1ybptkq0G3dWne0fn0tQWnDruVIuQLW8L1c81zjiPJu793Q0VVsr6lHzTTqvShlrmES0I9sAv0c
olJY8c9EAeaW26noPHggzl0SVsarfsL64OdEG6PWnWJDUNp002/aEkexGnY4ozPo49Y9iH71mk9N
35RRZAbM4uI5WVq8La0eZbB2x0FJ+6bSw8lAFdM2Wh11y/Z4jKX/RBj7K+VIJnbHxwU8CGcCTFCV
kzDA2qcZN/Ppvnjq29+AtJlJsXH5H0M7YPez8wKBkUra9pTboTTMA5gdiepWFhVzl3hnLoFGft01
nLUx1CaymkBfVDEBpQyu5yQGNA+qwPbf2tPRHCmCKnVpPDmG8oHWqEMmHdl+3uARSxVAgr8frEoo
+6CJ8CznNoB4yZ8Di5lItd2Oq2AXy7+3hqjYooFXAs+kVEhTvISKd7PSjNXJwuqVp3BuieLSmCZP
Zg8CyBPMdckn/L2zRZs0utMHO5Gpkx03i2r11Ol75KiSt7GVuKOhY0ozf0arHmh1UrH9Gmg2Rjdw
OjBgoYqu7XMB849mu9s6XLUK5UMP17lY2/cm6sOvRXXLTZZT973SHL1RoLWGb23XpQoR2aOikcWA
7HFmC4AGO+RYXND63VQ9CRJAZkzQ6JIFTfiXCsGUzC/LGcHeg5rE7y050WAW0eDx5SezXfpWpHn3
8cYuqeAMNY939SNjZkR504D42zqtFJMDlhfMrMkxXAfkHu6Ptu/7qb9IlFATWLPDREWykkVEo9jK
Ct/45hWRVQes9xBaGHpdaE8x/CRNT7lJ9s/a/YxZOUH8slNUQsh5/d40eCYfQED8uIiMgItCr/jo
tPx9qKbBe3mIc+KMt/Dgokn4rcsC6xhbWY47plwJn0eP/tLXwN6ayYgh/n3P179eDSTUrnj+WNb2
YLOyoMt3AkHMYxy++As2U63eOAk02C/KR8F4dOFKwUx1mKV038eu2GS4UXPiUrvluOgqvbuuNdn2
KbEC64ald6tCSe3n+DOhAnqLuQFtE0me4by/X1gWsl5jCciyj3y66sn8T57SqdPKJe0upl7jGBqr
83HZdniSda1S4ncxrvJ/RJl646BCyV8aQ9JiYVrS/HPqFd6PLTYsMkrxlH0GwpGcvXfHHe6w8azy
7Iemz9Ri1PDzn65F18+QTTI9xpdEx88a/xBWpCqWTk+x0r75Ze+6/oFcy93cgtXVYjtcijUCr/PN
1dCE0uLKC/WKrqq8vn0UG7PQSzGhF+zKEIz5vzT03PNFEGXU00OzYW3sG6KhNG4ude+5jlkN0o0r
EJaQSDrmdmc1kHFXNbKW3JroOLcjjJ/GlaOE9pbC986SSPFFUEd+sJ7rXXbWnbZpIqlYoVJZ1/kM
A4jy0DvTFU4U719QVCQIfizGNRRFTwBp3Y4jYN/siBf+Z3cH+9mMnmBgb1P9zT5/6dB3rbuHLmwy
n2qkt5iKLFM95yGN9Yvy7Jca04gHFNQ2zzxi4K+fXA66419SeLKiiIfw9t8c5q/xN+Sj9nIdWNsZ
4AN+L2xoOBU4z05ZcV5YaC1DD1rwPm8TlXh7YErx8g0c4GZWcnexJJRe6oXUIH5iDQOfTHzIJAsP
+7Ov4EkXUNNqLQLFKPElyrjlsm43OL7PRCj3d2rUEIFHwVKtxaXeYrcAd1R5pjLlYSfPVxYyOQli
nzSOzaHHpL8hMWZxipxPFcr145xWBmDtgAnyTy0XlO+4AsJbLrdX63pswP4WdpLogP4jLXFFOVJM
ztDLTJTR3u6KCGujRfbPeAKdieZvChUOzyVMwRRxROO0JhglSp2XnA9qGgYljZIEYyEPMxV5zwN5
CCrF2RG8H1VY4tjfFhxJDB319/Ti6UOCgfWpgYepgZSQRXud3zqvgUvVdTVjLLMEjiBocjckPxHa
daUoehyT/tZsQYhrq+hbvLPunoEsLw669AvjRDAOlZOc02DdyMU6xVCfJQrv54MoRtXjqmIn3+Ko
RE3I4yY9BHqSwNZOLG+2LIEqYMjqtMmxeSN6Vn1NlRwTuygPm/MDRXM6ntXgQP5+EIyYK73LuEik
+jow5ZApXt6rE3GAOW0oge3tRXXtKE/BdjyoscpYTrEAvlX3QbAw6memTHXvMu17+u6NIEwf1uFf
KqcqgM3dLThy4Rtv7ir25gotL2XsPOaRWfhb16itj9Pq+XGXzIxLZtjL4RjPinp8w0G1NG93LPMi
6cS+bPnF4FRozZ+l1RF3qR7gcbArFeuKJcG7LciNHIoPffVRngChJRQPvhd67e49BI2aJyus3PWw
2/Uper/3uZb76QhqnwJxP9SP7h4Q8fA96S7iQYI/hB0Ma8yw3PdgI96GLngiEDOM1twHPbDh3ZTI
qpYA4XzgPtPUqU4FbRNqVqjXviLW3KqnOT2HZn50yNeUW41svTkQ7ON9LzR2IoZeiraUg/U8/JSN
/DSDmjZoeWA5WaoWxz0w417jYcDraD3XdRdmeoEzl3yWH4AnLc1qLe5VykBtA8qzi7dMbdaqN+Au
Wi3iGwawOXJiIIl6wSSq2tWH8VqIdgp4GL+NSEnSJxsECLFYJu5leBiHue9/aNNaEV+z/CQa8W6k
I193J0y0EShd8gRANW+UV7shgSy59zrfFY/Vc8nADQgU8V8q3OymObcz0pfQPz7Xevz49NSGuFZh
29ELoYUJBF4OpZ/cez/UStYS6QJoekubdM6VGCTxKzGAZrKt/tHuNbmAQS4D9qI5+QxE3lVYs/VK
ExfW/1fAe40zh4Vj0l0zKNGxa6FP/ZOScK6IgPY9lkMfmVmG2Jgm7CsS/kpNPm9nATXein3uC+iE
CJUfMSO0ub7Bhp0Fry0XljSi6gPL1p7GXxigjv/+vQKsJ956Ol2mrYdOmVxUNy54OMbknZeukm8i
L8RPcQpLyL/M5fU9VcPWNMo6+7LvrPreLbU87Jckt00I8Sm08BxZm6RtiuRZGKJ0cJv9mlOl2KQT
zO8Hy/6wBxRMQAr0qBeC/n8MYXOMYLv5GF1dojD/MlyP9+KuX9H1chnmcdsehjHe5LRAkEo7PxRK
vpJwWQjRbrL4p6Y2LOD1Jrs9E6N5/Pyvmpf7K0cNujaFNlYIFybnx0GMbH4YJqxbmaaCFXm9CZl/
hJFz8jzRC0R8N4vU65kHsGjeKZkAbWKZ+7AWy3MDduER3MbnX30kR11DIZStxc4ZtX7JM/40QyBs
c+4X0OBlQ4WaIFUZDmhy+KIpNiS6ssL78IiHgfMcO5H62EfsreDmgGpQTwKg1Du7ks1H9tQgAgUg
1O7D4EWamAjC2NAiZBj7xj6QBsmLg3HfQ4QxEHQ/fmXpVGXtfDPVPtp+azcG7W15szl0w9IVlYe3
sYYAxdxbNVspiP11JCMc4NAh60D45uGbbJ2nuWz7z1GcXZJzMXzBMCp17fWqWZYEUs+cus4OkWih
aWx4/PwXKENH/+6qFuD5LOMuWqfAeNXrWXR7WAcX1LJOSnQ5Z2SOW1Ur+pW8HgpTn/Iqu8x12vQ2
2sPDbAbc9yO9FC5IfyHrZNnbjjzOYs8LPklqEQVQD0AAwxKICBAvDdoXUOdssJkgoB2XGezNdiLp
/PhuEM1etIoyp+TQLq9De1YWB5VfKf6tHmqoxF2fkVsOHVePmcqfgJdsu7V6ZoVjhXY+vEXpPflz
q8ZNq7E3zA+1WtJqmVcf8sNFPXNBfOWhxAOsWHZharaYh9yHb8hA8v4h/jl8G3a5ZY6AVtusYeOJ
pWSiuZXF50ccj7DlpBTpeD/g3QUD6OD1lSKIfDlh6HbNJzb0Opc5bBw734pGJx3sWWx+6QbTLF9i
panN9oPFgLvab4utEGP2CRoIpzerZMG2Mm9v94Hv8x/KXSRORJqx/QFjR2CFyPVYAqKrHLGVpNYu
RF7PKTF74SAnS58d7m4voGIZ30utAYYcE61XJDe/sZ6LWfIZLuJ/Bc7GrJMg0qtOrv3ntnig10Cp
RySR5i+GQN5JnFTy9vDQepSmH59naEFHbzDSPx8FtywSDEgx32AGDtHYTolKOabLufRGDZ5XFesp
R4SSfbQ6ePMORLGaRqRuJl/EBoBO8vtrj9YOKUgH7btVZqFaqyZnbmSF27ASmPl2pooi40O5WgDG
gsiDOf9BJqo80WJPVWTef0YClnQEwpOOjUh2IAtdlrAX1iBb8f4r1MDJi011SLO+ZQ577q/0Kt1v
4kT4tUlktT5SdfQHeYlq6PI4vNNfFsEfDNLIAvMZBON6B7YQIqOonb0OtV/UdGyFvak1YZP/9jQI
jcfmaMNOoOIojVLRZcf75o1e9iET1zzN46/zM9P+LczC/58OMk8ExaoaTug4+rxWMvAqus+SIrQf
mdktOvZ4Lsh0P/00Jv3KuuLqZoIxCp+nX4p88zBxY736ft+IsIzKlHrRbc2XYdzH34LcsgsAmd8E
5SaRvKyQ2E/+eyUz7JkqEtJfG9O5Rtm+dcgjzoh1YMLG74LNt7s0Ef9fAyF3qy3IS7cZzNwlPIko
ws63/KAbmJoBZMRDSM7JPri0ZaD8O8KMRVL9sWuSligNyPoE57A6hO2aadjCu8AwI4nFJKA6nS5T
BiK3udLu7NGxh7EiHzh1Q2M7+6wWtR9mD8wCA3NeEb4p2IFNpSD8wytEPDPIABLYilqmEKrFobzh
Uaxb/MxfU9B3rd58F3oSOAq3/La9ZrAg+0c1wGH35QWeUeUiE3+eZBW5ZA0Ra/nFjOvZdZjF+xzH
wHL9lv1O7BODlHTsjR1+YyND4N12SFnxksFN/eZmgRITqsvRCKMOEalS2CCinAMY99YSOdJ57Y2m
8YzMLU7bhDghRpkScSLjlEICq7DI9KkirTM9+PuPY/8gH3Gc8jYwRkkKefVcVMTopVHtk0JfZh4t
K7C8ra2nazGYUA+lnM0eqTKY2GHmEMtUulgvrIrpsGPUq3cLUF0UPtZkPy27m2Ut8K7GOCsjPlcc
50Rmq3wHuABqSpwVuf6ccgqxf22sb68OvPJ0s1dIJ8kQkHVb6S/QsOinKrRCUlPEURPVS5D9ULx0
nO2fxAxGTwypPPaWu/UaR9fvmAP0s1yuMDB4ckRFxri1WlX4UnqNEuIvzTyvInakToE/33gLeuhE
UxhlcztNJGLoGt71f6b6XrncmNSMlsTaW9HysYwtSJ3Bp1srOreulFhHuCxsGscYUNGUz2VvruyM
UpGDUbgkeZMJuxzXpAgSNzwiSx6ur72KASmS9H7ttifqenpyiH/uIThC09hF38eg/mBfrv7ViV3T
GUasK2UshOQ1JzXZNSSTd9N9dgvkjB6oq/EWQCjyXoZS3ad0pguuRichQEvniMN8d1P56OZL+DqF
bEcgb9W/4BQpRh/aVs+DgMZb6/1r0pgjisCMxzC+lv5vHHjns7YMujNO5WDabFllNmSpKPqOSbXo
NYpFmcG0LfpBmsmNXh89yvTZuUoemliSWNeveiV/vhV7jCAxl8JtIdYeu0P7Gkg2bzZAXq2gIQ15
EbzizLPB17HZCR94ISvdFd26KixpSpGgIpejBIXadECNnOLi7D8egKMUjSDT5pmd1WuTwaS5WoKC
7dLg6U/swr/KlSuwk2uPAzexSxNVwP64qBJt3SuuPFAZLUMOTAgXju9htZrslpsS6AlLcj2nJQaQ
fZSJwGY1yXvrELtN39hrSWZyGFVSWQHST4tz29mXLzUr7dLtT/hES8DcJACVE/qY03/kt6i3hCU1
vvF08SR7DxWKWCbvpBCjRvwvgkI5V8MjumEZyD/ypRIPEfZzq8k1Rx7qHOv2yopMPULTaqaa8Q5p
sTrnNxIqOR+dSD5TdOHiyLwec9nvz7w8FCN4qHQoCxU7UBxUQMz/7ZQDK0cNZDgU0gy+v782/3vY
yIr5LKrhT+u6AXp4xR56mqzPchocr1hlKqpwh9wQ/6tRPGjsedb9i+ef7gdc52shlVGcNIfmmINT
AJzN3mwaRCzyqm/1kt7v+2AaAkgZxLNPIcjftgIC6xYVOdjbOT327IqajA52iNn/84xk6fL1WvL8
D5BiJAnJRq9EaIWNAVd259EEzC8KnTi8dU6uyHzm42G0mD9RNVUNJ50vYmRk3fguFSDc4ZBTu2X7
BcAWzBU3te4eINeAMb4qxeWHS+xzs5apR+g96ET7dZ/2aOoXzeKQGE9G4tRh4ytF0J9Pc8qJ7YK2
AvcxiKiElQPnnyRvtM9xK6yGVIludKkbAMQy+FDWxIGprKsYww+Kukol+jrFp7RqnzmzQaMM7BJQ
Lw/tVeTsKLLcs2SOcDviXFT/ud6bRq2mgfR/YOztvvwojtYsxiVmFJiaGXnmqYCvlXDLZWLwfON5
E0tPjOWrED6oFELCzj/horiXup5PW6wVH0KRgn+g1v1JhvOlnYsUDiM05MNxVe8ci4zxYMMP35yy
lnWE3tjy9YTTXnTA5OZG1RKguV04zyZV4ty7T/YHNZYivalv3l+NYEnnA03OBKGJ3+zZ6haYdFai
Xv+dcVg2ahEQ6xz1zDT6aNJO4yeiKK5Of+Pjk2GqQJtLruxgrTMMVNB4rL7dtOS5TDrpCNRCXw8L
Iv5Dm9RxuJ1CySTwR74gun0yU90Ujab9ZCVMiVaAvljUQzShL50nwd+dkI9n6sDhLbJGuX2N8wQf
F6/z5u8hB1dKkcSdU51IqnsmMY7vajhkDtdc2LgpwD9irVwTsaE/nXEoHf8tWu09YG7yRIidklJ3
qgpLFtpU2Lc+IKr7Gb41jQoGRKPBGhcUc7bqd1hfOLHDapLANwKU5pACuWGT6H1tFrweTgN+J/fC
Gue1xuj6XBo2czHKhFa4EwjLrECoPJAPrQvcL+1PXepuFCdE6FEXdVbD69G8t1HUQqBej7AVA6+H
RTFo7dsqLBaWpj18tOUM+lO1UBo/RAlqiXhxWYJSxjP3MitlwhNfd44YDKr3T4pVixI46JGCWrd8
VqmKqtp1uakdp7U/seCzcL264DiTdq4xy2aNgL9vRWcqRmiSfxXVeWhPrQQbjDJ+nSc+wlv/ABhU
jrbQ49eduRzZ55ji1/CaBo4ubX6pJQJymKFcRUTwwZCJqSHXkhz8RIjo/8gP+1VoM5AYkVF0naGC
uQdHyMKp4KNpIHcg6qf5tb1HiBgszDt1dwg28tJ32GgXli14oo9p0Ffvv38IHRyi30iJmzjBdmgQ
1lv/Z/1LkEiff7js4Brl4+7Q0SAHPRclh62Bz+pAwdr54ECmxpdWfJtjttbzhD1rQm9B14SXlnos
X1zObEY0/Q9tlyi33dDBJ/mimeuOIDjJkx4lCwqrfHmj7A/6Cb6w76YgjZmFkhnLtTt/8KAj+9WT
QGnIYsk6qnSTsG5rxwNEx5TZxvUnVjDo0xaZGYXyYI90ctEvB0KwBJT+GXj9xS2J5oYOMTnBgxsj
F0+bbdA23hYU/97oECRClQ8XsnPCIy7F6hRCMGFKJF16qmYtJ2ARQJ9sJQ5wrBbpdcCQiLU3vJWQ
LFzP0jC4BIErds6rq5LPpXRUehZF/sItkZSMuOi2pnWJPdklZEfOeTHwBKB8FfbO9RBeS6c4K6MD
wvIwp97zlWkoYbktFGZM94G03c27qVGl53DgtTn5oeLK+kdKak4E4Y4Spbm82/L40/2xvPC0RWA2
nUZDe691PdMtfImKNTfGH3vegrJ3fhvPCatDQA7EtVI2doq4iqagZGupxTNNm1pYI2+PkjOkP6NY
+rb1AftPgzCFJoj7BrmsPJ6OMDKgkpNew3l9BkQPlV6jVoliDGtE9Cg6m6r+B9TcrJG/40q/NCfN
copVyXZ7P0sPxqtV23TEZ6/uOf+gKudguBCQtwVFiJvNHbrd9Br9jwYb5zDNSXxx+y07P8dmTZ8c
jWGi25DX8RCcV8ohr5HH+aFw5/PXKkVu8qUwxct6WUlS5Y9VyJqHIk3Bha/NgTnXXFgn+RdYLPJA
bAGGz4fsWuZDLTHGP6RD+o2i81XOcIHXMWS/uMb4V0HG28DHMhnv+r6IqBsrQ164jFMCxyr9kZkk
u+DDQE0dQIveFyCbM/OSPoc2f58efyiyxQ3DuQXGAdlPFp1Lo7+X3JP4acZTBS/YU4bYBUl5LAMj
uH573kBq6AUlafRYiL7B8mLkmMtQpDoQL/fh9y1OyH/b2yEbKRZO4Prmgg5ZB0C/GcuQrbeHNXZ+
Whg6z1q1l/SV++hXTc3lO7LTtp6TCa0CycBFs8EHcIN/IPlrRetyYAPMQsE7KDYTtqkX/7sRF0HO
Nbq7oKM4dZmJ7FAj6JXlafRo/H4jFv3nzNlPVX8F6XyupJ+ElTSSi1p7cHERKzXpsSpgcKshlSqy
9J2QPdoRvLSNivMJVcB98Y0F15uMTZSymFza9HiOf49tzrAuwXwTTuGFB8SB5bFgySkm9tyZ2XBk
wj271pe+bylijXK+4z2ULoN4FqDRKKJBFTNOaL3nTWLc7+5s1noCFA7fvbGOz6th81K+be+P3TAE
efvxawDhQwlrgrOSeJuk4K2YEnPnJ0rChMTp0IwBzhwdn4dCtb0MF+3zJlACpugUTDGPiQW7Fm4j
SHh42GQzo+olefQ+idpMc7dwEP57yZIU+KktY650/bZFPJ+Jmf19p8/bIaFyuKubrr6n+T0ZkB9s
0A89xII0zlUi45tk7o18XBTxl4ayVd7hctSoIuTjx029l9K/K5+SEnAVQaL/CxkaV5jYrov4iHNs
7Y+ZvYOtYcb5ouVcGv/vtTcaWsShYqJwCkaZi+xHyl7HJyh15GCnxU3tmCIFqFVzSFOkHcQGKByr
Gr0+jiqLMtbS/kitRuW+HFA8W3rrH2jhJ+1erzXOZeyNuwubmBpNwYfTaGj+dLbIFf9cPePODH2B
yGK0nNzU0VSrpEyCzL2LbNWceoXB2TqYmhlhuFysoVB9/sUO+EpppfeEnW+vMTUq1+cmQCdx7Rrv
iIH7Ie9RaRSW15dB3AyoqE8rDm5Pei15x/BcsAZvAwhqr0xwKqfSkqxq4QQxI0HHITIzI9VxqC0L
WUmwLOSe8jXw+AHQLDbxO31vxb9xFbm9GiBkpQfMnEjkxAPkwhXTU/IIvjTpEAWdSos0gJh6VBn2
TuptV4+Rfswm7HWuKpno/NdmL9EAWvoeheeTygmemAwrm2dkodGIUWP54qSD8YvHBiz/LPQIsKRt
EOO+byFo1qaHOQq9tltfvxxWtBzgpKWnxNVjhhedW9qTFqzkEgioiryvBpJzkqdDSKabC7TyMKQU
AjHVCDqvEm5Rw5AeNjCq0kcT3k+QPeCxCRhPg848JmAr/d8LgscREEfMy+zTiaKVNZziYbyZqdmp
zY4GM4iqhfO4BJ5yEqFXMx2Wb20Dk1zylnE6VY25qdJH5bGrsnPOV0bNCauwBy+roouO2y+bTrjh
z5+0veWEFZV6KUXihPFNn4KXGbT6D66/rXvnllCXfDex9yoMNi/JR1HRTfyO9eH+J15MSzZ0h3xU
qd75UGTdVBdOYbZREgNf+5rhpGFZqJFE/UsG7Eq/2x5nrEKpAPxyPQM0pUEeOk4c+4smSQiA46Ll
FG1i6BAJo0vfJzl+Is0YDoE/34rxHgHuRbkUZqKDlpU9Q7hScepnwINe8DPBYnANtBSams1Gmu+w
Km90MC9EpCRZoYr6DRky7rwS+GnEFp112ZDqQ9JIW29+XegAiaXdHZDomy9H26zHVf/3wPNnlw1C
8ZPPb7se3VZmBVHEmV7hw0TittitV9jk7OjYsW2CEecrT5UfQJknjLQQrCw0OwXmu8reUb1e4guK
QXo17I3WwUms2ol1eHf3G312LygXfxKGsee9ibColeQcZEQYuVojXvRGKkMIzavgRfFu8ZHA42sD
AH4XEeYKybd/7WN4xP7D6AWSi07nsAwfNHrH0/YmdWM10KJE1PNsBIqQdMum1pqC/KLYaBUCteJq
v4lO0BAXIXnH53xvgrtZlMD5uODBHYQKOzqSboTHLvltcs448lmRFWjG7mYl9wLUtzN4gOyo/mrX
raJBHs05w8dcF7mQg6B1OsdN2Sk+Oebh4Dg8Op0e2oUhfgXyRLzhsRe23peeoyja/KFG7WEF6D0r
ktlGQXVV+Za38F5lUyyXjRc6NdNEnKI9D/BeXgLPSXWUPPcblTSnzOLrD0wAXcHm37Mt5LOvbm5h
tNmfnH890CziL7yCVnaYlO9DsAeLycdquedOyoxpBbnruvzef1B+eobQlYR/++yjsm1Kx1LfOe5w
EaUcNk0Js3OMs2e5BjtDlQj8uKz27ec49u+51nyYPEaQek1x1+fs2CVkIZZEkCVtzWWObJWKAVuD
4PHo/1azgo2/fOhibaLf/PeNEyHtor4xieLRnVbzdejBa3dfMyLJPBmZYnolTwsA0JijCS1wwge8
tOT1/IUnPk0Z5HhxUh/iLzeS5dlKYT7vJAucK3OUZDB6OcVwg3CGBEf3OJLS7A3YhIqNgmBcy4/A
oZ2+PtgZQkYNCyBnHiZnwzyPTvkWH9qX9GHM12BWhhzVz0Xpr24CDVOep9tU3W3NDJ1mgXFq7Mcw
5pD8lUF3dK18KLmHuDHkjQK7S81nxDrx+rohg/QYhmpvhCNWEnRT9E0aH9XDPJ4YLpd0fncapP7k
8Udg7sIOUK2z5SrtBk6Nv4q9GhMZ5ouyU3qp+pLzOGrDX/CJN5F66U6wMHEzlZJSX/qkpmDkEolv
LfPKVBbEF37GKxnp9pDhVuTURQhrQqwVdunoylu5cfdxhVal6uyJZ1J3YVTZbAHZht/NggKcFvpI
4ZPhVv4Z7M5ZJfXWvR+f4ZGnxrWYES1Nrxn+a8TW+6Pn8x8CTxcvm5rofbLGjdqVf7JHI+sma0AH
0dSuxylfQIegcbfTq7ZLPSK3iwOc8YeObr72Emk56nxCXLzNlIUGSllBJVS5JtHgjptVJs1x5zbZ
owAddEcio7dPxM2Lr5mKtG1YWwMHoTAp1UGBYkdTi7m/Hf6++aTU9sXyxJxwNU55SY5RGyYHUzcB
wUqqAxaxGpuVyPRFlPYmeP8fOrjiFL/tnb08fphiRv6UmbPycwKaTnL53pg8RM98o2Oy5OCG9UiA
pXva9sfNMuVEaXYHtUNY7YiXQTMNzNe6GR2kluAuVj7K59E7E9Jz30TkuN/LnAQftBUT9gFU5boC
7inWrfVe6mEOdgdi9ai+vz8Q9MxDtc0Nlv5myDz4hFPWkMTt/QKHd8TnXKUjdRgJv8j+Dx8EALWM
R0kKgYwhVooVSXhgEqwKCkk9YKi99tklbPQFeGj6tsKued20xXrWzuiCzZih0kfCcFHizp0a4YqF
Fe3NnzuNskOZssdmzEJwbiMKg/IgPcYiuoX7jLnJ3I7P0IA31RSajeRaR6OSflNHxylvFPS+Mdno
/c5bWcXYRDwhwSf/ub/a9UyzsIrfnPkZQA4J4bwS2HZ2yhqh7X+HjTJs/nqKAXhbNBpTTqbENPDK
O50Cmg67FfhiNs32BP2jDjugaKzliomEa5jLQMM9btjRvwO5qnyvc+HzkTxmGQoKGtpgjc+xxXP9
ovBHVTyWDV8b6cxv/saNxo55NYpXFYuFtAIC8omFTL4LJtnEzdOw251GbpIrXLDxTKMyHjXC590J
7OBPBjDFVQL1u03FfUXHeQwgoQTuIuPIAF1J8ALEuoxAj7DoeW75zvOGyMeI6QsswGqZpq8rYR04
N8rgy4yvgkjyFvQwDJ2lEXcnJRfR2/3b22qrvruJnwd91CDFQt9AkXAmCIPwofw+YdZasfZoAoWx
d18i+TseE1jFkJReL25hGAOWA1KdWmIEkapzetV8yST2XVWU+0eVhbENhEYhMk3yWU1zs+XkVNOJ
pELBph65/8Ecx1Z5kr3+knC7zpiN6z02IhHBdct5hg==
`protect end_protected

