

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
I93D9zAOqgF5xhkIGPbl8GJra4lNAzUCqWqwUKHPRswLTMNB7+TgCn7D1jE7gWMcbnC9BUv3Mx9K
oaTY5ZseRw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QQKJOb6VFqqG77ztBROe9vAN4TIbb3YHpw7kgu/5jUIhCNPRlaQFxoG042Pe8wBygZJ7zZGLaMks
3B9y5MKz2IimhFvAAL4rqgQZ531fkS5xfSsbWqEpJ9FjQmAFMtHZJ6pyshLoql+rjOPMO986R9Ul
mCT+rwL+hUXiJFoF/X0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ULN6geEV5Nx5kceSmM9wvqfbf++hx0u6GVwH0ft4GQVO7fcMuhUWu+U5R2VaMC8c/ZnwPFC1TwXE
0HFdjBw/2TJT2r6RmqFwEljM6I7iAM0ScDmRYoSSXBENvwqHI0goYU/SAGW6+xDnhWSgaZ9NbXt3
l48DQ5iRhe5lA4ct3wDZ+XO5oz4idq5yrKf93QPFS5A6rlNWPLnA1a4ATeIcDAdlg7MAdNn0si8G
h0IlfCsnk0X+fjYzQ7Uek2spxfDgGcNKcMorlJ9jhRuuKPISwkTsJo+lx4a/4HBjR5157XWRsO2g
9ZI4ZmM6VXmODBYy7xEmACJk1RYa9MaaqHjLqw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UrRVVRcmL6e2jhJjoDrNfIr+b2UsaitDs1463qkIPPDX0gZHSkG+EGUBF7zxh8t58vFY4bRd4zOQ
paHNUAu7UOx0cjQFieL+Hfl4TPDGpcnCXZeWSwFqFHxoTJmhwWCdL1ejkVLE9J73pomraPvva0nh
xNx9s+ng96T2SsqWeXntjVlSNgQhfajKj+oGmZfy+XS4v2Lzowyo1xZkAl6c+c8PoAhYd3ffwwIy
KP48nKcw4RX3zRDxLuiPyrdl6tcny1hIpuSw1OJn3jk18XT8E7Gm+K9vzhWM4GUDyPbM3oJBLuto
z0HKNj9a0nNztwlvfdtk6LdP2SPupPvbHpu1Tg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V2R5QkNtdP2r3qCMkHPuk5SL3rXpOUln4kmMrWXT6PzvlAB6j1k+M8OLBhMQki9X3e3j9BOl10qV
wqN0GBAajVoSc3rI8fh68LiFGrH3sHUiF1nFXSuBtP4x/K8PP4hpEdQv7NQRmPKufOOfKKiZ+4yG
PaifKxzBQRFRnzJlqA/BiEB8zeMzgjk7EFxlwEqsStVOA2RDDUbcD4uUM5c1z2EvO4lDmkaAqfTB
n3xASzgIaoIWDW/uUdMxbCIazQpE1qKHsob2Jk6vWnhykaV5mHiW8ybndPtiWbia7YYcHTT7IAI6
2DWeLpSoe/Ja3FoCG4IsukXOb/pgo4sdn7GyKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fsLjVl42s27fKDlNsuViqofNZWdDeIYLgav9sjU9dBfXdmwtLko79oBgFYKuuhAsD+2s+lxKpn+2
zVT74MvgYH+EnGZU9TSpgR74YdtZfvM+yf9sVHAbYRfX7euNP/HhqxUb7DwydlCEeYp8JpVf/jB9
IbGzhm1CjlZXLIQ6z0M=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JuW5jal4WpNHeWpOjtgpJFIASjjcUEPZ5TZN7t35dvLYKTzyvP7E6C8Afrfg+gWYO2Q4ZEeeo5hp
qQ7vLWjxQKGGcWI3jWcbqry5wNiQ2BSFIw8cgAxr6uXR/dPKcKJSdSJpsDUA5QnSDS3rQfGN21If
41fSkewwZK79CEsm1wzDE2+n6+4ZPHB6x1LZ3YMvjCo3yu9UJ54k6S0w6ECfxiyTgSoQ++rrIFxg
DyJ/fYmTZM+6jsvM30MDw5wX+7jezHaAkGBZZ3KiIXiuaVNlCp92JzroAUqBV1CD9YjeuFS86pOG
CG6HyTo4aiC8ej1jIcTj4xnPiAqrHY5CI9Jwqw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x00J6OaKyc7R9A04ctRfw2tpES4TJRjYemxLPGwNgVC7tQtzFFSpQvV1uu7MbHc/CbkHQQm0on+b
F/ZwLIDGgUhVBsG7bijWO08tIELcW4pKhrCHjH42xxueIezl1f/AQeWjafSvZMUc+TqGLDYHD+UX
E2T18ZKQcelTfU1n/wGtEqhJIK8hgD1hjbufk7XTlHZGiaI46U9LnGuslGX58RxUeyE6D1sfW0fo
KWr7KaqlcLpaqgIC1T7zJ6HwBjQKA76/Akfy+bCIp3fygfUHd1cVkl1pmqTD7zDbFfvVwpT/dBql
JIXQ2pM9Y3TLo9gJsCU4zm9O0vjgaacKQcewtQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 719600)
`protect data_block
o+axQg+fZOIzrU3FldSdH2DDMM4rejjs38bfZ2hPjudKO5HKHBoSUOmO4dXRmFnIbiLWe+CnHMJ1
fLahgEhDUDImRHY1GCem0z1qq3k0ZyAwoQ/uPFt9CZAapJ11MyAFaDL/rusd/zaYBMdNjLUGZTo+
LFvM64RYBIZ/vp6DxLBqTRUQ7Bmthkcbw+oJCPu7MH0eVdse5uy3Gt3k82fpr4HpIqW2apfNoErZ
JYHPKQfURpdPv14kkJZx62QAUeQCvWbzh5LV65DdkSsLosxCNYYHlCcMwY/yuEH7FQkBI5phtPEk
+PkcQMiD9v2c8DdXKl1yG1wpceqwKOGZVnZctaBH8oF9e9XZEc7OHV7wJOY0tmlWktKldsQWnpj2
o9SQVGGuz+Foq46MiL0nya8ZXU4Xp7HpO4Tw60VbwDqTGR9RsCR8nyj7qHkn1wk3kdROHz2rnU7b
m/yJpO6Wjl5eYE1Ff5hMIMAjLBClwx3hnL6v7VMaDltCglBv7kIZIm30020I7K7K/9qJEBf4Le1O
yEWPWKt66H9yYaa9lVGH0iRfzD1Qyn0A2Zedx1NHm4wC5+XzPNF0SFX/iZwyjGp4fEKGoM9zaGKp
yzT4GP7TY2KS8eQkN658wCYhA2mTkjuQnWCJVAa6A9XAd6fZy5CYLff+eH6Xb6QN7H78jLL5sbOy
J/fvdG+JVT/OoAArQ18/4d09Fa8UdlR6hhxUbQN896B3khPwY+T0IqKYJVZGGU/lMVQZdYk/EqWo
MxKZelo0AAGFCIG947vxZsua6s8rSDZd2Vk7g85pj4GPX9T+j0EVLQxcgp5HXpImsUOufUI3SKTy
SXuzCTYovZ2Odk0EJ9yzxhQDREajfFw7L6kBegov2ESESQ1QoIXMyHbrtHNU77abpZr1b9dgybZ4
3uZLBvNl6AKotn0A+pJDgie3cegALGRhKBpCAqLmk4J6JvXm7ICYbBfGuFJua8+42ZX5PzzerPYZ
jWUrirIvTJJ7ViXSYIVu1ZArvQqUzeQz4YnJLMigIs/X7H6F2oFNTm4n19avWjFcwRGgLEBprcpr
H1WiEL3Q/AShxUew263wSu/gglTNmMwTEAu0e02TvlVByxrupa9nrh3oMKaKVEK7EsW2iVKOrXws
C9s+ex21nq9VOV/v45PxVHBOJAgmSG2hO7cq3DtYGLGZUyk6o80E6VreTjLvuL301FteuTBRboiI
0aTJVldJWic2Io8jiqN4NlQCMHmm1oERaK9ndb3DUvLbbSLbuGwp6r1wVmlfrqNYGyHSs3OXvXeM
Sf6neywdhgWbHD7RN47lDaM7CYwOmhTORXbyGqqCVetrT/vXdkNEghe1yrVciQ53AZO1LCwiyKc0
PCzNN9Zm9f5iXh0gYE75MpwjPTtOEGUSi+SMNPSaRXXYiwAJi/4UYsiTPDf/OSJe9SEe+BIctAZf
zRA0DTi5QJY8bm4CwXAuZQ5owPHEpk3fkVtvVdOTXdFRQgEthZ5LG2576/ofj2RGDje2gyVLW+kN
ZXqID52f/qHLFD6PW+jfqUkX3MVVeMtzAvAlhmuRsjNa1+AIy1ecK8pLhOQsXj/McU8VgwVoCi2y
I+c4zO6eDtBJwKUPiRTBMcTi0N9xXve/VaN+SPlUZ/BHGv5xuB5ahkBrNlslJWXfBlus8DIutMRx
BBY4GPAP7D1B6i4hbBwLs0I6zz+J2Y70c4bzkKyB4ncdroKzBdvJo5beODDEsxtjN23mWpZ6KTaH
xS6BGkVncxR2yE4TW2PvXgW7+MAGELEawJZW4nuXKh5Y5u1AMpsBxEGA+ca8hLpxylxna5KkRRdP
1XuiJKtvAy1x5Q5BN7HV4BTg+lHLn0LtRVPptrQtH1grOLqmDVb/t5oEl1bRxiczpd9sECKbQ9Nt
ChKyCNRbKByOpHfojGQCvPCLUcoUD518BZwLm0r9HcClWDSEFe4IPOz+gRqG5wFtMpbYj1f6UsM+
dL/7Q4vbnAnnYNhfUaOHWtmPwOeDYnd9Cp33iQC7eKZ32uMVOLi9F5QgYh27KFpSRILg2gymXsY/
LpjxyYAcmnMU5SlHVEiD/KAkVqF0iLvTdGeLJkKtsmFHCdwNgaVzGMMG7jvfLv6VEA0hnjFw3mMD
HRA9eWz7xpTH542280sB7NW3arxEYqQjs3JWn6R3JGIXK8Am5wVzjK7lWgB7MBlpOBK/sB28Ipcv
Wag2RA8OhOYy00sfN+UuNHNQLG0sh+I6LsP3nyt/HuYCFUqL/fZuWeziwFiv2qLBi9/dMzDg7irC
0dN266MpQh8Yr/M4pN+DQReOr3JEvw8FmffXA3zUZaStxmIW94hKyIrBFVcM/RVkPZtGeJB2mOCv
H6u1EmExncdX9WE3qwNvYuWP0aO7pqG64jWAyHmzhHCgQIJ0Vh/BfHwwp3elML9vWgIkE3BFewOS
1kNIgznCxmtRFb7k/PNeIQ5sNHwEfp7T/cobIua3XDMfXkQPMjpfindhcJz4F0p/5xxSikuYOlag
1tHOwF2AVzvMSw9DFbX2xvqrZrGD3dtNU0CBJJafBt5T/OS6pOKY+1bqZpeDbQwXPdjcmbjs4Vo9
Jxhw6k3cgoPxKMTMkEjMeyAWtZoigt5Pd2VEhuhNzOQ1AH8FaMfRguggTiSCWmCZZtedcnQfM339
GvqWjzAVJGRgHZA3H87E71eIa8sf5dWF/ojjDs/cHP/4lFIbaSl+fAjwJPRiRXlik/V30rCE/r4W
y1RTHVHZBleuqh76+JSnIT0b+6V3Xbi8ExhRHi/ljxibFb4XLxwnczw+zhmJ+GnPsA6HJPGC+pnQ
4Uc2Xxq60aW6V8FHKbS41k2bEXfmy2halqu/6CzkORcT9pXJQA1lugrFG5s+hrIN6TBKZ13jsNmD
PKP693uLVZ5zwTlPqCP83bL3C6dwD0qhVX3Yz+XFE67ZYRVvQbnJ0DbyppezgnnhW82EVCy9reN7
Ulby9lHX0mfZ9Led1znAugH/+3M2PlV7quwteojpQLK51qZck/vnnwdlpS8Z0+XQjmyKWw3p+NWY
jf3OvOuARA5On+QKRTgUG7lxi/v/Aj8VAErvOlGJ+QV15TlVzj2dJ2ZGUp7S9gRBmOL1CDDWwIl6
4UQF0Pky25aVv+DTyQgJ7ksu32i+276uDDzi2SnvyFU9d6l10D/Obt+LWBj7QrmBRVNJWtGQjhs+
iECK05MZQY/kobnR3kPULCDpzrNfuDyTrhoNRZWnnlGB7CyRcnbChReH5DJ9d9hAQI2EzatKH/f1
XPbjdcDNbwTrvWN+uL5wYwMC4HWQoccnaJhBkMbNkKEKgPxfRqRcez8w4At6UCzQMwRWwP+xRCZm
qQA9ai9Qtftt6+cbKuOBxxVQLeEet4/E1S5WWrgoDc1v4j5NPAcBmH36e2ZNxhAgSKZYUeQ7fMIb
h73Vccee//qn1zz/OhhO7sMY3UNawlMCeJYUaaTQSCqXydUdd2axAOG+/fKnA1ZI9+oqPz3MK3fd
/6IB8WnCS3mLQQCDIKbyHW9QFbcprW47T94rzIIl9EUiXEGqQsXPtZ0zoRJxJtyT2qg54zFCDbMR
ITLcFmeuyuIOqRUw8O9AErBVw4YedCB0OaHl5h/gC8D5dnjP4e7zF6CvpmrP1VmsF1QXQFoSZRya
cguPanHLi0BnQnkL+5LH/GG/So+DsGbbx1tJ6m96klw/4inKjf9mP7iZEMGg5DYX+eLLHHFlIqlm
RcmuZuRfSjZM743gVMB9EI4uFyjFPhutlwGNWmTuWR0Ote/Iujy1v+rCfz/fTxR8JlmShU3hPSw2
dP5GtqOo/lO1Vq4IaZrfBizYQR5OFnje1ravP3JgOjOBURzSNJA2VI1oxeA6pdMk2z3PGVkjt8D5
YbJR3J50874uH3Pt3ecg/DA1k4Vtus8mI7UznhIP2Vvs97GoPNy4cd7dVm5V0LgQPNjzxke3V3Va
HBqleIA/pKn34JD7qtqDkScKtdUz/ZPeGVuI2vQGuFFsAqPtKlY9wMwe7rb1KX4GlR/RXSovvis9
+XE614tfRBpXTSNIbGIUx557o6Zkpk+ZTBxkXmVmyJJxCuib39n6ulMRpjM62bncrHY/EEGe01C3
vD9EFkoa+YSg8pI5NEVvVIC233RBvG7gzhU7UfIISNECat/NNFqXL7NWMcDE0dBJNcLLXxodzhyn
H3sXlrZ+69aTXkbQRoO5vllpR34AC0PG1YWpK4cU99NnXbySL78pL9ZUBcuLM1wTBTEjylmyT6JX
hIF3wGLtG1aK4ypXgMfL/tzls6q2CjF6WzKbE8PdS7A7vRvOidmfwN5Wmlta4SQ9D3/9Khg0Gz+A
Ppy0JZJEDOsSQP43U3mUZc9HoasxJrlW4q2vq0q+jxnEcjnC1fZKLUCXh1WAyaJXYqZW8wIyrwfr
60JL9W2zWaS2xGbbjLaz5LRb8BhWG6l3IYXyWZaYcUndV42DNcynlT+1kcwIj+jj3BIkuXhOe7LI
GANxDbibGkPy5urfeGD/tiD9bWK7pbbIZw1zp3ZTgswqeYqCvx6uY4+pr6zhPmtlaahSp3qkpNN/
hRG5GIcNaOpMzqVWSuUUBp9hQQ6RREYON9A9R2Q13yGsXv3zhARlXJN+Sut/IAtaRdEDmZuxCgNh
HzZ6A3CrJIsw5lIlzNwKNWpntH3RYAFS32JE25dS/bz0TaL4VWfKzrhn5oL9Y4w5D76BWDgOsqoN
ja4KjJJs70GJkV2SCMo9BAlaAuimBYn/HbatsPm2oXwZm96dElHrsA+TvUSz3fzXZBKXMkit6v4X
Z8WYsXKS7KPsEfZpGlCeVR4pDJz5bK+l7ndyWogf1LjdLnOoDHk8QGG+bV+QvttWoe+QvdjKASWu
hClSeetQ44wSC3pu3cLSBZG4PC94NuwZuHw5121er2F4jbIULzVNz8ma/x7oxnJIWp/14cnsgSoY
M8pz+J/loAQiwToDKnohEW8+3RpMZ4g6tkm2rsmLwEMuLP5TZ90CjOmqfwICBYqBCUG1tvOpfPL2
v5leFDENea7krc6XDn31aJQyRy+g9aWw+hx6JlG6P+e1fUzCz6w+TTtpOrn87Dz14AaP4X1Lu38v
Q+nWpotVnkisymj+n1hu9Hvz0UficHJWSSv5W0LO0DV+lg4zU8uUjK35ymvvP75G9w8Y4X8He+bv
FAFJ6nYHJiHK61VyZRitcwg0admV3MXW357HxN4pmEvfKM96tQt0y21KiDLDn0lzGKx/mH4K4V1e
zHsL5P2ovSAXrSNBhaLxCwQcFU2CnOHP8myiwR7WJtz6IT5sCVUY6HYHbPExNajthF6UwlrkawtN
nsDZdRBFDZARAze6EU5kK+cOv3lTWnqRP6RTFAh8rA8v2Zg+sTVQzI2TIyRnF1leKMA83h8LOkLy
3Xf8Eku/ILUaly2hwVp5e/asj0iE0N4Iss65WBPrb5+SobPEHlmSSdyuj6F/bnG3uPvH1RtCAIYA
ofu6c8C/Nq6R/5vYxLvwOZkKrN7LpZinL4DTt/65WcOX5gg5kRVxO9M57QNML20nvEg/WFJ6F/ED
AmuxeTg4DlbYvQhHyl/5PlLeSj2Gmkf06OoSijjzxqASs0COSKzPqG2C3UHc0Va/TKrgKimncCrj
0H5c31W4VRARKJnyWk2t5M/ZGnrQ2KGEDk8u5f3LSPKCkfUjUwjhvkpbkDV4ebLYVaj/lQZmLLSR
YF/KOEhPHQI9w/2Wj1jCSxcoa2fEsOm5tp7EtpocET31BvkNcqRTPEiY8DDnhuEr2Z4s7FlLIQj+
g4GXILZTjEQMXffFaYALllGQQTNSjpKB60qNww9y5kcafIL4hiCj6TpKWnFyYXGeC3vuvqz7ETNC
YbzYqsm8zgF44fVowZ380LYFrXa72cJj21HYO1fuAFPLSbbE42ydlXb3Qobeq/l8XMCCimJu0DAD
Dxk/DpGjCQgeNFb7rka7X1O9o+Gpd5ESDVTUkMuMKpEaB0INR5/hZ+grQi+46QS/9SjfqflEwxvT
bBYRvsccri9yD4H09qQAFa9k+BMcFyL0ukC4v8tPlPNDWkpHh0ogXXRwxDDVhqRCCX8zUt7NqYNM
JwUkI7jfff/ODDRtlTLNJcrGWVlbMkZEsTR2nr6tc56VvfEOPY21xbqrAeSC7IW9S5eBVMb5nmHT
UQOjWRDbb0PVLb3BoRdQG/qReJNLVe+LqFe6mx6raCJ4MVNlReD5jn1ilY06DG2EgK9Pcd4lqt4m
fUaKrx5p/Tpg6ouEUzm8/c3mPNBvjVZjwHcep28x6Xy2Gc+zUsZFLyaw1B8AFtAluay/U0kbPFOb
kbeIVVBu2FyY9+chd2EQzZLnilSac3BODyPcBLQOq2XKPE9n2h0d8wZ8II8IFMP5derY9n/66fbi
4EuX1cCbYukoAf+3qxmKWiNr7JU+55iSm2A5vf7CKEsYgxywYziW58nKafNFilVz8MzeehD026vR
mrnFIvdXOVg62NaBO7GrEnhafCDCh8gHMJJUIzV9ZYkRCvYnIlOFO69Yh+SVkkdli76Rj8vV0ery
i1enTKYDGQQDKsrPUs4uzmGbpFiYT1u3jKuGdOBD51inImSK3JoXx3JdbpoxkAwHtgMUp31TIoUF
gfj61SfUWgSdjelSDjD0o0nnpiQSc68vdLjwAIywqLvjkphy+Dx499vKseWHdgi/jzUFbb18Y+ou
+qICcBs94kQlmNlkby/LVXrK37xKXZLFsSxQExOK1ucI8vkkwb6fPiZSFCiBJB7SqarDNlES7sFb
YAr8vw2LwKH0FtX56X3n60s520EFNg/46J0zkv3yOQws49Edwcx/3iLmtJboWL81eG1VuSU4vU4V
KIJizKO4i+nDI1kxI3YYlsLQxrNviTcku7NnelVkvUDyg9tpnzjHrwWMtuy3OevxZopCRE8upWEx
I8QCybQSgNRIY/Lcqj1SUGy5V1Ka8wqpxlN3afaVMslPQNuAgZWCFld4T0ATUMdMlVhbpzzwHlpf
5m/luP+cC2mp4jr3OLKZ8rsJlwYFFxoI8NIbjQjIQv9gqOtNgumjjZHsJhVnaKwtSOkP0jldWpzE
wOBWa9bzTmu0RjVX5UjFiKwMvkUC4fDoQ6KjOPT35N1BkHBd8fNl0kvLE+I3FMhsgcrn7Rl6tzsZ
N9EH7yaOVHrEJlsqDIqJ6oqQkqQlcTxJZLdg7LhaG2fQ8QxExkMVPE6TyfK1KLjxIq4M1YN0iAsT
xdzEjg/ofGNd1IWyw9oy1VwU7LdVB6BiwwKPs34BIm4+yIbQ1Hw6vhJlRJlC1tddH0xFnLIlenwR
S6nHQV0SUtLEjRSMgcNeRZTK/KJDj4Uf4k0t3BsYtf77uZLZOEZ5jl1BpMALBJgphHc1WYskWvfT
z1k82Yt47IEuGUukvWtrEtNO+du9KXWdJSwJB8CfV0i5KAYbiFRNc8kzneEPKV2KiILNJPc+HuVk
W8NqAvGkJZHElk9R0D60pAIL1BY3ufb8DvSzEiPlLBpISDBRkD+875jvaltJlKgBUjKAn3kf79QA
Vm0QNlvqR3XLYbewTktgJYMibtfG3/Hs10YxZ0/Pggr/6X3mXhXOTvpT5IVFVgTNzIrQzkY5ogms
8695kWXwYmWynQ6mTsWgvOZSvbiIhfc/NTA3307iWiQCE9SeLGcMXzkPsJkYt8HPrAOFb4sn5Y7M
1bsIQRLr2VDTux7ybq+mR+BxCtO1MWg2/GojPgV+tJaqzwt0xrceI1mzTfjDYcpj2N1200oZj4qh
j8Juox58vmrvPHlsQPK2oY/F7XFOwNwCAzlxST0mNKz8XGDjWuh7XLIMdVwEwxDsGZ2uTjM7U3Wi
ItABCf46ELmaEOGE8Ly0JtEjfSvcMI/3Jm0N8w4QDRZYUT8KYbrcRGZebABJcNU6wVl5UDbL0/yG
sh1lyTgwvc0hyemGCid1TCP+GdGURUECtRmWc8EUZRb0ni+00tb5UEa/sfBt9u5EsUzkOP5uCxu+
IdYtU1m6vgSkAMgJaI/IMb9d9rKeZWrS7wOidapzR6UKt68ZvliiUiBTCl1JnKwKsW4TgA5PYNLU
FyJt2cyd6hnb5LF/OEgASZpbGrkuATxcw/l9gjFAM9z3oaN1qktRk6H6KokPbnoOQDTnWULYybXG
jirvOen4i0gK0suYwwIKpD0hmUgubb0oJ8alR6TvOuyiSRYZpjSKj12h+gQUQJz4Vs2i6VT04h9J
yFA/P//0vFu7pNFj1+biLx+rWgho5Uv50Dprgi431YgViLoaPVMZeLe8QFr67Y//DrSNLnj1sKLx
t/wg0GE72c3HjGKVuKmtw3FkJTlSsicNlACkC8Nk36rWQoEBRyovkxg6Z4eXMPI+KnYDZ25jfwJ4
V+WZXtdbg0FYDqMb7R7hoLHDaL1P5a44L1vIwGcqT2JyK6vLWleeTdn230yJ+NGCeEbDKZCko+Tg
ekG+gEihyZjA61hkhNbrixkKLP94zsmmbnN8mfS0kQWBL4a+2xRxyc3ZBjKNCxvkRmonAv+SKeIw
WTy832GXZ2Sphdlqk274YIczijDyFeTUiZjZzLrRZk0gemkCySunoFfu1MOPXgKu1zcDvxhu3aWp
DMzPmmgNJ/CK5hi4tWxcyiWLU1JKje21alwrStSupnk4TrYBsxAzykdd1TwC+ilkGgN6K3en0E3L
W0LIb6yYaqXqctj6ripdQDvyjF3Z+pLymzJRQRBU/Fv515+/G3wesBDoiBUp+bMOHP9lyLeSqoV4
4+sVhbEk3bO91GatUHYVf/RpN4hK5cEcet8bkR4WaM42qyzs+X331sxjjAEcOryx8AimeYrx6xYU
flweoiip47K4fre/3fsRC0zDHoxiDvQI4ux3nPWaWcnOpDHTfFLNOE/SJinKHc/r28y0rHpckR+o
fSNo8v8HiWdrD5wfLCgA07E6uq70IBH5N2pRdfbEAeiWGrbDPLmyYRdtA5yCeoDa806LWXPeZDBX
MQtLbFe6c7/A0gtrLsb2tT7DPwP9yrq93KOpW9vrQ8SYidIpnIjptvsCRd9X7v8JQN/t8nwAe+nT
f9+bdTZ9HXXNVjbbooF/hFJ3MXpDJmMxJYCLFYsvx8OWUGOIGPIRco4aY322iPdq0WtHzdHBv3mo
Xi3J6uPivGbGwf9No/5/yDZEDrPyddIJ5dbmNw+gw09nWXDROfV90yEG4HGEiwjhSVlRNz7jCAOx
sA5EDyRB5RiCvn/QESmvmFSz1bOGnhel1QtzCMOspzLSqzM0taC4ur9WpDozxldJPn7Alb4QEVpK
qjNmee3z50o+bbknTInKXcsTLN1tdrAUnEOoxKSQeshZ5AEIWOBedDYaihX1TOh/q4uQCS4YYKz/
tSW5I12ZUW+eoxVoWttjjYZf6IWWvbfLyECxeSkvftQKKkrzzhFOFuhXezZKdcs4PyXDu5CnGD/H
9eYEJfbd9HgwGyBhcoHM0F1/QOVbFj1iQfCgw3DQKv8JHhRVQ+kPkx2nCv1t5+d2dgTX1yBvrLgF
MjUyi+yJXgLh9P0OCw4qZ8tYXR7Oo2QDQFDVx2VZu9w+4DJ2IHrCeu5qzCcqLI1FW1gYLA4FiDsz
FnUCLNIome7qLFkM17b0kMx+gnk4+ekbrLShS+hNqtGyjYIhsc0nhaW3cznaI7VTyIojnBQmRHqW
7dVd56lFWjWG5lMTXpxCsEqfWejDgXyUnPFajQIo2mmm+IRCQ4Qfr57/hQHt2LmCGvo9Gah9oZFz
kY+O48K7SJfdnD59eiaSNoSdMfc5TYLkNwIiFvzwp1puB8AOsJ59lrXBceMwF/G/SAmJH6enjMEc
RyCLZXsLRLeRL3eTox/3h9GTio/bUKEvlHnXAKs1G2lLfPo8fJHipgIJPEc39DLiX+8gYDEImvIc
Xtku+d7O7OXdi4/5k0HG8Cvlwh20cKsv5Ikf+FAX2mT57GKRhDODFj1MGEOJt0/Ti908f03oiMSJ
+8IQW1wl6jkHLXoNqnygFu6T//96Vx7JLR6LoAnjJzzacnPs2w6q0j0ZAF26jQg4M8BZ7vZKiWeR
u682wiljKeV1HU0Vad0cbEzXSrC9Ht0Uw3hvn6hDzrpFDlzd9XQ7KOV0Y+UwLzF4qBtmodOugJP+
0F9GhoUgTm8WSG4bLD4a2WRPyGuA+dNRtih6WN7ghH15mdFj/Ic8xXmmpKa8B0zGRU+bb79hVOaF
9Nay6FIFwBzq+zzokqughqyO5j0dPJzJ2KY3viUXEjm6QTM29fCkFx+w60QsqqpouXegEEd6VnB7
xM+QtS0F5X9uECz2mFQsNv/7kGXdYJ32hrHQSUhkZHuZv79KjrBdgMYJOFNNh9U2/ENK8VlPNoib
cRNb0IfbXp7cJm5xb6w6abE9bZSqXWJpj3P4kUdp9+1Ekl4ed9W4ygrcrnEykBWySBNwCmmhnt7y
3N3Z3NWDAUu1DGkXvPIOU8h1NnRJ/zjKJntqw5J1SMLOqWfeb7Dx8MXBAovLNn14SZF++/ZMrf1M
9m2myppYinIUEMGxGgC/aQMfSqzITHVtO4NhiYQOWbbeMbav4wM93yFe+qdWseWoYkJHTNHxbwBe
kQY4JNSf2T+7tSOKTpDGk5+Jv0idlk4HwRx9HGG/zaoWam5Hq7WqVppAvZds8U5ESUWwuO/tPxA9
YqFYTBp9KcByUcf/3HnVRzYaT25iXmllJd8EzPxj/iqhEXwbXQhwRKOFMGbVpa/qE9bvmXWr7tjN
GLQtONiQwZgaBIaWYINi8jMo6MeenlyUyaIUm6A6GiLui4qTImPMBwwKIZ9Dy3I7ewpRp4S2P/Kl
OJhVqJHc30H+JOJvcxKAFah7cS5VRIMNGvSjsm5AUYr5mCnoBsHAyuOQSFtK2/uJ5kBX/8QDLWiy
zD63Aqqt+p30ueMcNOmnCJuhnxq6iOoxYnBZ8/RXli5FU9yDauqHAiE8cAh+Q9oYywc4ryQtQ2Ia
lp+fkBAutS5egMLkG6YNV1lK+78HETwb5YqxBHJshpr+JfkIXT5vgQzq9zdro4vXOCTJgUoQg4FZ
1WzNj+I2ZLHufRbOwMaEmtFHXr9nucg4pKpnLHLP1wmXW2Cm5OM2+0NXnYfGUzY5M5KOTuhVb2g1
b7WHB46BS/2g5YROooy28AbFE4eGa7Lrgkm4m1NSs2v0nimeYebgdnmwJidToHi+nDMpjVsEeOzq
IgQbYqnyDcgWvK5x3dbtvk3V5OQ7X0442aYIErHzIreHzmCohMCBWniz6OAcmQ7hoIuI4/RFcAlF
doPRjzIs39Kp4yyKGdXgQ71u22EmdIXOVOWNzHLezkJ0PJu30d6JFlhJ1AqcxKGGPZbFw1HGb352
I2Nom0GEV9t5DTyazg2UzfrJfCZMrMqSEIJ1T8TJV/AM4XC6jkvSP8PAyq4O+nKMSRp8v6EXq9v1
Bq5+KmO92v6XOEX6i8T/y8R/H3ynGS7Vf1zGWRDmtZnyaCb6uERrDovluqLTahJo2MLh46iCHmrm
2JPEHxktazzmvHnqhuDjtys7vHEejhu9Brfdbx8lEw//pIzA4bOeYLSWN87wCthxtk90P/+lalzD
Ug/uLgvl9IR9edcio6WB7rEyZoMW9aOV0aNbiGOeyuk32q5tEZBKLZCkUsCWJ9cG34RDhF0Y8ICS
sFtWcUL6mzoID8WapUv0wNmcjayqeZrzZ+jhhegZYwxRgw3Eu1ZryV3Z5qfLsxDlHyMmjQo2kGF3
qJ6H1oMN3kYDiK/AI3+L9C89O6QL4ctmbWhpN54y8Ct0Ps37Sxlz1x6LamRCwzG2KDfNPl65pOES
mpe2K1FlK7UJsLbKEUYeAcqssW3DIvO+8t3GscGQb6kfoFKXhpADFGw1ZQ2JZtNMUGYHiTEOkW19
PgYnaoW8GfWGPtQ++8rRijos3pr+tFBtUNEAtBdeg8XZtX1b83GzDbdb6RQsL3rEycHih5LA8WuA
ptG9ueOcxxYpUGBRWGByeX+2OXMd5BrMWMmZLyn8aUqicnVxsBpxAEwVrk6v3ZM/RPJ1NpVajnDQ
YZ9hzKHB757H414EbovzuSZnaX5rnBfalscmwFzF4CPJHNjNYQ1Bpsho8sXqTKdPINZ1rKHctp6H
nvy2SVUv8umvM2+tTJmjrJaql6ytzGVdCH5KOoQEefl/jtwLY51/onT4uI+IwDgaUcbDcRU6uzY7
eS7osr9IqHQdXwlBgNUqjbdKL2Q6WO/8sjvP573e4D9WEpUrixkqm9P0yLk3CVwudob1IkLCNOlR
sMHFtPPl+Pr6GNGTRrcRQyyXSRZ8V++KrYtNyP7kldTcJclNDTEmywpOFh7bDIq1utwRl19yxmXt
ESrlGQk3Iw4uZ/OtgXlJs30/lUdO2oiIlWjeCax3g36z5KLDpsws755P3ndXgLZAD2cRUmJiW4BE
vpXLptrjcnqyNdF4WwHTjACin5N0RjpPzMluS4xj2raYOc4c04H5a38U3d+a17oHdDb+ImvioDmA
lwdrl/7IDclVqxK5cOIP95qrlEpb5+SKfVK1JiS9tEMRaMF53pSISAwVE3S1GqahX2CDono+rlT9
xLpzus5BGKv4kfmYEJafu2h4Y9sBnERRPR2ScSzu3FDXxmloiN08F4sw3XRBqtI6kSD0TlSiIph2
NqKgxoITjE5Uhg4giEXKfojQpcX/VW4AK0KRtY1t1TYafTzAsd5eSyhH3cCzRttshxq41M8tI5G5
9KvZe9MYGbpFrxEKHsz1FZPLHhgxy9AQmMMJ75AZ251Mc9u9ZuiNum4jOEWrF+wyUARvD/GbqNfx
PslLRa6cgn3KixGXsIi3lRdLQCNqO7F+FhjHjn04kF4543D1JqKmOuxcowXuiCnzQ4zNbFIwWG8z
PWJol3K1RZyp8tYNGDvLLISGrjpmTCNvgf26Iuv3B8OTQLQ1DLyKRmADi2gNsNLnfToFNGfdzBhi
g+AgKuce/V0pC1BiIDKop6opCPXZrJ3cYzD8d5d7Kxurcus4t0qwhE8oUaGIVI7IYMgFAohDFm/0
gQLNTr/ZVqP8OFoDrS83hpv+Twogiehig3ahusPqdxSEGH94QO5XgBLHzyqOXDDkm6my2hKEtP7N
VomSbgKtnqBAUUZlnawBDWz8n/roLejFpSU621KK3apUuqyugMCxxoIOqVesabn0d6Hq1hYGaFR/
p+WIIpY+M/QKCM9uLCd1gSkm2Jx1JCccIwBRyVvUFQjBXveFxggzv/Le8eQ8o4JYMooXBPJT6UMF
vfN7PzULZ6HMLrsTPAU/nrkM0kGoyGAz6s34QQXx+CM/3NR2OXI5fAjRaBKxpsTUXYEjAeiJQNy/
AIgaJdd96+sdcstkzJ/yvScugZQTjhjSDvxIf20bpnkospEwPI/DAdldclrlE19S8I2vbUjwrHi7
qkhPWOla3Wzj3i7QqTeoI/ICisW/bynhJtuNQdjRvHRVyk9eQS+c/rX7dirAz9FLfeHLuVbBV3Bz
smLIpsVt8dT4tBMvPSkLMeKsUZ5VEgdTLcG5C76YUH1t1wwG+7g699dGKN+e/jiFSq36in+obI47
gsqQs7zPG+GcVOCrgAoO1PUWPSa0q+1uxGaW6b1fho5OF96o9NO0ogIgTHSMp2vkGwL8cgZ38x7i
FPFvPPRIf5kGru8g/X034LOD8RPD010pyeE1PXhx+TriH0hHKkhKYCDP6EWjYdSjwrgt9usFdVjl
vqv9nUNlVmcf8sKrfhkQ/Hm+KvXK7bPIJzFdtTh5O1O2PBUSbCDDFfVpKwPhOZ5zkm1h3zZ37Vr8
ltTWRd1MVpnNmhkTemlcuGflMG7hZCe+7ryEksFblCEzgNqaUqK4Fum5MbeVtSpnPVXY2YRv6UJS
5Eh6w1AAMWdbONHpKgjIX3tIsTAFhQWRc9UebklCzf0dXEPgkLTHiLz5g4bSDTOsvVPWyTOziLhz
WYLuIS6C+CfLIfzJ933azY3p5py7YZw/d+KMXLSdBPI7eApOFP1kfzkEnJUtICbTnb/OTtIAOBp2
bSOS+LtcqGBBU4VjK1UMlRthiYTnDy6J2SR/A8DazeCr9cPdlhdSx7W723EQIFoSqpYnr99kt8zw
B6h08KEaXHfAvEqQdSTqi3goTgLqK6cIu/TlTpdoi8L3KTTyOMOCRN6BZs+8K4k7qrtVAAKi38Ge
be8AT/C7iE6JezOdz4a3vrtl0eMyR2ERKyMxQlOolaalj785TKAI1nAnrp1IrTnELRVoT8oHmCAL
s+1GG64jNHc7JDOEZG2sarG9lSv/GdEzjKEURnXubH5GdmoVmNGKJv8sg1l1gQXyHUe2AUtn0SzR
y2yH62DkdGY1j0+a9FTUmJxBzp0vQl6klUFGyXxCs/G9WHG6l92k4AQ4TxaMkj/b/vFouDEM73fT
HjWejwRXu2XzBarTVdVhi+HfalpopYvNMSkIlgx8BgQwAgmqofxMXQ7DcfirrenqNKcGHtyPbU0h
iFnIadcHbE0x97OkytlhehGeSJKxmwPSs6CbTQWQpNtJ6MICNnfwX4abZ0sdXaJdcGQo/P5M+yed
AkxZYd2eSe06ziBaSHq+UM1m5r2b4KY3elW08+VWLKiT+hSYEG0P0YRyP8AdIQu03nRMndWVH5bX
asmsHEZhymRCnYVJM1c2tnXwCkgMHMFz3q6Zpfy+SytoyK8aZ+QAiQPywpozMtAuiA2xL8K6+ypQ
LZEWU5kMTOZMAd915GxOtr4DGqMbASgngMNf8QbbuqyuQLbzFeTH23tmW4zeqzbec06ibI88mCUy
o1cszVwGLkLtfB++bhDP9OO6hFMfS/+qQiBXOa4dvdop7BjMRKVnz1JTPvxnBrZjw/lOp3jIOsdh
kVEym3iHLVXaIEfONblUW4GciLVzj+C5ycJs3u0DgQesFJajBI/s/+aqu49igkSXPxsBQUEDt8R/
uktKsLJzz76oHC+5ADNWvvflBLpm/4vcTe6Hc+NBAS5AZgAHzabmsHPiqRoY9zj77rEVwenIVCih
Dg6UXibPuysjT7yiC6OI0oqbzezAbRWk1WuFt0ONKxQc2Qc/YNBE6n+LOIoCtQ2k5Ab9yIyKjzRn
D7OfJ/VeXb9KxGq2r6x7rwEDAWXcrZizCDCh4s90O3tFmv8ihPwO0Nmw5qdyizUd9sErDEZQhxmm
mrwba3wLgO+iZKgrQEvUltCYqLYzo/dF1p6UM/qxTGcT9iQhb+Z8cM2eJxBUWuxHVL8qBtIRroT3
EWpCnh1+Jksq3YL8AK3jKsj3xEX59riWxHN+PZTFVNMtblb6jXayYF0TH0OT2KpDpk7/uh/aMUuv
rCdrUwJTmW8WE/BlBUADFxQvAGhzDno3eMmz+aZHYnsaLpStLKXAbVvw8TN1PUrQUAVbc7D/7FAV
GRTPCa7lnrSeln5Lut7uGEeSxzuOCPghOSG7ZxgbvYQJJUmdcqUoTNthlSbApEgtbVRrytIikh4v
JuQd83DJdXlyq9f2eya4BrEbIZQK8/mr3PjKPBHhMZY9hkR2c+fsGUKvHRP968znpOwdpVakDLyJ
mMrqvJLAfXQaYGMzX99CCdcAtOaa9uGpJxr8Ak1lKkjYC/bRpGjenySgV5gWxRm2jGL4E9dTxO5x
8Z7YKILTiAIOvZPJ7nKWKA/3ATrH913KVOu/ZiKzAB1buBoWnxjo9HbMbIfg45ctPTGUaSi6FCmX
lUFJbsnp/y5H4DXmNMQpiXKK7A2+Z12orIWkf6//ESTh9F0DADMgjAu3+9Z3ZImxF7antK2Br7wm
9B8/7GKM8f4YDt76hYJPyX8bRBPz0Aq3yzHhfFFjhrxubAS2Vsv0eHI9RUDM662XUKpRhhNlnoTA
iqEJlIX/r/hYhYQaxXdM3zfejdYYlpAJZ2xSN6WzyjRLd6vVu9RMgvy6DYr6Ncx2rU6wv6FFzGH+
dGqQRS3Bbg3wvDR4vRS9ib3/MS/D/GGQyKL5BbLFUsjX0xDEy7RRxYjlO1J3ptWHE/T2qM5+eQIa
fKzZYkeggLGbfHNmG4qint4CN+dEgT1RbWwHwV0p4nuCiGG/XOJ68prLjHMCzG+48800JBzj7+0t
Y9yg/77CT1EV4ySUUkLoWivT5TLaFPfNmFFVyYmQZ4DYlMA5vamh6y9rdkYsNowwRvWWfPOdJbJk
FqJkdk5VDOZTLSpvUNI+MfqPZLvxp3L17yxMhqtnEUtzuPskkHZh/7YG1+IbhGA7UQ4jfDcFWo54
EFu1CIOoYfn3ZcbE+bbLIw8UU3iR/vopvGaDB6fCGm7RnwOVdqojQyo/gJqsKfteCSTUuXChNkWb
JVtnDS7LhBEM0PMFnqeW5duaec3Uchztgjb49W9C1WpGGZiNkTad9d70pux8SniJdEoBsEmZe+hL
GsWHVOONHShAEj8XjqzPFt8RPNcXqvcxa39lW5rSTtKtzccwddsuket98aokudUBfUeNomnJFEGZ
q6MpXL5Icm46fNVJnts81OxIIS1KDNevcbes/hiOy49BQhvyy0IllWED+tDaGi4l89QT8/vwMyC2
fBWrCzIR3eMLufdIhdO8ystS1d7L+TiZ1fryyTFy4tWZgApQky1MkGQbQBOE5aFrFiehhLod2gBl
4C5GEa4V8ZnsrX/BXwk4Pdma1SDlP9I0/lF1GhdCPUiuG9htw4fHFZnOjqMB5kuxxfJZtKktDD/2
qaoNvNYTpItUXglnRHF2euhjazmm+XHtlO28qoXuap3rs2EIY7P+vBIN8CxuJLSoUF/8TEt1BZyG
aQkOQu9x0QU+0yQIIhlUlOejCTRYzsVNDU4yb2JbhIrZDNlN0J+X9+GhccRFOw0dBdFDypUAnCJI
5a1MsKtF7Y5O+QdhpnrxZWt6c1x9mBh8gsC2AITgNlk10axV1kv2sppvfY/jMLf9g+3qakXkjHId
C0d06sUoQ42y8ybaqECaYr/tLp2nFUx7xEdJLJhfolSw7/sYdXvHXguUsxCkM8xkrNSTjDZkYiS8
4NaamWNqz9mbpjpMQBg0hr/LerH7KctOc+VZ2UUBuDN8AM7qLll5NM9cTV5zoEIjZZzFymobEf2w
r9/5rzoZZarvFIFnNjGosS32k/ROO08ZkzepnqjZh1m0koFU21YO3BaopM8+TJh8mzoGOs0urLkP
EPtApqVuSsAQTYM4oCwjVOWQ9iinFLCwiA5i76sv/M3duNRi1ZqD9DNhrnItdiTYLqFilDQ2fFKB
nOHPE6fknU1nCOUlXizhVj+tLyTv2qS+QB0Iti56rDiGPA3IuuGdv4whxZQvLwUugw/Vr40YZkFO
aWzRyAqQBi5wpV0tXC3i1+WvEGm6UJ0MsIKINDUkxXPlPY3voHjlnDtxqtCbAKLkB3sirK+m0WJG
2Tx/fpMY+Th4RhaQq3VaP1lVyNbcPkLw95UHrk4xgzltSap6STB466JL2ffGuvKIA5gp/1EBtjyG
N5VA78J/G9Eemb899bWGDDwdKvLkyXgmIMEKmuDKLGfYsBm/f+MYlrHgSWIAP62bv9qO4IbcEkCo
hxA1rPnNkk5PYHW1tnNGQwWpZUu4pz1bIOHb1JiSdGvRoMYREfHi+f9u5cwI2aWyFUbXvQmRIgmT
60qiNCSoChY6Zgc9C7+WQ2v0i4DcIY90bDAYnIhL5UOGLfNqPiO1Haghm/JmvqvpeQHvRYTZe2vk
HPqLKPc2wC0QpN7zVWbVOAe3K9dIZ5+VyPNzypJd5arEdNvwIfAM4Oj+9gEMApYlErJwuVdWxT21
eJkE1lJw6QJZyge20E+VGXs2EZb69NUc+Yi3yoRSHloMaUFHlRaBzbcItC7ZjlCPn0a5AHYK4Bs1
MrR/gsxmQzJ13MjaY/gLEkhvXJPAz8ZdsEBNDIt9Q07iqKcn5cF6ykCOsWWD4lRC+tNsPnzgcVJg
RjNsZDzgyA/AHHse6nEA39AKmNyr8hZnV8rVW727HZG/UdPtvnqVBgIRmdsBwAkxvCnZVB+w+rYw
u7SEcIwu0qor1Ei5K7XpKnxR7hJYzXFEQ+28DyKYTMG8AuGPVHODChsrigPOT14ZLGNC1b/Timrw
f2/+ereXRWJx/s3mMkc1+TQK402ZyloxyHcb1p2QFhWuFF0zQcHCo66vZERyw6+Psy8jdJGi+FGe
ovP1mjD4POLEay1+F+bDCT2/GZLqsY4UiUr1+SQGvERvTgZxoSppEMBv8QYKqqbOfhQPnkjD2ZY1
KG6O1EKRT/S2N5K515efojnK14mJLsgrPJSvIQDDHzmxZxRcu/Bz6zQiIwlWYdpnpM7E6c799UuH
4ljDkce0SNO5Z1VZsMdkTQjyxTd4wUGg6Nve9bgnFPo6p8wiS3bGTQ8mw3aUpm4+cSegkmA1SYm+
+Cumh19nFvQp6DP8U08hhEIgbkoyi3TKVfiQ02FqWwNLMKp2LkAIKgZ0ddIFN/gAG295E0xHDVcB
Lg7yOmAV7tiMg3ZjfmsfmZqctwIABTh78RkLsYVakRAEzuZzZSkNixQ3V3Qfsu7i/TNbHnN3JUrF
/Gb8g3nJDXmMDcHpVe8jnxHTBvVtNJHQO/JV7G/LzwMeBD0XhrXhVO+lvD/2qB2IERIuR7pdCQD+
7WDUE/DS1N0Zgl7WFdOiJDM5N+l0ZZnlwrJtVgvtnJ/p8WOVDI5h7PVimdVnEYpdPLsrJM/WgEyT
35eVz5vb02uEJECttzPRdarz7nv8+41pog0Jlsd/hEEurhGwDdee7B9VsCEQ3480OqBh5tz3/+DN
v6fctqZkgM8zV+8t3I0DCkEPIWNfAVQycSKlPGKcZvY5puJESZPvovQVsHBxuJcX9/1Vz3MPCjEp
79X0/OjM7ZPfBsUpVZENAs1I9q2sGEuonJ86IbPUgZp1ynQZ8DvG9i/s80aHSlQeNAVeeJ9GnIw5
4fNFkrGkHgB+QUzH+uLkI/w5shAm6Rrc8+1RjUCqol/McWkb6BEWbOJ1Zl+M8G3/QlcnLhDAzQjD
+IUtc3cJ+WgT9MllFrWpUjukg6YIPwelg9SM15BVlXK2V2RQBYG7Foekt49PWWd5bNITzhQre680
LdIwwiW3lMUv78V9WiqSTQEXRZ0Vb+YL7M+WVS0aAwlYazJekcP6EBIu9m6W2jY8ayNzdYGqj68D
5NZMK5KD4lBcDQac3K/uNDXiTePGl1fv/Q7sAt66SI1aCTAyQChqtdjaL/u+vV2bvlryiuO5P7gW
sryHkYKmlGjIT9L74YM3CD3clp24zzFK53+vkTuKXgSA5daeozWajMW5LCugxFJyyz/EJenHrU/N
oPpk1o9hMc5GRAvtBbegYyfguwTU7TNPAwXAotSQG+DOGTbMtp3YE7xaLoHgIXOzfKjWovdTKdrp
AGxoDIco/TyXxTkRTLjN8fYg9RvFdKGyJjEEAyUuCvQ7pyhKNstVOh1IdDIYdpzM1tWd9iJaeGlk
2sn1qjxoSsV5tXa4f+OJCXz6spzYLDbbSjpI0Y0Yqw1bB/QXGVaqoqMGSheRiN8EjY+YD3FXzINR
vNgGfteGbdinMOVbYA2/c8yPITrYSkJIC22pTButNZAd27QfSRTr0Ep/b3yGOqJLALxVevdxNhOH
MgPmZpOuDYHmegXw0Fn3yB31t8WsiSMC7ACK+/iQ+StVPCs6qJwo3SQNTbKX8tHBBSSCmxcZVSQL
heIFErur4rbu3GxJgVuKzYmaQESUi1eqM08nhx517rZagOysbAlCUL2vhIJXKO4wlw5W/0tPuItl
lPigi2WqN4xfBscUnzJBAF7kFq9Qy6G0lnbvQ/pEWThrC27acMbB41zzcWvOYkBKTUdNLoeLzJ+Q
FSnAsO8KIMwjXu7h96YT7qjnbYTsLWQuzb65uwj4In6+6sjgIOq7vEY+9Z4VNJgkBAxVDzEHGDgP
SxpA6/AHJqiQSFgFBwA4WrUN/Sn7pRvebKijhW6jZ9uyX2XFSf8fQqIG3+/4tEuwvAFrYFSrPwtK
Fu6n1P4FnM58lk//ZpE0/U6ZH5damGmGC3FIxREvJbjSTo+1uceT8u0y8uxThdpGng0pLgG4oR8f
7G6S7HYRtXFLs1W6CJ7f64etCOPTcCOS1zY0JPQi2Z+CuHyX+ROA6n5aUaZW8TZoai7eOxKS/xJQ
jFIR3bKU2kr7xHD08vvpCkOq7ZkIMeGU9WN8OEiNxrWqdUuTqOfzEb0RWVVcCoBaJ8f4OtmgsatX
84ymX6srt28dIGSNP1ugFSZaKffiJl5v32+ZcM9OI2w0kGaN5gtevzL6++Om1XQ60aB6h9spAFjC
cwq8QzMo0yyuP91Mfxg8rDVBawacYRfA+QLWoU/4RR/GDztnLAmQsCZjgK5a58rZRB2BrWLq5/y6
3vbsRU/v8HKpj6CRqq+Zg0Se+bz0TaaL8bG71YXktt7cpATiEmwLAu6xWEBGJElsRBG2s4mNSPpW
TEcXpGwGQQlD4QKFdE8ZhmewxCLfFSo7eaIGUSkTLEfco0HY7KdMZXm/Me5T2BLrViThuZLUwHyK
AN2/jvYXYt8+JN0f0vT1G0MboF9EgaVtGmjS2AtsRFzCSLVXaOaWWh8DDb7U2uKBswxX0AR6fukm
bWmIbj4nb3els6l1acdY6krNLdXMmGUMdd4j5krDwsnNRUmFsCxfddFJWJ6NBUngJfrszBif8o4H
C+MEZCktghkobast7vg3i+DQ+ZcbRoHAdBIEX8iEMa8Ai3ujfniD73HayNXG4tH17hABMYIH4spi
ORlu+gxqZX9i9FDm13I2Q1Uzzvg5T5Olsax6Brp4xnQwRBjC4FnARjB8IxaiRC5wEoFz3VqHVJey
vcMVCHPDF96E10cBr1r4n7bqHpeVcyh0BvbWFvFpWGTMScm8/lTnarUZm2+xnDFeBfDvuNszTVCR
CcTJOSx2/EMQbXDxAeGmuQMGvVbCkKZUgUclBizqv6MeVVdGbcETbT4+yTm6aHRpYhfqY4Egi1CT
wFGTlrbqBEDSuTxNVD52JcH67xycYbxajMeC0gbUcB75Juyb0JmUwyEePcVNNRQt/1i7ce4LGgur
EAdgZbp7Sg20dXJHeNFbLhroXuTSzRvMnn74OixOsuW4u4nFBNClvr5A/F4LMGADtRYcdMp+jzIq
6BRRqCi9vhyRRmPIk8bhideHwFR09CAhsphbmkWtZ4RTIcHGbmB2ai+UCFBtZDQQdbgd2uz07nJe
FcuFLUDihauIqQUh/2kO4q1c0ly+R3ymdw9CR+StxREPfBX75+R4NsQVcIBTguqV1fauuivaxLln
X6vkff5cMjrTHJ9znJe0YzvqYuqPNZ2nvhVRycJPfNyItOlbj/bVsEKgComZ1+WbCYCelJpjROsD
leORjvSAq34gYhg+PhPzCQGr/gU7hX0GoTFuLmS945AQ+WA0IxEgNDTJo208UOvLGrAMYQKKQQu+
88o/1MwYEDrpfpRdkbRiLOiW5vBuB2YxWVYF9zpsTfEuPEGsx8TwqkLWXWnlCAQ+BRhxmjDMCoWI
69nWQAC/8EmpAkwQxNlnBMPE9qgw8on+5EBzXFUyOClNHmhCbRaiZyqOb4q9M0D8EJxll7MlTL7Q
VXbe6J/JLMsW+KjOcSjc4vbcxaVKwRpAiZZ0An/knRv+XuWgjUevb48bggWy6Uzp9Qw0uOjVjv9Z
DJ+8fqw3Uhl2WdtgAD74GCWqGoN1QWBrDUv390cwhcQc0iyEwFZwt4U6YDzkVJodwfXPtB2frhvF
ERJqUtGLIehNzl4isII2w1s5gjP0WmAjy6SwHcHPxWZd0Sqy47hQx1FC04EUeFVlO8zg+SnkqWW1
fblmF+fG0kLtFKfZcNPXgOZwxKXn2ZIOxV9ZKZb34onK4iSg9hpOBGxQZV2wZ6W6CZojx9DaQs7V
ONOU0AhxNErAVqrKmS6HBjAFIEl2HDR2wjuX7LsrEikcBsMhiX4rsx6iOi9O5wEbPT25hAjcOZti
cAbePaFuhKTLXeolVm5OES0Dhmvo7zJaEis4xdCvo3eZ4ozat4SbE3B2d0gNZ7gUaHb78atEqFVX
diDRRY1RL55dNpgg3rq1EMOHfR618iaYZ5KKvQEu8Eh+D4bhGd10JWgiIN3T0+2rJkG6wW5DAMl9
+dV623vwFfwtCHk2aFn0Tg1SGNTQULiNaEweP2+PCwYXFD9BjWjRd4lgKBZrjsODWQwXHGZxZ9cO
7cH6kYCHp0YAwbvPqP9k0w1PzFSWLqOZi0Mw64ttYBzWVtkpLDAoD6TTlPoPkx1gwSgRdxWSsTfK
hBKKRpvS5B1vPTT8Av4JzDIefaCUzUnh72LgzYZbuqb0tcNt86RtH0Pd4QScVgvNrK3pCYf/fLIq
bVXEpftmn3qgdVuRB4idhfrvgEidCzVSPfvS90j+VXnewfJ12fDVcts2VzF0clVX5cyTAfqW2b3r
fPBsOywP/6tNPuA/fnXj6jWD4Yr9AVhFStUL1at5mJ3Psq60FTQwpDKQUOFUqPnG/gyLF1eL6PTi
PcwCvhk52i6FgAIwhlbA2frBA4Gjfo3UiUvqJReZLkTaa4RbGfT25AbYD45vJ+fkqyzOiRRap3DK
qvTGBArPh3Jv9phNO8Y+oAx3MCJsDQZRgRbnfG3N5mnCHbtdbn375SISu+mAYtx790lueIH/aNvf
OylbOuTBN7sf7eHv5h/6euA2iwqp6yKKK8NBzSY91rKsxYbq+jfdNhgQVJyXDYquIXPAiVoDLLer
7y0XtaZtZnqefzirUNOjcD4jTdNVcHulvb5LNL7aTDwMbApqqGWIJ4XJbqK0pPp3nfP/BlNGemIX
b4XP0rUR17uRhD3kyAhEHuD6CWGz2QrkucKaaG+B69h4Guwe2lEsIEcuV673CevvNubjYT5TfC5L
LbiGhodA/N3b2jiyysVwf0i4l4ZTd+iIs4h8ceR6jR2RYQTO0fVGEZj6awiM8U6tuGC7HxyrOrDD
rEJqqKAw367jG4TN76cmfdKKkIb3H4h9gYKbwNkKGACDUei6SqyNx7bOXag2gVptoOx76qiZViM6
hKMP3IIuZcr1q/i33SLn3KwFpeE7wSWigE2Oenl8t9yGecm3xycYplDOlhdJWOBYN+ByZ+0bq6AG
rdhnkhRUcRNeov08K7qwg9tipDvROhAE3fsx1LeiSrQHhi7Mrv6wpFBXKHvbUBBuM9YumSgmvEX8
06tJRKdRWFIhJXOTY5Xm1aid53SkqrCQ7yxvwTNhLyH1wU0u89ZlRxL69IanxbNNI5ZoHVhSlHIO
n6n1sjUgRf1rfcKhy2evfJKCRVleRylf40AwAH+fpWN4bnBlBS5SdXHdMi1UDuiHeFHziLsZM7Y3
9OzEp/Y4Q8/QrADM/4ZHcnP3Dt+OdTL2FFAcAI5f+61Iy+3N4CHAc5YR4lt3z/pfg/e8UISqB1qC
Z0CeHW/jt5S/3b9N2YG4yCs5tbiQDQUZlMUBrxn7lz1B6ivGhbDx/HlZeBAxePyZdJxbVFQ80eVe
uYnf3mkQksJT2pOxj6OFk9cEfw8+/dU8uVj2qWTr3/NslqwIzvo9ccL4q4aV8pEF+1+Bx5TyVhZR
gEL6JsXvKhDOJ0Xm5FdYkSjB049poV46/lycuXAfD3Kz4UE2jt6JcDfUHL55teqb6xnwxVux3035
N+RN6vhd2on6OEPtvicZi0khQVDJ9pe81VfNsLsboYd6eiSkKzPVeHXgh+OPqUVahKa0Yrt8C97I
nQI+PLr9R8fPyoTKbczeJ8ZPjOwm7GRgPHUVV6p7cvqGUctWIvsCmh3UALQPJuoTxPxKSMG4NBWi
bglcksHvT93+gDj3tULr0lCmJYP9TyXgbsL275DFqQ/2VLH1/cNlUQFXnQVKhns2UGKsBiiTJrk4
yoRs5kuU05hCh8HpVQiJ/UiOQUhoHdNF3Wvt7BZBC9woUlZ6M0jiApN+J1gLA+nYRSjYQFe2lEhs
57MdNBQH1M72uiOd45t1xDn7SHDCqsfXB5dSixt1t0W5uS5rM/Mc9WYcqevt6Hvc72TGFIOAh3l3
mz2OjICIQEfqgU8RbjQUKptv6LHDWuwYpXHAA1hMjEaJixcwB0kX6VGpFhVuNqKKGib8qmAhYrdQ
G6lfXpda33WnaL0cDlugf1bMjvqwnhO0LUmcfSdnKnSqPdFbJFxaiOmGvTkCvidt+k3jM1PBc0IF
jkwjRYfVv0P+Uxm65pSahBYWX0EMEnISJcFml9shePeokfDSYXdqiv/HsVROKEfTzZfIdkWUV/uz
I8RB4e4Nsg+FUW1WyNncele0FlmUx2oamYXnLT9UZ43NeRpFaH5d0lzO2//DfcBPyn0G/7zwnplm
fQjfWRM2ERfhueifWSeit3rGbI5A/ZpA1wZusc7+LEtBut49nln6Xzo9Kx75lfV4b43EqcU+QGag
lSjulaISAlrr4doTpGkujbPc3mdC6Glj6g4mO4mpGHPq601BrSrnIQnQBtU5PIzDK5ZP2ORvajp3
B2XGOSBgFQNkx1WB/biU4VeJjJ/SXdwmFvXBTk07i79TO05YAUTAelV9fIF1Lj8GyuNuEeAtBF75
iiWgRwO3djnfVg5hVj338qyP3O0PNb1j+fd2k8rMIZL4aVF+YCOXJx9rFIPT0dO9S9P+Y/Wcs1uG
NWn7T/zw7n8u5QgJHzIbAIClxiCxFDlCzBuVX28mzGdmWUj+inIy4EHfN2RTF2QYR/RwidbBSaPU
nKAERQwN6YYD3iaSezYrnHJSBoc8xh/+qaigN9Ty2mc2xaA5WuBqO22jECB1AX/PUNG9BmucjDfr
eix6kJ/M5KFOMrytUveNSQNyC//tD3YtA3UHk3PFjsACEuZvyllOcRTxsoubXqRNIq0XCBVxVarK
2hCzfvTiJ9ip66Ph4sKVRDbXxDKZd5Bd/s25ls1bu/mclTxp3mA8dT+m3CS1YAUd1Ny6DKSU/obm
NItqV6h9CgoTgNdNpbtFZA3AB2TPMTkN48QLoh7kFXHb/LDP7rAEw5qoYwzNKg1RPKfgthXFXM53
FncuKRWDQPI4vAloKpiemHsXQA0kzQWYCmxvAryKcWUmQPYaCtE+zV/E9ylvQY9Z6puKvCupurjs
+aQnr5W+H+sxlUZa2L6IarXz/d7ZJKcgbF4SnJcK9vbPdujgYXgNdoHhKh71ZSfmRrqmQWCnAYX5
tYGT86aLcWCsaFoa3swU6YaLYeAKIA3cd+59c9AHWsMufuR7D2aF0qcvP+D3qTW1f+XW/YR7LB86
Pd3HCwelXvgxzfb4umuDxtqckf9oxqVh0XnLOxmCwrVXiySa8TZGDz2kJ0Ta39w8+wzoeHgBf5pH
dUGFq+sBZR48GrZ+gjGVnwgKLKwwl0LVzoB3oWzOWh4mBmuGACz/ahsozuuw02XOLzc44MpvuGQ1
+fpfGaThrYCoRmMR68RFHVQw+rI5/WaZitkRsJhdQLOpLnaSCzKhSVjE0pmj//N81aEz0FrBir7E
GXBhrnSaa2LdV25dE0HUscffK+6fZQlozPllRNL5MgUCs3LEL0K+720GsXiFdH0TufWs5MWAHnpy
rNtVsPO6IRlnUQaoZJPYqL1hGgcJgxXejNq2LrVgUmKCMqNI4vC4LNIh/6KqoWVXSb78BMZOyzNe
GmGpdyKvzWKn11f3xSgUJJtJInceoACBDWldhR0+T/sCnvMTVYSGUFVCLqO2BPMJ4nOCuKrokdDN
82wx5CHSAMrE7PUAQEqc5ARn420sSrdh/Sd2ZsTQT2R6UCD6ehwzRLTT8fZACKEpQmQMtXkweDfM
OOh5Ewh7RbJynlbkMB+SwYQbTrDHXD/5+WBhhCYsKrbspXM07nN975R8LEH7u6LKF2PbZnpa5jsL
D/B9bbipD8EUz3MPabo6jb/w1aslphd0ZBsSrLyCPZJq/KxafJ+/ZUeVL6M5Xv8skTQtR8XNIhka
lEBJH8WbXCviXAMVt0xFos05eq3WhEl2QMgwNA1EileqVcbIR4EHa6I6zRYjghqP8BPwNAWMQwZC
/Ry9ONmcrrxbq5XZGAgFi97CLUGR7MtQqbj/6wPwWo+WF+cgWMCEo+EZMbvmrRGjHQxrzfDzoTyh
Uap4hhorQ+ZyrWECthg285GeF8sfbuOoShkpRuazD+HS709Pgf9tZSOL3l7L2mRinfVq1DlR2qoA
Q0+IKnThuzjT0YIMrw6BH9xGbhnZbdWGh5Cr1BkLBdwAkYO2sVdxWpGnFlq15EXNkK6tW622nATX
Oe8bbzt5Q/qWzCD+IyVERtv0YW2ByV3vFeJXya624rly8Y7T0wHot/XVCypNUQyRMFK2WgeQ77wA
NK2Jl5UvwKVQ8hmCHQmrUovWQb3S/QmAKVpHMMD7/MGflcX16LzsfMxs9lkNwnb9LNqKuwObd3Il
ecsrRtuZJrZ2GnxXsm0vT2w0ffwWNZ7afcs/1/ua74Hbbof1HpBxqEc+ie0rEc0OmvJJZqCVb9qz
iqei66cUatvbMfCzGftO8X/uXfiQFCtcPEpuiA4vqBylSWrn6uTGBuN4fRDez5GpR4RAQ5XBeC2r
i3eFs0dxcwVMgoAU0hf+jyV24D+vcL64II2AyojInGaKLIKrMAwPgGKAHeEpr05Laz8Ds16fvDg2
rk5QGJTzVc7XYpmJtxRC4anFl5wnVfyXNnEJxbJzIOo7SimTm4nE4OeM4HOIDRqZLoBt5LedEaS+
he//Pi3+2iI65T8/VBnNZZ2OnKv615HfEMBDvLoKqz9qhUm7FD4pEYrEt5Tw+MGRdSwcTYG1oa++
tQII62Yk383Zb/c1D20UzZqfAe8qD5k/DYxCWhESKcLPG/v34MOzVg7XMfTwb46n+jemNSGVCeDC
XnNL6+oVZMHhyQuw7ZXB6zqI/Xs8DmQ53P0Bb+nIk6FQWBqRAlZQaR3usSk/G1es/h8wufCsCfMT
N4iRQOg7HFxg3jIXE0Xu1LR33jrya8dsSqHaNNUBf5Kxe38o24XdVOxt+C5CIdJfe0QqvbRWcsjr
ccAtR6cRgLR0zfJdYdQ70NZZSaNb8IVg+TsBeqM+PVa4yeEyajNHgWJEax7AGgKc65ljvGx0kzFz
w3tm2YTvEDs6UEZ82XxFbV9MzJDETVMSZ8H9vz8R4rnFMVV3VtUTOeELpIhIo8hccHkR/Njmd7ti
WgOArMj4x222qalYiPbqVENi2x0SZtWWEs2Bh4jFjPnuAQh0nUBmJj7u376QosMeANIsW/BNyCvW
GqK7M0zr0Pto3SRRPmNegVoP7UVnjIYUWB7GgqlOyoL/S3PSOBxWTAASQ5VvJEofmUVq7b6+e2Cl
SP2AO0noff1Pgd42gqRrdXEKNoHyVXl8XZ45XEz/FCaB2ajfV1Id09S/Z006tlHjDlvp8s0Rf5rx
PP6PZJjJ/oyyTgbAMAqMDt1Eu6RFGupBjjb2yo2ulXykaaufzOuVJSlOkcWmeEB7Il+6guI7oitO
rmpLKPD4/etHzNt8HrIiOaMP0GSPTw+Mi2Xm/t6PM84pBuBPjFmsIEtYv8HfJPepKvnecwnaYgri
CMH4CkKGcB5EFpIwfSwP7anfD2xNgejC44HCly76MJKD6bSeBM31qFPz1O+oE6ABzra1OKuYx06h
am16sUyMnCb8onBafzwZqVWeI18UVZjA6fnNYA+YwljMiKr25VphX05ORsDtoYB2EsTdXE2FfzGF
AEh7qqofQZA0+dUKS4dTIN55GYNobhVfoRf5RKFlUbUz4kTSVlAh6WweOrBbanLm292npSbPc2ne
Wal35WjJVwVxZ5oONxHGq4oHs8D3QsCUb124d2IOHBDUz0F7k0oBlfboo+hQF7Fis9qkL4k+aEf4
oAuxX8GAy7eraVTojs55pnS89+UhFGd1+6tEOZEabcKnJ8k9VXRsU28tvScqFgtpqJJ7uMGx/LCB
vA4W0jYG97NhOjdPV/2+5IrRjMkJuUH9tWmfNK02ga0pjesHQ/qlrmdmPAwm1lJ3wqyCOzh6tCpW
fxXAIpaqRBZJU4yDFyo3xJxz+stYtm4QayFVsTgr8o802S7LrWvlljf5oF2pJxQ50pyvj+1OsyQI
SRJHFon2/f5nPVFa1scxchpt8zq2zU+CqQRzmIb/ggisZGFOMaf522+CXfV6RhKhaifYVXLhet31
Kw/4N5TxQWdj+lf/Es0v3royLVlEcczVhDz+4jYwIKR4LgBr66m+sTOELlCpZdYKUMfoSc2L6amB
KD/8uyC0lpmeQ/mP64UFfbm4HDd9cIMllZBHYoCVC5P/7jzdmrYlshGLrbfHOlB6C3a3yFMSyWXf
6QiBVcxmShk55uxmwHS8lSW/as8VeO7/9LejnM6eh7pb3N5dL4Cb0xS8kI5xrxefdhqdXGJXNQ6H
tZbMNOE5ffFq7UIoEtBAVGOkUnIpmQVIvTF5zPadbuu/5q9xzZX1qnk9nOirqh2AmtCT8SE8nX3r
i2AexMJ6twQ5J7kArPM+iWQoCikMk6blu3CPOW8PYGCzsbKgRPERomXOIf1XB+CN3mhE0Tc9np/X
07T/6MBu6Fn0ky0iqE7yJXs3TV67TPG4PB5RK/87eK9jw1tQb5fK2bUkulvQq1xzAhuVQkW+qAa1
P1y5fAZqkiZFo+txOxjl2rNhoH+1BY8VWDLG7YJYlHsGuUnfGDb7sE+N1s87KBNrG4XzQjS19aDm
UoGwJQUJkPnehcHO4Qq9HFEbcQLEg/t0DfhO8tqHBBnwxErCQ33om7vwITQlCFmzAUFwCoyweE+0
5uKZ/OlJlZrxBHLH730exckN2LseOBfxUIcJmYtZirKI9jFxFPEUsW+iq+oLPEYeO94JN3835M0h
j+RVqtsYu8HMYSZm8D/SWHtmG+ZDBYZMYnpEiQyk7nabI58kRuuXHjATSy76yQnUdl5UkYEy6hPx
Sc9qbIoOIHkT3oQKLfqSzlSuMuG1JMgbtjRXxI5I/HgB7kRfDJlnEAqlcSKDkF/pCzGgzk1iDe9L
2CpAaHOdokf9SLKsM6V2H/PilQ+cIXmoL+KX+fmsvAOMHR/W9ytQgzYQwXhbxhL17FS2PzU4BfYO
LWETvDN8Yc8TiCr9D/ip+49oFcydPvdCuhqf+/kbOa20T+s5z4OkjhAzPFV5cEtisXwm7/bMNep4
x77xV7hWRLieE4bQvukOsmULylNVu4rPDcjxWnHa55/sEQpYWenI4DkyqwEk9tMohmY6WAIRvVQ0
SIYzi9fkzLqpoIT4/mBmsoQ7Rmkb4EOuXudNEbT+OVguFzN40Xjn4cxe1G/APeuR+HWFjmYgB2nV
wCgmGV1w+B1B0THQJwUQPX1umIEfa7IQC3Z7Attk96G+TD656jxYU9ZU4iMKtOF3KdDissAWOq/q
raH9H4PwhU1SbXTzc9muuIuqqWuE+e1mdg9VetqXjCeG5kZvMpwJ6qeyAz95hxvtoyRhoqKaBUhq
+hShERJE/wHVrx+eFh74U1X3KqhcvEh1oS5h5lPrlqGvL+SUNeoYLhDBNNv+hAyDpum1FxI4to8l
XbNt2FzCi5KRuYeEvOpC6Kp4gc4BIOVOEj9Bgf9ZAaKycqokXg8dZtMBD9DpYdcEcHJp68niZZ4G
GDzhfxCBb9CeDDfDQgQUGxW0WT8A5wkMTwSe0fjFwXwLJgPFQEwS/R2aH8PNkFr/hYr4/Go/5PCk
Tsi+WkU3k627XMwCCBD3HqhQIMdkSJczVPliTQ5kUbzmJHbr9Ppm45xj/eZL5NpHcSanyqrJ/WQA
BAzNd+90Y0xpcV8QjuXfy1VTJTqaIdHCQWhv1sKyqitPo6eePOQxZ6OMPSjdB8fAJS/+/t9149mu
ZW3sXa064toWHIt/e0yr2A2RSgktzVWadZsj0kIjjh8Wh3jtwSQoyaw5TULvpBeMyc89YS1W3sNf
9eh74oZrAVBWEgrBGlqFe1vMFxKSmAhJx5TCagleIRz4xgUgC/DHJgD3CBxHg5m1fl4hFOmIwdtw
arxKudc9xybP941x8km5mhwyTcme8l84K+YYNzjwZZ+RXNLwHoy+Xr0zQYhj6ABqRC/e9jLaJw5X
r5pC9sN1WRrzfN6pYVeAhLHvuciOddO263psUUG4Ryb/d8eT/xtNb9b51mVlK0Lth918hnyvUZ03
skftE50WPRrmG1nXlMOd8vHZiPETORcEts1EsYMHTB3HWSv/OBPIW0SY4vnXIXG3Qp+ub8jiZ8UQ
tVaf/+8Q1TT4NAcxZLorZbdSqJoXWltSv3JaquXG0jaVvzsq5ODgbrcCWZSByBMcXd+dI+j82dvU
d4c5QFDRJS5e4bmV0vOY74yaV1a7x+c9GKS/Rl85wVve9qTwPoU5iN6bOtwqlYgYKldS1Tf61Y41
mhVe1RSg7u+cJe9gmAXM4MCim/L1aVsG9BnuXKEQG5HU4ubZ48hv+1c130Rj7ADC8811Mlnjb4bZ
YRQ2v1L9y/s1y4o1o3UmGp64dfBNx4M6zl6rUX/wQDYZvKEaAbF80ddViLuFS+GyaHV/Ta9NBBty
dyUbzBA3N9+nrTyuuWa6HvJ+eG2LcTOD5L+LO3+s+ckOk9b/YszpqX4j5ym1mG8VJmI32ux3Xk9t
3hvNtumVT9WY2vt3FkONl8w0/b2AigTBlko0ZlZOF0Y71ERs//97UvOGli6LkIYYi8z4ONYLIY6u
2CouYpYz9gYy2lDfs2m8tU/iNMHvLHL+SJHYaF/rusbFwgvlzQ655+YUm1PPyWpiWlmx1T1wHw6e
891dJ4dwZvOnKd4egSm48BlBBcZjTSaHQCWyTeyds0Qjljj28iVIjPlU/8NMvuB3rDz9eAMs0MeB
+Kot2UrYe9NGCCbA/TATEFuHLeQ47oAaRn2TrHbIMi7CVaSg9OFlH39nFtqlS6vPZt8+Jam7UOxc
Mlw/h+oZ5M3RfL1mEtGsKcbYi9cU+lerrRE0FasBmY/xhI84WKm2o7aCvxtwjZBT1ew9TRK0QHo1
cpftV3f3UXtWfdxVMJUKhd5Voxz/0jeOOq0HGBAPCr2VQ2v6BAMagiAu55VzhpYleVeHpZnskmFc
Nmj7EOnspPWTLJ6KnwdKKBW0MJ0ogClomVKmNByFW9vQKrgK7d/o2eXMSeG7KYiW4gM72p/o6paO
KbOnNmLP7dUio+socxvHzoslUzF2I+lC3pWyDZS6RgFaGmkuSNMGp0oQJoOhjNSr7kpsZrUZga0j
rUTNh5pF3jtEKqe0KooZVWnFU1xyCSdK18mIvQYSODu3qSRpVvNgMQoz6eK/W51oMTPWMPoF7z5A
iikG/kBka2o9FcLjUgkg3LJv4qRsFGKqQ6U+pi7KCzIu4+OUwbIvIg+SbbC9nDEyeXYYPx6HGo3a
/e1La681tHFplyTgYjlDIRDWmW+1Z59hq9rPTIq6+H/7A4bN7cqS4SrTJjk1uyjjylpK6ynOnVgI
QSueV0/cX2zdqC38eTlK0lQ4vU6AaB4M7jkRPNUdB5t57XwyxlwHT5mgzspi86PzQYskchcWkeZj
rPyxX8ytVj46+DmpkRk86zD5SOjkQxwWsxqAzH2mE4wavGKZ+I0BKcioh0HuXkAVJHfKy3wziSzx
q/7EEpLKoF7QRA73BAKSoVO+iITqu85NLVr7MQlbvEBUSGA/9dgkhR0gsuhq7OtvsERGGJ1xCRf7
G6rJBHK1+/c089TFgVRpfvDET6Cpk9aShnIF3ZmoINtFQ7Zb+o5O6djRKLsiVVHo41jDg8Jue4MG
nkpYHYTKuN2qyDZ2HdDNrslcuWHPpC1ZcsN7XPsxt6xw50V5/5zSkliarfcgpLcR3JM9CNdmNRQD
g5+dHZLGwqIM2uewgN70KThHy57HPNDoRUWuLtwVcBLx08HlB1i/IwufCjuj77Xnv5hb07VKkdoO
ueHZVTiWbmiweWoBk8X/aPo9K84MZudeiXOI/JmnXmoIOeNxHy6lSJL4DPqTIt0Ow/mh8TODSWc5
IY3InpEGcj5CTxEXJOsfbkImjcyQsutZ+84mL6QVjv43ml6sw5wSrmio0CbXHIEbKfxS8doiVImn
/lgDB48pZ4FNiyA5bHS/UCAjoh5Jap8aB9KQ8Rm/67v76Vg3dqxqtfegs0zTAgqjeze3td/ureFQ
Vum99D9becBHTLPW2ArkjtX+UBzmLQ2PlhKRbXIS7zEL4gcSqexgWU/tQQd1xN5LXxrHIJ1t7zss
vZXigXdb2J3oi4om6y+MWNaq2bIt/sZrF7Or63BbuAxnJLVihvEBDyHoiL4VxR2Z06Bo0hMXGfow
/USd5el/ay5//BxEEzLOdqo4BPwvL/F0RR+wyrQ3NkND81my0LvVcKUX9AidpYj9icHf358lkAqF
gEN+ot1n5vDCXTPPzKSs21qXwAsfV4F7qgFiOqEErR/Vkyu+IWI0zsRJ+UhurHpdPgnkRP8cCPyL
YrZcAHWUbQ9Umlb9VezIFhRBSrypgunb0CS15ftwcmTsCpMoS9w6SsCMZzDURWZ3g89g6xEIePzG
1iUESdVGw4ieTzIEwZEZJHuqY4SatyRw2xK2TlHR8DyaYI7HA1nfjdlpNZkYz5ODFGUsEriHiEB2
NxQqp/L0AoMdEXyl3AXSUnXp4KiUnostL6O6x5V36D+oum339XjsW0HNNeYh2w9aEyYxY7tstvke
0r8jM2ljEnBXJE/xZ0Mk9iCj3O6zPS7f3jL87U3tgBEM4UFRbD4U8EuQyrxJZfoVLlLEzffzIGaJ
ioeIm6IvcWhjmb3cqZ7MeSJkv5gU/B4hoeGN1tvK9iouIsjctFLaA9xx9KbeYq8p2MSG2N3b2xIB
wsWxhzIL40gotY8AJuP8s4INGVvfr6SRA/jUdnxr3Gf2RbQzk9ueGjdNLf7N5bgi7e3fB+WEZEt0
xZOjTQidTg9d0m12kXVwvuG2J327Mah0PDgV0mYZ67UF2SHCEITm8/3dtOIlL1t9W1g/Sn+XQXhj
eRMWIAMAXouo0VAVSehSKf/G7/0a2AIKXLXX5h69OWylwMI0fdSzO9Lt0+Gg7LCXTkm0h/O9lWic
nCqJIX9+JmRoKyG8oxUKEiCeWoJcKX6tV1vaax2gbYEFqVaxI0Czm3O6gDLfjUDJZZQ5qUo/Os2F
s44Hab9oIiKqriY1D26yxU9PPzzmEdbIQR0rRZw0ljaI3Vsd21CyWra6YefXRvnaGjQgh3UKWIl/
XC24Bx+vR7VxT88/W30i8DMg4ZebQzbYPhJfo/IMlH1+djr5DXxZKpGQHFHP9/2rqzXUnNsvaA1n
WBPJeGeSYJCM2vDHBpYMbwuekjxm/BCX9ixXmkJA7UjtxGoiR1KVpBe+UdbdiVR5QZgvtnIq1Vzs
fWHl27PGgy7292fuIilCa9SOtDaMsE+InLIJwsoQKPcfAWVXGo1LyeT/gYPMAWZQfkFHJvJEgmzS
f/vZSom/8LYv/IrJzFtmf5/OjTaH62wyLv8kI/9oN+hIGG3dnFbTMVWTkuqXtuObqce+/ENy6UjD
NaFeZuCQPsLxCZfYPxxJNvx1UjIBBKAwIm5wMFzRFLWyLYyhl/NcMeOpTFaaHHxTW26GG/J+PC2w
yflX30N+c3LfAhd0GFsi6zORnjtqC5tr5NjeYZPU1qBIQebrCJOkL9ytmlLbpHbC6ZspQeXsmj6n
Kn7K4Jfj1S3rljF6fph0CBrau2ASsamr07Mbr7IRWWGKCkGki7SfLZ4U5hfMK9NgU78tv1d2qgom
xUieMshvF81VMrrBIFsDxWtn/QtV8erCTjkzi1y8Z9A9n4Fq7bJG8zZbOdU/SZRcRVo2bKzO4Goo
PGDXFkWR10t2dqJMCi1I26EVVdb2/PqOQOccCB8JKH70Chf4SoFDsURl1z6ecn243Omjhmzqf1P9
0d9dtlhfIF/euTteRMitEWE4JU66Cw5uxUX+jCIBORBrOlNr5kZp22XiDZwAslEp1PLfqnYZm2eM
6Od6wmOL+xiAs3VV3KCgeqamiBVXUYOjp1vsXlxOr5uG5h8dBKD41Qf2qEPXuit0tdaQIbN8J8Sc
qvRReVKFLQSMt/KdWfYKF3K9kAOn6ks8SQ4NRbSfdcewQnwI6LPMu0rx0m+W/v1zOHsVOMsgaXZ8
+QOeHsC0D+Vuqss2ThbbDr5ZfGR+5bhYIVhoqusD5xk5zrA7JtqEFVdkix9rJfMNg7qzoQibEuQl
V+bZImUo0hZqKXV7KS8x+6TVMQ621CoVU4lgibIp52ohQPYvew+zhosjnQLfgjOTSy1Zt2bZ6SG7
RGlQRizdI9DKB3qVpDuwicB4fhEXAlapkPcilZ2BdS3i8kf8aD/Iz6dVskJpLxK3wO3r3sZIlWNq
DsMot8Muv3XntrwYJwmI79YA8+boUTNSLS2/EbUfqdJfKJ45bO/h4lX1xGGbC1Se7kYyixRr0IMb
9JLz74P8L82RMy5nYmLdQjkQyCl6PydyxwHy/mkOuyxpsvIbVjSjIMVsYmmNVW7uZMK7o6pG2q6K
xvBridQUNejWZ6t+LKigum7KWDKOupsJ3EmMVE/Q9h2DO03ysTJQrEMaGheiN4P2X4ualMeOjK34
6qTDiFQ2v6bjp1vLccQ8M19lpbkdDhfKBNXhVZxbMtFXOhW7kn3x/u1q9Nmm9RcGLFLnwKjZAL/v
M1YPrbws1zQ2u4oOmO6zZn1yjLHxvPU6w1IzPk/NXuRjA0P9vIZXL/2xXK7KWW1Veaj0nazgp23K
lnHEL/HzKzmDxFbWYdnCHOQUwsLcOEULuc4EyDBNVEWcGmITshVcCtTeeoSd0t5T4A56FZB7dV7R
/RvmMYrRJMCs6dEjkVRoA6Jpd1mH82DdSSriJX8OE3NlvKoy9TO8bmDeRkpGyHj1FEg3OKSRf6VN
HbuH6xCAB1Rl+zBgz1jtAIozemINSnraQvUK5F2gDieO4CgPuaraf0yrMnZfIZQX8J/Cde6g1wsh
2wYN358GusBtClURwud8mlqHpWxwVcpWysl+KW2OYi9su4MbHGWv4b7CCaLHhWfiS+vFNdtRGzwD
6cTtZBfXddMC9dinY8d91TWegD9PPAi7HrHtmgZ8fRv65TI6wthTNU5oOq9l1JUTEeFWbz3p1cds
gj0gH4m04xaEQDvTAySna5rlTnqTiwBENsX/vbNKZrMthM9R/Hkqkykp48Gg2LYPmlgi9WhEB4Vo
exrt/SdhEYyZkuX+P1MocEFWjK3iw95dxDgl5JqS8Z9A7skm8ZZs/cL65nN/4EQ74GTf1Ts2vDco
znixrv6n8NRl3FBZfyTFlnMqqdYgw2QXsx/A99c2iYMIBxCswNRY4DFewnHj1gCIFLTIfzG8avEl
CgEzgPGhx8BbvClNZbMnMCzaVPzbrtb5O9vKJHURuSMNiA4fY8ZrbnUev1g1xvHK0rwbl+F+2Ojs
6eqMqI77DnBpW3qd/5GhXbEuJBoeX3L3F6Lo6dZDMDeh8C32Yapb8S9Mf5Y1OPalH/OH+yiGTtY0
YsJLOlLFkGBwPPCA7gNFheFdl07QtoBRTeBXQKvu2tXocZ6rPmEZoRH3K/GV28larpyBdNWWy4Pl
MR5pF8kyxZ+oiHFsqdYHP2bBY4ZoFo+WcIB5iM8BwGao80RTopJwmqPc10uDgKUEWU05BBZ3wpnc
U7rNsvbdjMysQSqVLDA0kAFFKl7Zu2KE9MqMbaWA227x0LJyzkrPjLqQRJfLNhV99FwgGmtzehGt
+86aLp7V30k3qFE3zSQIzNROawlgtA0VhTuomApAVC2nwT3C4XmY34Z+299zT1FDTyGpC6qYREF0
sRgn8ErEVNmpJrJNKsZO2DKyvblQ18WVEtmJsQFnLjGvdtwCzErgixbTl6EW4M2XZQQK8yRmsBD6
bwd099/3V1Q25dJVNvxnKatV7BWX9RBUgjutz8Ln36UKWso5wu8ibEeVlx64H9QFkcmZhY9DBhGa
3cABgj+uJIfdkeuQJnnyKPh27zzlKzMG9aOi1jbBT5HY43SPEOwje/lV+BuLZIGNo6nE6aF8oS4Q
AkIVmHqjE1heuG2BLUEj+2H8Pv8a0aeDm1EBpU6VsumGkY/HgmhumgB5fCT0EhWnidOlMF3PKBXU
R3t/BfW6obgs8hHNEztISZwFdrp8EAUSTw3nMnL7Gyk//so9zMiFSFDIbknf80NrGB2Yc+AuZ5Fj
pHkcUL5X7zUcsb7mGL+bGxDjNhvok76QWkXpisJ5/d0W8ptXC7zjTix3Fm7WXs8Fn5Pho60l45mY
lHFG+Tigiwx/4VpVEH/6aHwlW7ZbHWZtrWHCAtOt3+Y/zPPwZTJixPPUXlPS9trnvbJDXOzIPqlO
C+YksgJhoZ5UUFUAITY++Pzo9/jB2afw3XIdvp0nEvoMdoW0BokbDKI9k0fBhnm4rdTAFrPOe9SH
LjadvWn1VfllVz2DV3ksFXzjdJNvnBnfaFnEeGlTkq5f52jfRJKida7rVdgoJwyE7B/nOp13cvri
ZE525ONQsBYnOPeS+ap6Z6QRNJvJbGjo5DsTCRoxd3+iPEXxzNpDdhBtiIHqPyVbkXAWX6Br77c8
hjUoPmtq3t/dRCA4TOtVIuiglQX6YKTb2tOlJpXAvhaToNqKmNurFVWigZdsuKFFDFiM1PqRXQxE
EuplXtncdtgDWc9FSN07ftVcNbjy5F0ZK3qapO1epNvcYFBHhFIe+4HDuHE+8MMdkG4u/TrDGNG0
42KnW6o8IPzi4wcM1OzyTwAyfOUkuxGNUrG3lJoCouHqwmMMdvwN4swm0+8A11ltOgl2LrzS7uJi
NDhM0R49vSR8O27CTLxWHGzzBkD/6ALjc17Rkvj3ybiU0ags22fgYb6f/7/+2OnQAqngA/kARhLH
4GIebjopBFZ9dE4w3KRgCiEvOoNQfn+NvTgOF4fJuod+V1XAgaXzHUFXj6tyDMEABOlPIlO4Z54y
4QdPsG+hgd0lSY0sktk01bB3rJj2xpqw8aWiX0Y57Eon1fjjGZoP7fXAAlSnGc0M27lFej9K5Zkn
EA3k2MF1v9E9NCb8daS4JwLeucRLsO0oU807uyT+4lsNUWOSUhD4G6CRXH/hMVaX+7XaZ2lOloij
NJTYhS3PnRjN+uIT0bFso4+Bw0QlwYpfceiDF7Nc2nK1/86E29t3tQbLMS5FQN9y/2MszRPGNK/D
N7u4IBZkKw0gHz8zYR7Du1JyUNuwJU2ag1bI+1H+8mXRC9bk3FdUyQmhbDtFE96pdQzE2N7KhnJ2
rIpDkzY8x0TV2tFqGvSIdd/TttgapHt07NBPCePmxljrGnWlH5fC5XXsnPNYLLqmKcqP/5Oz/4Cm
YWosqgdMJ6SGrgcPWNMK/W7Siz+tuhj4B502+i5Dzxch2WseUc/flo3pWrXHTz5E66AUdkf1BfrX
rTRmTCbHEpRdgoCpPZf12NyqecKHA6UAt8hZrSvXsuyhaNk9dRCsjDeSSuYfkyatfukC+7fnE7fU
lonjbCwet6ViKjHWUhc1jM4+rT7TV+rGyvhYwmoAWh2vmnqy1zuraLS4NWMzH4UvcRHrMLFhS8qS
i+5pjz7ZZ8ekjEQ2zn/iOQWFYyMb2fok29I9T3laRSoG/4i2aPRcWognFk2RTzUhmA7pMY0nEffs
djAtgbrRbscnNRExR0Gxzdmk+i1GnzM9lPuX2jPpjfLCcULtu4ZiQ0yw+pNIv70eE/CWibzRTsIq
ENJ3DjD+ZPh22d61l5508+BOdvpQ7r8oqqtQwilO3QQKUpDoaL6HBklVQDkO0VL0CrChRCVjS24O
Ecw4aLQDj2dR+yRBT1KsD7zgcbe5y1K5zo0DEN0gbuXYXXwMBnc5RKWOV8NoxKplVFJhlC3qXqjf
qRLX85qrNhzpeTsEVkDiaQ2bCt7GRq0yn7OIlKeCMpS74ZNLZ4+f0Hk5lGf2iRQZtj2AHM7V6vZ5
nXsCcR5UUiOsADHXACaIEURbS6hoNzN/agUZLd2eR2rqWH3ADf6XLg0ENQ5MewEo1JIUt+b9SRc2
+ZFsGlFKx6S5npx0T9XN5kqFPx+94Sw87JpCIR3rlfFLpevFKQIX2xTpnWWs49gQCk3K0q1wPP4W
Cxhazcy3RIzdsnrjJw9viMkF601Ow+E2w3l3Kjt9P2TYzwLc5FO7m8m9lLC6GkOjgUIsTWTT9l8y
2fEO7DGcBM+En2fGY6kSArPEmymXfstmWKeho7LzMagz2WEP8IVleDgwXF5B9XvIlU3QyFFnnWuF
QjayapTgSAerDN9XBPoYKCmIDRKCsp9fOlxzkswEAi9dy+cOSae4V+9RSw6kOqyDwzXbOstCaDm5
6tOF/ZIJBp6GZdLuzsz947wendkqbhMXudY/0dwHiptdVBnVjxPlfEbbrH9//k0Su5+4bEu/2Nxy
QRoRyAgy65pCyBJYTMsvokQJC+i7jUWmHCKpb0JfvYnyuE2Oxpr9SATD1yc62U76+IsOl7xQxkD+
t4AxjE7dGQFU2gszSl44hv6yzWsOfPu6xWC7R/omiObjon6BO7VIzeTlha6NTnClScDwnI6wCEdA
C+vrDO9ZEHAVndCRkpUNno+jW61nwRlViRdFreC3sPj6D1PZcbdpdLdYrum9jsBp8AFLIp7is6R6
E+XKw9VWdeqt5Ela5ZYpzjO2PTcBGH3II01S9V29R8D0wiwv35iHpk4pvycHx9YIdp3wzcf1XA/O
4USbaaRkS0p9XA4gkGhQtyQyonLI7RxxCTyoTJt+NDZespHf9khIyAtChr/RC/Ly5dnnZgo1NrUO
TkogexTyriukYdSVJzKWaDx59t8l52PT0t96ATZAjDPL18aXdTQh7Wvgam9Ag2P9my+A/QmGOqsW
a2rE1LgZCJJRjTYoLYP0YTO6Xen0SxhgW4kF9xrvLB+3HPxoh9wN0mtUer7uYvbyko/Tc+hcC1Kg
FrlocgL7+lAElDqX6Bh2DtkP39P/DjHXzTzPIamPAmbSmltis+EBifZ2WH/dqr772UVfSWrhx/BR
ASAtqHNCPTgDkrpeUTa4vh1Q3tTigO2DHQdjSF82Dqs58/1fJ7wDDKSJYpylScAbec3BRU+pzEEk
Hov3f6sA7OqBAHSVQgYY7dZi9vAA306jpnMnl1KTaRkbski4FwY9E4+jtovDlY6rQvpyhjFgQacu
5i2ulTZrdoWUfqk1DneeFHMbdAVlcsmznVsBmJRF6KTplB4XGS/DKMfFpYEVwW0iMPgz0FtAyzqv
g1qJG5ADcxK1OG0TUCm87tmFEQ8MpyV0Py59Iz4OVbA4TBUF47AsTwLea0DLaS3BIPFPbhJolcAh
ollQ6B/hRNl2XDO4ZSFwbFXZ0Ui57XIqV9BSIq2x21Vju6fAEBTo3+6g9zoF1TiNhNJK53Iii13f
tHxWg/LMtpVbTTrljR70fqOWaSzDjStMEn6Xn5Xq9pgH/x1qO9UE+eNCK9ZYEffOWuX+4/y9VLVs
cemPIOcoihjkRHkm9O0llzskjq7ozj/G7+4jUvrhTI8mMMkpERT+YJQBaSD3q0oqgAapBpG61Q0z
mAoXsGPBXn+DZGI8i/+ElCeAI5bjVOMY5oNdn4EwU+bFJ6KkK4oJcWvS8BfCHpftP7s/BaJt7Uk/
/Hrx5EdzK7oWnvgZrrws0ia0NBzDF2q7ZjSRWHwT6vmzCSMRfqIGNGsL+8KTuzPyIJArTtamNpo7
fE8ZjjFfNEsSa1pwgHUvOFyttE1WYDIe7jE2F9TT2ZDkB2Qvqlq7qw/YQAOxfO3xRuhmBiiOGe5j
N+U/6YfzZ581d4xuzWVtnD3saaovtWu7hc0GJ8cVEoUhMhdXrP7Li/QTeWH/q1f3hKxfP7vpmUve
UEjiLDlP2PjP5e6LFVYwHeIyr44QIMInIdgbEzs4HpAw/LocsgAPV1vQiAasMgF7CuZpQ46WOtb/
U4VpWY/YafLFL83HkK9rC5v+flKOc7MC6KFVv+Ewsd+ysTC71/4+g6v5yls4iyVrAhgtgV+Adryd
0O9xmRqIRXtWZLmS3joNYpnELeYvh4uQ72EuJi5PL7Cmzr3BbbwRbQmgqiavSqD0ar+nCx8u0kM+
NvFCqZ+zZUDpmaGAMVLR3uWP4gFQCnzFF71DkoCAZM6gdevzq40IyuNzxU+uwrWRFLis4y62ouO7
AIFlUvf5ur5gFrQcW7NC/vrDXRqvyj1+Yi6u56nl7KDFAnWUFjznPXIJFTbx3YDHSSVTlH63pvsp
EZ3O4pD5Z+n1TSJMh1xa7qgFKoe2i6ShVnK1isuZCeXqmNvmYX1/bXixMlEq5j+kPlXy2ILHiNj4
jGt4cIFgf+X1Rgyb1pvkQz3o5Iq2066JJXfZOM0+6DyQOVuNCwkCoaXxajCoIejI5elxacYue5+c
tSi9qsLhbwrj58le7DgQ+zMCEWlZ0NbtPJfbhs8CBZ6PXQVJ5cK5wXkJiWty0xASMTl65xkbgqiI
46HKHB6EFP1TQLXZfIjUc1EfPpWKnf93o+DvAniITcykgy2OoPQNaaWP0NKC5pgUOh9f2x3pvCVA
fNCcE5T0VgvqoGjubPQttz2IUQLW5daeMiHkrpio9L8KrwF8EStQ3fbTw6C/Ax3myO04feSexKkE
ovBhvORvSzpSToFdfZ3l+nihyPU+59GP4vfrJoFkM3al8QRyaIiHo5b2CGQ3cefHVNoAQlA7sXsd
bZEv4f/r3pC9E4qiOAEjNiZOzUUxz5jsI4L1t7k/Ax+e4S7aX11ybroluW2D2YvAKxuOapXG3j7b
5IsXJE8OEDDHL5y0P4p8SIqMv+N14C+AaoYOJRruk09xxpPp1cEUTezJzgonrdcaFjPVBFka5CZF
UTRLWQyO0ulP7p6RCiENdQYQvk3dbNpNCyQQzjdBrpGhEAuDmKqGtOKkc7R2Y9CEeFrF52VKwjMj
F7u5oX9WzS6IMuhv4TEIFQClP5kXBLqFV4r131MP+rsGnQLVGzWAOIswuCQobOlVtkJ7upR3ceUw
/6TZ8U01yZ5A27taFONBjAEMPsHo7J669oEm5FLcbN9qr75rCq57BheGK4EYXdDokvzdesrapWOo
rXtd5JWHeoxSlo32Yrz2H4RXqqZY+7NhoQbeWLZACzV3ubX3cmelM7DDViStvBdgctf9hdYyANg/
Fw05pDNrMFAj+DPvde6BITRG+rwhjTBOZEGUI6Ah11I7SDXr6lebWDlkshJ+90TrbPepKKBxtXMI
FRPLkMzk7pIDg0WMJVEJfq58bXZiOa5fW6em4S+rfaifsNLEJfgq5J2z7Y9ZIO5QWJ396irxOvtk
u7MZ43sS/I6he+6Otm2DoyC0EVd9DWMR33EC8ZiskNaTJ8wd7EjDa3wwaydkcsxee8cmVef0wAd1
IYd6zgeSiiR1ONIFqxGnQj+J0cxgxo+mcp/xQU7WyrR0665AmGR1w72DP9BXLKNo582UiIWlW70B
SLrler8STsXwD0E8pBaeW64b98R04Wu5yV1D1d2ZNKm/aqevc+fz4oRX59ef8veZOHtCadt0ltJe
egU+xKUeyPCC4WFAxxiW8+YVs5DWh4CUhUDQ20UUHR0v25G0aU07DXUa1+RAhbY10bNIiapso5Yc
mS3ZOrdN4wIZEj5whHtQYtpi1G6/iuj3fb7lJ0cu+5YokpfKZT3rllIOHpbd+vQPZCq1alx5pBoy
LyWDwNdEozAySLwJYYFXNDy0J0xVu7Z42UOvQ+waHjWt9sFYULd53B8Y8/CKD0HlzRhVKxvt2mKN
VxU9YRDlh075usXrCE5FE1KPu6DAI+BcYDtGeJcEZVS0RcpQYV0hga5F/PgtRgDsV+m0BGwEFV/8
4J3oE/FcuscGLcMg5G6TTYDHa4hkNfTG2SaCR4DVn9g839XTQP0UsPle23HIsCo6hC8YF77Zmy8U
uNlqoPAR1eLFNs+rBr1l1ZABIQfkUxaytRIdcjoVIYL1ERyvdEdTJwy5PeTPe1O5k0loG0jUuXfZ
4y0AbQ4ckjlhLQDZarWhkfxtfKUTp2QWlharF1+DiMDdEeC8kW8H3CHY0S3i534SuI6yNhDwxmLS
7OVDUvLmf61R7iMZgW1mjoI/DBNPYiIImmZ4fSTeHl5V1Zt16hXSvsuup8segShcjdC2GIJhOFwv
UOsWdnFmlnSW0cxVeOd4LtaucRGseVCFtyB0z2nMgxzzzUcPt4R+pDgi++e7FQ1N1gfdIADOP+gk
T7Nx9RC0WcDi5LAhkhU86QBKm7pVQyn+voJkW9sF0JweEx1U2SB637bWOp98ngNGX/zuziW+RI2b
hEULuJYoqiSv/oOvqnJiDzwzlRzmr4UiDgx/mq4UKIiXvCP4gRtbROnvwQiAnSEO30O/+pmnMXmB
Hx1XDmRh5mlNvXik3xnKuNgA/IsJIor5+C1a36n+ybQWoMszge9RcuY8bxZehfPZ2X+xBEa2DcDC
F4WN1mwI/QzXnBhWKI4q6u9/AlXk9X/Y7ue0cmxt3isD775VXNRSeyTn+bNFDHrZfjhWa6q9Q2DC
G33KjvU0ZpABszuNa8eapGdvdegM0xqlLBNQ34vM1HymYeSmsdo8hZkX5wy4n9hvnJo0xazko9kM
HD+NkH56TnrOVo2EYj+e54edfRB4tOLVzeoT/bduVJ/lz+GjJv/m12YpXlevy5lPXTRvlYKWmehV
sMcWHd3p+9M+MzNl13eO+pChR84tQr7P4j74NXsYl3ogEMhXUFaD+KMBRTvR0NC9liLZJenVXuIk
5om5uRPh7mcCQkQofanQEsgTta05ub352IP2aAwgv6ptOg5+B+bLxh9QUSjJRXQ73TdbVkV1EI4Z
+wZjAl69+h4YFr4fHMDHbvEjopHRUWoWErVlTihItjC5VHiqAs8rZRU5ZwEELgsH3WLOoic34nrt
KBMv2GeEYOKH1pblBhilnl3AhyM052kgfyoGjv+9Fs7Qz/SMYqHFmR2jRdjuhYfPtYVIH1yFCfkA
IuljtsGfDakqS2v2nY39mq/UCWiPJ+WYQmERGHh4/lpzZ+0tUo50fu2FOnASTfGH+S83eV+agCII
y5lnK53mhAVrCve4uaHmETMcE1YSZk0jsxjIFYKn32R5W5Xhzi4cNIfvz1NfCOis6LU4V6kjgOFq
3MZ+TcokeBmJ9a4crneksjG7+xWhKsrKehF3j/YFruAJAqwu9MSWr9QZqFUi8E68OHR63HFmfsKt
2drbKhae/4W9ZaBi3VBPXNh5pdrEkXoelAA2jNxLmVWOO2lXJA5y3GZIRmdeZ5xWgThZqONjBJUD
U4tc/w/q2kUGD4L00YxyttRjgN4y2vIx2Vc3IEPZcFvo9dzuDoZBaySFAbALNKoQnpeABCbcdt57
hTHDkx3T0nUrZYLiqeM8LAq7zYGxZtynjZrSIdpE7Vjg4Y5YjIMfPD/C7HhT3hWLAaRQ1X7G0W5o
B9yhZAcEI4McQonfaEe3ieD1vDXv8aHL35COQSl+U20qMPmyUTdBOV0F2dIDxI9wR04bY3Tbhbrw
/3afczosy1ZXUaaeRZsWgFSqHoerUUrOF3kKlHmQmTK3bFaW/3Q/6QSTp8B3zVjE8T4HCMTAyNn1
ft00x2yq5QOjvqquk87COEEZn6kTJxifhoLD56frg/+O1XxiFawiJsWiGF5HZWmTOOHGRgzKMrYQ
YXj5IsWK0jWHnrVpJUSo3yi9IN4bwW8tuwyAm1ROu2BdixgeN4xWoZpF1+Vl1xqxtYKQHNiLg/d8
EP+goL3H9po6w9h4+xWXqNRuypPurkqTzZh36jLOeN8buJleoVmEEtyHelrnTmE33s57uFHYtkBF
d5X3puKv1Ai4JSPw1Pqz6ruuqxyZGC7CzgUCSNLbX9LoFTHviXSSev7EjaBPrcxsqnLuDM7pkqKO
B4W2qO51kjkI+oZvssJDyrS/vCkwJ3k00mGMUbmjeCzw+Pxro8axRCypa3J6vXwTTXD8EShtNG73
NjQk0Zy8wE/y13irya9cabO4hhfRxIc6NqMqbdrJtYlOv3C5Bu+Xd41ydknyTFUeEq1OR/cpq6oV
aedQpqUl4QtS4v1SBNEZ+CpXgKqjRCgRqfb1igVHnWudupL6uZ6lG2ryg/h0DKhdvApYR6ZYE/1q
kKCTRG6jRoiQAfrpr7rU8oek4MM9IlMUO5YNbio/F7P4VK9WyDyNYVm5ISzYr1PPcyGbWST6HM7+
WV6Amq2elspHxMBF7cn3YtVkl/m6HRO6LdMLFgCGxfRJgfZfwJQKW/tvpfgnIjaCtNRTzCxRahOW
Z1DZa4QEPmUJo1c3lIYY1o8NlARgtgQmXLatQSbsXPegivUF6szvxI8uRrZcb5S4iNDzQ+HHKYaj
oumDITd3IVeA4OnIkKo785dSK4pEJfZ9NIY+SEhFOnsniyCPSWhdOZpyD6hiqsQbK26fFGvGHyzi
A5VxTlFHT2+sjdhPBpXvt4MZZSxD0mnsHC/SwdzYuVRC88Nf1v3NQsr3K11Kl+IrhVZpZDIkyOHz
V7ueXsT+dp75CERGcAaDxGn+bziEzZu1XOWVCtovayM9hsNcW/ny6+5GsPWFs6GXL3XzKfbLz/YI
EUFXX8y2qL/VAA6SFe1voopDGuRBHEcboCoE2Qx8kJWpI55kl6KZyWEtrfvGjUUd+dHKK9ZolVwV
9IT6PC7Y+5ojr27lkkZpO4lvSA82ZhZuABoCyWD/RDXNTkP9H+JevnOoxmY5lWeC0JrQtR3oGMRD
Kwa3Y9jbwMr8fukdJVq+xY+K13vjRUeVWTW3l2XewMHPDQfEVc8D13E68qsR1rxSOdAG3vp3etg4
mHhKsFBjljRPqPe07bkSHY4nrFOiyiJkbhJAlZAquoXjKb6pxuDzOlz4bsHDi0ch1NWZ9nVV6bwF
WVjOAK+bAmTuO2SbeaCZrXsoePgHqRITTnnfqdC07lzPqmArYul1GmzP/4heHN5zLJz7MUE1Sdqi
nVJtNyfMHiUfkNJyz2NdlDxIBWbvR9qRidWtZ73chVviQDg28KUzdmJx7dhhSsQf6A38tkOzRZ1q
s2qDm9iuqPF4uyEgVACye2yfAuCXVOnu5I/7n3wPP5tJzNaBsc46YNUOK5eSzvZU7OEmf77/ByUs
CoNtQuxiHoutVqZ6/EdSe1BSUdRX2uud14azjpo1vlNZo52zS26lumnZ2YvdOnpfq7CHm3kyw76Z
004TGN8yoF3bkfA4ja+TUQn/cGhHGUvC8gmkCJlnVFSUaPWbQ25MEYRxU733hXATusUDUwNxF2WH
rIF79cllmAxF4lTB051F69XxQDUONjrgnPq+BnRQRLdWbbwzHENf4NikRTf4ahFdE5GBYJiKX++S
c3TlmzDcnG6mcBUgiExGtDeEeSadpkONvmcn10gtvtVp08zLMG/mnDngp7O3DWM46/TCAQBamjt2
KgvlxqVJOZCt2RjSJzqFVtDHUbCeCNp20CGcoThsYod2igx0f8Y7o58rw4dng8RvwTZ4v2GWCVyA
/cwCLFHjjdZ9x5EViw15Z4vPEUGX/9IAORA+1ZLGZ+Z9ekWu1r07h7ONrIUNCQ0AJFINe0R6doXF
eLXUN/1aiEvsMa8N16IWbXPerdCGPmXm7r9G94WUlVHPYOCioEvrKoVns2yGJVGlLKogpqzHqVqU
xdegKRB40oAxVSSs+px/yhSOBQ28p6vnGj4JNTje7CB1PZGTxij/1QXex4aUSam7cF7xaLwRCzHJ
iF5YUx/qcNGxwb/SzTY+gHYicIhlPQrnMvsExj12EHHC5n35XMoMPOrVEUj/2IuMoKOar4rSCg48
7uaGzHdvACrTJhTy+o1XbfjLf3flhkl327ayz26u3b1Q622D0CaebJH55YxiPEj6KX5NuUy/FYPr
fLHT4csFoL/o9HxVHSVZ9sQbE+cIJF9U1lqBSu4lqXDnTgyQu5y/cc81TPVfvL3ylYTlMH1eCPN8
5vyh+uOSOPW7zyxeqtknD3N8hQn3g4PZYWJDwUy8R4X1fP8C6nmlNThudj9Kp1JRg3PVVTZBmjd5
SguUWZtE/mPFSf1aXugLSkLvnQBUpx5Wr82dx5YVFNGZBU8Bl2QY5Y8d0nQukFiO7q2FBja1dLQO
pw4puehCX7vDPgIAUZFio9pkL/xnru5zhvriTUbnKAWepkCuf6leBAGNqLlEMbHSi60w3SFRYJGP
YqNniLi4/Kl6ehtd3Cx49m2/mSfxW6hjS8hjQWTOcGq98s0BaV1vcVlIl5pA4jaGWJ59KZ2MXt+v
OCKWoKwbeo+ZfIWv9YMTllt2Px7B0s1L/+51Aynftu0a45uC1CCIxEm6xkgeAjOQy297A0xKjgBY
3GLcMtCOoBa6vYdtND1j/3xIeR841BZJ78VLOlK+Eco5DYBPk0U/025c/NKDt0AbfQiRLngjpCH8
rZ0mN9gsGru35MMgslre6mg1OcqBEBL31HC4H0LCwR/HyvNUexv8+uD/U28jA7xwjrc8EBkNVXJt
m4OD77XB+1EvZGswSzVhPJbomQCWd1Tm78GiK9cFKKiRr2W2O5+xidxbW74JLYClpg2Fg58/nX+J
X0KzAhyo3XUcxp54ZxCf4LW6X7meUGJOgMr/+TO0UnHRbKnoqtXi7hOzaS9mLI9Pmrc8MvJlY5OY
8MmdtPv89e7oI0A7Yqu3CHRhspq3sJp50luveQwnQzyfl7+hoqbgEbbprimbFtbH5PQSrMFpp++B
cRs4HjSF4f1LfNMbG89p7iyW4RoAuwwSCnE1OndUSNkuKIpYeAKhWkzXtIKTJ0zV5/di6bVcgheY
VhJwiweqpeu+Rvu0atPut9KYYAJZNrqARDFEd/Kg1ohiiDijWKuKnAtjY44nDXm8tnsdFbc43PzH
c/TEOWLoxajf1RqWbkz7ldJ/x3UgysZloYkt4XxkAzynCq0YnV7Oz5pCM67qeVTSwJOMNlHnb7EU
mnw/GukXykToW9O8cY98B/DXhoJZ8dmFPv+MxdUcaAuBNPci5DRCTAnt9821W/WIoNcsstQhklLe
9f+bGkyyoDM+tqACxEJWw3NPebHF/BKePD1M9KminzTxEKS8XeTWZgyP62ofSlFiuchbueQmTUOo
Sfxuk4vxR2G+h19GwdR90w+LkO+8ksf2i/7yr3KOieEaBPJa3WJEh/jmqrUD4VtcPkbF0iJJsYPO
+/RfSjdhBRQDwypY/T9RXDi7mkSCni7sE486o4sjVlZQQXd31Jy8UmiEcoaANyaw2/9VcMMpZG5Z
UTxpVMqdNAr5ZToCvqlTyHYmPd8fM9VtL2MNMDyrbXqZBJrEpPjLVcm9CFRaLKBQySbDcLmQQ1eJ
N13YDtWaoj8Z8+2Ig1on/nXXbUlLFyPRV/cP/JniqgdOPb8tVNNWhIarJ1a7qLRacVSN4Sk3aqs0
KUO7WgTS+ucp5EkecJVwU7/qKwATv/HK4+J9qYB60cZV858qh/R/Pmc6n0QTY7cWMFqAE3nS/c/K
iaXxX+7Sab3qg/j8Bl8YH1w9x1T+wRS1K42HnINrZnBVwsAzp8wpXdorHwMmONBM5akl9pLYJZhD
o/6ZgZLbYxmtKFdzb7Renbb8qoO7Gh+PrEnjqw1w+qeZrZWJvNQNiBcUcO1WAT4qjFWOIUgOqlmG
sZTtqTIO4nKJNVbUdqHsYZDRl+gfDOXV/68oYcvpr9HLJUwhBfMusfoljtV/S6eJ3CXWFvIXcglM
vDVuuhbxP4Y09cN9nnxjjeTGqRdyE6RD1DWSzNBAcGe319+dqXXJ8W/prFmTFFLXJ6ESmPkqI0cr
varua73OAsNK9XkPf1o8S77UdkOTeNbUDTfENIlksRr5HxykanBhv4cBdoe/Bw7JyI/fnkOD/Idz
OWgI870BuBz3vn8OCc6GymOgdwS7uljBPmBF8JSwcjA5/lvdawfBYQ2jbzjJUMnekx5b92TtDR/H
NAf3v8LvD1LGVdKtkVGnOxLFJ6EqhtHIWtOa/hUmzgsQFqtVoNPPKuk2uXOMrrd5Q9wFfpi4YPTi
qMqVP1OOcaLkxj17n27rvCJIlvA0uetJuBBiPCnzADC9aW0fCTO/kD8SHXbIopxT4XT9Cn1HHjBH
q51jiAPb9cSOSDdfXpi/zBD3rr7oPHRS57u7uir3ybcilQn0E1lOIjjeUkKaQyh9dJfu0ZQb4aUd
RsnWuEKCcXyHv84WMS6k2sXkXMTHrG5TRJBb37u86QlzRWw4pzLf0ESxufcQFI/qub3bhI1H6u6X
qM3BwaAPt0KEQuDKwLvpuDcD/r02uAHRSINxUYymrPVGaKog/TWzO1WcaQamYhhpOoXrDum81RVp
28qz9SrKMsy8IpWaJ3ERONjHnTh1CjD6eBngFoktv9bQdTIU9UGrHsoqI5WXaWqXnRaZaeVCnUWJ
UYj9FcWHYh/1TabRrSzcDkgdCPNVdIDvvTGxtnlDm92i8Fvkx6xp4Omui10739pZkPeJWvN7oET5
5aHLWcLo37KB+bksqnfWQ68PjqxGdLp/lrH7d71ljA7Y7h3tWcGmuygvvOcTREDdhrMQxXNdRxug
vs/GUjy6ExvreAGYwM58YUuf95UR8GdV5Ok2v0v52dSstB4nRWk1gS5/JaBRTNrqfoDsPCAiexUt
8XSC9XkxJp6WdnIKQjMmmUxT7JzpIleKB6DDBeUPLoAzdYlmA2xIFmAx3a6WF2knDhPdL7TDHKVb
XJC6KXRhxsxeo5YA3vusvi0QwXhqOK58k7Uc6oacmsIcs/D0l5DX+UJW7yRdkKDZWCwibJkPLCGV
bQZJqAP3wgqIe40gEbrZejlnmF5m0N1tFIg1eR5gKCM+DJABIvmm/xnohFyMI37vbBWskq01sWVH
eIntLYHTdoeP0tzDasgr9SArNLoS33eeb7ZnMjOSSLrGkFSKkxFjNXcQoHY3g622Cm/ZLpI1m8AN
CiRZGT1Dp/scgj9quorXFsP66FKe8LmlWC6P5/uh39OpWF7k9gVg0fICbfAUCpGlokVM5clVHcwD
mEY1inykt0jxaeoxhrGaFNKrHnacxvcqg3hFp3oaqciWbeh95oOoXHhFyMTyDKdfFzh5xpspeH8s
dyksiFmjDE/caoCbDC9R7dr7mvp2spgb6+f+lm08jCu1akNMk0vc9Pz1EB7HrDACcIRL35VUR1n5
QdchHYZ9V4IzGWw5J73n+0UNTQwA5d10L3oFGKJYkMzHj0/H0T1pc/NGXu0sVco8quVbBnoLz0dT
C421o8179/2J31XdhPl8z+pZKPOnCaebLTqxmls3Bmzq8pH9cm6pTvLP+EkTXh9c7UbqLawBSlX1
4Kz/Bz/QboXlmkDwj5yhf9F7YIUNTgKDtzUi6PWlQ3wByGT6UMPWnfjjv3XL7eoZDy46rzMbs6SA
phy0yMxNJyPa0xsuuBNTcelO/wy/mUIkiAr7/DObhoTAbP6V6Y8VQEQKRrVY8M3ppX56MAijrmqP
ilu8ZAc3byHs9v3eL7J7PzY3sDmrMexGRgvuTnBCbUZYcgP4KOuwvrJ918msAcVWQ9L+EbxknpGb
pwUJAv8BgFPmUGd4WqyuKJkUITABSOqGLvv9kGysBrPJa8fEdyLkEemTBc6x0KO+//ztL9XMXnNy
XICknUZ40rHTVQVu3hSES9lsjcgDOVoQ14Z/R6buN0qJjuzjlVjCA+PXbQx1vnr3mD7GGnVRinyq
ZZzsssmxyIgJATRjzt0s+cFReb+TwH5lWk+vK6tI3jGGmCr3QZe8JlD8HINTEH+VIBzH1tCr+6C3
W2dNba+x89IP856PI2sg8b3Vb9mhVfGcSzOT0J8cZp5AUcSCmGbnhqlwMeVN0dK7bQKkMflrcOw8
Ao6SmutNASCbbLakU73LfiUFRwEbTsa2iATqFCsLm6BU4Em/rTrN2mays9nyqCQfJ9oobrF0G01H
Cjfz0hOh5R0mGH8Nja8wFIOW08zmWhdHSXDqwT0eojR6wYMDa6zEKEMLYBzvVM0N2F3v8luPiYNA
s/92fmFnsL7uH/upAfIWXrF2ur1B6/xX7o3T0OSICUnlhnrCi4+nmnQkybkmt092/Es1idqb1Qnh
7O0YcQTW4t/iAORVa2J41vXI9lyS/xv7VXdEYEvRCG2BeLZP9bn1/q0cb+/RJIDRapVom9RwHXoe
h5qlU1fhj4X4tL/MoAcL1EwhbFUZ2JWdx3rKfDyB/u3ttSPyLbTqzNJtiCA6FKdFCr7cJSM48ugA
LG+u6ovBdsY8rWb6LhxbQ6T9v88eGmSHrIt3GArbzIM8VBsJlwSEUeOcg8KqHFKPbFQ3DiEBIT6E
oSDfKOwFGRY0JL26iGO2a3JNhokqDrZ8jlI/eVlQzKc2C5FvblRAmrTSXEykiUaX0TZY4XYranJQ
/Kd5XcpJaEL7zICHmUZL/d5vXe6dRIk2c0WQdSObIr7pPNkrHuHw8eJZ7yb/aD6kbGp7ji9/rSns
WvHdfeMdxAcFGq6oSkdt8lwxg51YfLpPpxDJfCeau8cmtLbtT5Ap5IDaJn2oUW41SyXOpakFac9d
PnbzQMrkLiwrNVQgykgHyQLeJaCr1IWuKXVV05BxbybnyPsDNdQ6s7WhQ/ig0aHsbFi3oiQckRPC
0thptwI+ffYxIkFfS6nt776l8piy0+1z59BgARssPeNq98GEaAhATZ7qksKvZg9G+6eBM/De8w2d
kwecY3Ani+1JYLl0lOrlAif6sbGt6SNaYIXzXAKgA6jmS8QmYGjk6kdcu/VF8RUVD+CnW8ppjSGw
d7d+7fjGLAZT99ccv6RStWJNthyDW9hYXyCTcxneiw5N7oMiNsn6Bbil3O7cqjnFLWQNwlst+Cil
zdMJqpUCayubbY5yqfKnYvGIR14r+hsAUewKC2cX8nl+q78cbFIDzhDeWxbVO3uBEQK6H4Ua7LFW
1//ZC8tmyEdYrIejAWQ4Tks9EHhyxfqUXW0OX88t+S9qvy1Z/pA5k+5wO44PjYwALXhkQl8ZT+8Y
ib7UdktafczVvNmeS2fN0DSig3G2SQz+UUUGBjG+hHxMMmKN4hQWDLX3KuqHGRLZ7HE+O3NcBHxw
UkTmY/53CM6P5/+EsG1qshar21Yp9ChjmSmbOjH7qdaGIAyNlAlng2pqCI4t4w4TXHAji/nWXNBD
eKFrRw3Absu151T02cd9u5g62EyzBPoHF14JDB2mNIs74R2v7XHhIdpmXT7KSTodA0fRxLDmRMCJ
40iEAfN5At5pU+Faoqzo03vfD3mANmaG8V6sTkE0EN3BvDZ5byVm4/dLsK2gHPG29RjVxQVn3kmR
nyJO26TFsMqL4SE1i0eleDTmJE4KAqENwq7XhgRp/+nderUnQOzXgsoLiB5m3W5fo3uSBeNAh2zi
Tnk7owBV/a/1UUh1YBhXjxFoMjvb4WoDEeLuDmVUcrj2q+6keudXn0YDHVHj+gARsQjWY7T1NX/T
KvIjiekaX1otL/IjtXHRiU9otK8aHHwwbjbpJHObIMof+zSwK088zymEfFRFwzmmyiQzviUtQ0GV
6GS2Q7Yb2WA9tt8Ny439O8XHJw1EizV8qglUwaGCXGLXvJJ0+70q6h04bJMqwZafP+IPQttD5oH7
srNHwuDKBwVvl9ago7pjqCsQV14VDqjQvgdUbnUGnQgUvTZF7j8jsMg9gva0BTG3z0e8hr4G8kI5
xYGiEM8nj0YRaRYIyLLcz4PWgjCz/qKRDZqf7PmDLwRxctUkhbA/IfrI/TE26KH42u60RqWhyMvc
oRFDfnkS5ssDungUQfq4nOX6kTPWdOp2O5Q58Wq69yGMKLUT1ox8uZXw2Dwmcg2WBbIlCIvKUnCa
Hjg0G/JOqA7R27kwvqrDbtdZrPIDMy9CtSJ17ONA+gOTOHBZK34BCdUkVk12ADmW6/bySQAJ18GS
Mstj7AIR9rYEhoNujLyD+MlVOuGFxeKZpFVsDaXtT2O5Bnf/rS7V1PAHDCoUvUgYYp2gG8GT2Md/
OFf9e7an6WFMVNNWWCYI5pZNMoAmNrIN9BWCcq5MNV8isxF3s4LYqM53MhE5wKSqU2llxHask5ml
IT2+50qOyh3TAoGGYtWbvXT+LVobyxQzs/LK2hk2xnu/rXLSQxHuIIjfh2G4aiYlEvPE2oW1fY+r
INoCZG2qF9KnJ+QXsKoV0fKYybaLK00WA9ueJg5+OrVoAthw8EOS9ONN8IEfAq3e5Dp1ELOEgKIZ
0zznZvtjbiDOto5yp56SBL79R9oThNQIAcCui/d4XMyMXhTyo3ls1QG10gDftIwKuFZbELYxJTxg
JHNP9dtNVQ19HMTL+F/u6IBpFtNR6qlkHWKdXPMCEOj579yzqm4olgIaVhJTf9BAem3iqV6Gi56u
pwPAwZMhvSXj3HL5F5NI9tZUZlCKYV0IlRZpf6lVv10U5Vm5fAdY6K4wsYnejzZMOYdNN8XP0GCb
sGI9v1HWfX+QdkMnky0jhq+wQbUYSRvLOlAt9wd0YlBl+GG9MGK/LRHT0RL3LA2y+q2RfD8VbFGg
8e8q23O4HoMHUDn3PeuRXGWhTmbuny6wnpNV+I1wHQjjW/5rhkhuht/t0aIUOxgsSAeFSIaU21VB
TptxzyJAAxJGJdF+Xj06tpdP3Fm/4wOesTaPfjQ+n22n5tcEnTPrUYRkVzvowZ7FRQggIJ2tZEEU
Gzv+Wqfb+65+Ey4IyCAqZ/Oiryf9f3hhY0q8dosf5R7amgRm4RPZjaE4L9Bg4OhveNppvMX/9qTA
LAYCst40d262BVMM+KfTArA7VT507qA6zYkqtEfxVplaAoy0wQZ4rLcQsmP6k6dvPlEwlBbnfW9w
6G9bJuODz2zNd44LsZcXaF7NO/emIJrC9+rARmEO3XIJz536LrnJFFT3Kar5epdduxPEs0Fp/Ghv
ZLSzwJZ7a2ACMZtAzLaPV04K3m3S0qkZGoYADTEkwY5aNpC2pN+gsqMf4KXFNJ5HLq09A+u9A8gj
Rs6ToSon7N7sVn10Xi0RNXO8oA2fSeo34QjRT+EGtXZwV3zkX6aqZ1Njk/iQQnRSSSbOmS+d2mLP
QOUmJzTR0NacAFFiaevA9kXAudNMdF60eY6iEIV4HmFfDV2wPLQGjaSKW6MkjJmj6xQXOLRjlZLg
51gvjIyFL369SUGh58X0GBXYUyzLrEf+4JcsfIdu3N6T5Pp0PScZ+NVPVyQP3JwxdednuTR2dyyF
OV29RTEs+mnOadxEEZmPvULKTggWWJBtlGKYoE4w5U+WFnsQ8MY+Cl7NbCcSz+Af+24MDONtcBFB
EmjUwA+3QwYnipHEet7jK3A+INtGRKBn92pmS9K+whGTIYrhPTR8MYG/SsKnUvqxMVWP1Tt13IcP
ItAGoPsSzaklWBJuUqq9XfRHBvuGPUacLQcL5s0eR8vjjHSZTomcbHcOsoSN0WbCCIQg9zRnKBZU
zbtiGZSszYwLs/LjYVYPQL5Q/F1uNIL7NNx9CCCmh/pnjF68YF4Dh1DXlr3+I9NYQNB8dMIILDMR
KnUTLjPpbtDC/1sqGHqZKgHEp/tqxXJS3ecgeJVoubUlLuV6VYHM46iQDp/cdu/fYB5YJXIpC2Pi
tgMIDvnbNBzgrEN6XvzeqD2if1bFpWCs5fElv8hilETaCYV8/z/sXclaUjJxXMtd+nB6r6lqpGFM
dp+oHV1Zxs3G1+o3Ax1rMwiEzwZyy2oxi9//cZm/H8PB35TOj4H2h+w3mSBzSMIs07N1WEOEX5/J
/3SDVHzQ/iwHWaGIH2FMnVHiMzpWHlNFhqTju2TnppQzOtgqH1SThn8D3NwbhBnmDKZ/08zrRX6j
YBH7+GbWgVpf1kUMiCbPlYU/WrZVdF/SBTahq7bSAc43Lb1o5fG2IDvSVOngpASiUB4vaVaHdSlC
V3hM/IU5YA08FRL+a4veULjAoMoxBysc+TiJJlLLGb8ITK8mXwW3duGtDBtjMJAaxZt23yD3zWbl
oCTtCdvqBwAtkproUnG8b4JmFTzLHjtp/j05H/KjPKejSATHoZatnSC0PKcbVo8HtovFzgAExz2k
nWemFPq37rbbB4UUl0PyviID6Mw1BmKjNfcqwl5zi6GdsxL0VmiSVWpLV2YB3Cs1CaCSLaW71p/q
N4gmP7xUz0aYDprg8z7nWeesidubbvJmhBtUyXeLBZGLZIHv3WJRqTzfaVaeKfbqdFSua+0oVSIP
oc6TC5VCp7fA5MeV8MlCA9P7IYnPbNNYqn9/bf+l1hWDSc0qndSatIaCezR9Bvc1efIuliilFt36
R506JE3plK22rD+20AztJDvRqxDeMuYx6Jrg7aQsyFx6r/rzRL+tKkJqW4KgGNcTifNzKSYinNVu
N8YZHDHWEmTfcnjG8rF/t675zB3GFFw0WwLWQnjTQxvImsIl+/De3u2XR+8Ct6mkmmuleoUlYIyI
7ovnk3dnpkfjtYIk9BDjXLf87K0pYrIsKB4y/GyiJruMBUwNeD6MfM85O3vAvW3yVxfLumA4Yfyo
C96Qf1oyaVGgZ92UmWeAR004jlu+tfpPbxhWr8Ivz19fdswQAY8E8+18HDcdlVyr6pQZZalFumH6
K7f1Zeqtzu2WvwQbl5eKfmxVFpTFF1DcvfB9bs4ihjkj4SCgF//1mbgKPFsDUZlIG7gllCBJVevl
NtCmxJ1fSkezRMveOOtNRtKRbyYhxVGyrMENfxjW59PfmOuZO8CwJO+TgEi7YkJdN2zJ3n2DXOM0
QnXHLIXFg5wlZxrTvgUPddLoyiY+xky2J1sDzwngP34Zh6Y3W678+zafm5TCaFBte8bf3zR32/GS
Tp1lb9dEFoEgJZspVDf/yekdevUobaEQsBpR/axtuzfOt/d2orlVZ/gtzL6NpNJFz+RbyAN/AIOz
WnwsGTrY7Fns8Op5teafuUlualTxKsabhoedRjPEIlzJjxtOpCfW9booalCDVhXmsq1e2uKPPhMc
v5qM+OsAlPb/18PPEzyTflZYVBX3NnNFIEhYtnb6nX6nPKoJThxxictTfY9yVGO0CXBYLcCQgfD+
DQpoOCNByfXKLufOGsNwUsGC80uwML+Wl7EbWznetjsDn8OFrSbLHayJkhhHzvEz9aqWPHcm0D0R
LXZ8YgZdEfZ92nRn8lhZhlpSr6aCIeIDOEHpPp9TNGTlIT8BMZe6pv1WBqUlQhE2fi1SQZq2OCPx
1pgYxbs1x0rMjY8GcZh5pq0c+sCXa7ZeqISvq3p9M7CxtFk3LcGC7jBpLhvaZrBCA89iq4HGOt3+
tAr7r9uQf8HRSCd/Th87tNDhsEqRgpntcD2CvQJGjQhSbuGhF2sSrNqMyeW/TaGYfun7+AnzFiuZ
Ok4lDBHg1kHgv3MZQOQqrrW9YYqI5FRG3drSCyDXpcZNfgguzkuK2NxREZEdI6ltcAe0uua9jJUC
Ov5yKbKCi62+H2nHmLS6MgCdmEOL1nGthZ4KQk+ivfsq8hm7WQDjvEOgKjjeSAUUwRHXBdTXhm1A
OxAfGX3hTvreAQuWHAyED/z3R51JJz8R1jcZccO9y6C29jRUSgyctRP+UF1XbJSdh1CR58dgCeMO
TZVuvR1P0uWr2+XFpADgH1HXD7mdN1JDfXTBmupVNW3CzUTscFPxQ+yWb0fDiXrK2N7FXW0Uftus
T5N/l2HNegjDehZTUyt7qBVLpKPwDumyNMyn1Ned0tnniCz/NhNaUu8/vVcCysz/au/gIa7rM3BE
aSfJLfx/iw1Eu9ypz2WWSaOOPYNnw5X9PGga2knufR9CjeOUj5JV4+kVLZtVZ44rbg+fArPlPLnU
NZz1jVsgIAQlb/feOXuGiytR8r6ieXbn4CEfb+4Kk4aydmw8W2Su5BgkRarneyDCqfmi0t3aDK52
4qYUXcQpEJJFsHmPriZUPOJU0e8ZOAHSdXbw//Na8WxYIbf/lv54CxZQCSMaZz5xaoDcV3RGU5ZA
1wCzWVt9wwUTPjEA6ynDQH/2s9QFju/JPmmHOv5pKE2R75Fl+2SpYVmFnbYD+xsIOTOzQzPfgCvp
lkf8qW+AFGxQ06woGi75sdBpaXU8dOuSzA4b4K5JVHY++ntrCegBlo2xcMxGOyTitut9e4FOM0R/
/HjCwuzSrZ0iwtVIYhb9bpUCQ0cqAibF0bzSnpQU2ywb/Gg7+ocw8/+d9kK1wprfY9QLSw9P221o
WOP9SIaxuPOG8uOZnDGSaAtpgPu7+1B0Be500LC942nygC/wZHV84f/6RVvQGSA/Ysrg7oYdcqYf
aTPl2wmyYHOzy25VqxmIgmvdxdrtqqE6Yx+aEPU73oQfGJa83r2t4DLdghQ9tAYhTGw08W0k+CtD
lIt8sV7h6PmMFMfhDUnEBr/kaE248jzsNSbfMmt4mHb56DSejxzFQRMavCp3m0bslhyS9ST8yua5
tpwuRY9qiVHSvNZx5lrrDqwVBxc4dBA+rlMyCzPFxE9ceJQKgz+suMs1jq2YdIO9yQF7hxcwKRFx
cxQ7/rvFsUh1LphPZlsitq8Ve+T9AU0wyre9BaZmC1XFgE84ZgotjNLW0wMkCoX6418KgVRCJ4SW
eRBkHIJDqQfo9oI8zzBNZHavZ+ghf4Dj0JLaNoW9laxWmRBdlW73dzS6pT3v0wqfE3vO52ETE++i
jLn7NystjamwXqFTOwsvSjju+77T72x7vJLHNCzeN2o1YL8Ouo11o4un2NkKFROe+gCzeMDXWuKt
dfBCL6BMSUNL7FXAQBYhQ2MH2WQADEAXRb6KkCQrEchsoZHV5UUthzp6ki1H3f63fxkIbENPDqTi
HP2agDjuxMUO1Mzr78iS45+p+wODFxmckGCAiWuJEnBW/nVvwY67z+0ZIAhIZschNdcUAZuWBdTn
q5FyWRvDbXKR3HEiVzKv5WJ62BTes7aczhfY0lQGyTLPWO26+6i5aQBYcqlMS07I3mo4DqQBZkYB
DyXitNNFutDZedImo0mDQsccqlPl2qNgIlBwLBTNgBagDpjGJ3YexbtTS9W/ficNAy9uSyP7R/f9
MCPu8TCuHlSVZYfVg8pVlezzsyOnXnbbqthFYNpkPXkurq1qxgxRrq+8p1AkMKJ6T8wFmo2VeIzy
1qN7crMzsXDbXCsL38wtofMRZrOi/ZHTA2G4ClsvAtzRUwSDkSxzq6vuJtahM7LpKu4nwKxifW6w
XTOZTLVk2SvP91h8YFQZGXENyLM6hVIUc5olHqpXBBxNArM7cJHlvv4tkDLatkr8CRC4EsxOKEcD
1tB8Bx2nM4hJeXIVMPi2OWLO/hwArOrqt0+06xeME16vaZzsc5VtkM+xAq6miJ/osm/vCWb74M/G
+0XGC4vy0N/+O0sSnVMBPLnYcNzGqsLiVrFQ0h9oJkjdS6mYr83fZUsicKYZKF6DT95AHbjJZw3J
TLLUPg/9hY+r+h2nFeAPIp4SboehSS1162Bpb6lxj/dF2ZwIGSXUVcU03O1J7Smo1lP3egHL9yi3
J2S42ZUDwCTuDwWXmjeOxHe6a0gs+qziFGG9cOSbzDoFQ3ek94WgaolZTVGP1nQ5QE9iCndEwzZE
56WRFH8LsIsYBqXS1+WO/LPrWZSI1qh///WiQleW9OdNntp2Kb+0mGyMBUgERmJNJnIrxEVWVVmz
BwW7JbTZv/exvT8uCqj/FJK6ObQ7HucMe3EhsGt8IkO4svfs+G8q/jNate48BwW6y/D5EamXrWqY
2qRzYh8+G0gD2R4TCcsHpxrXMxQ4ttmn/KzvdpdzoUHFUDXFThQzrpF7u1RluUqwj+ZrJgU4tlqB
H0UCms9diBVxeUfmH/4bu/IgdT6NM8JFA8jU7ZEmaZl5OhZ6o12cv7MnfQCpwj53YjU0lQxmdCr0
CHvv/yuc9yhOoHG2xWS0XKKGc9W+gSlILhxxU5hV4+jinjOQbxAPw+R5YO2IdIjq5OBgrPMz1m4L
MpwMjGMpNJv3iDZ1f7M1zLUmsASAqGCRgQKjVX6QjoHUdtlhQN2jczKKLUosFgqQMbjg4jsQ0Wgy
p/gp90bvhA2IF5U6wjeWCjXEmTG3fIWexJfMI4OHFMviwl4y2qpbkJqZQLW5+6cvBIgpMLNTiHgv
pZuq0WaZKx1YZtWKDWz6pKnX7gHccIY8NIHNLnvzEZeECxbznW9qOTwVds6aYmHkg3WIFfUOlR4c
nH7uJUuL77WqkgciHmQcXiY6niN/jccgf8dhv1+4J1a5APIfpYUChPCFWhish2RXemQVrg29WeGY
Nep1VUcLp2jeK8VEpt96R7U2NEUq+hpFqhaD3lxXc7tIRLAMujgxgIIOQ70Nvy8vr0uTsJFx+a3g
2sHU2VxB2ePZBi8DOuADfc5kKT7Whr8bS8VoGA12fiEmfWODKX0tFuSAsIqHref9j5H0Q/LZkkul
3jjSn+TqogoqKwyvpMVMVDG0ZvAAyqhgBTMmVGdcHjcyzTBFkGTV5dw7MOpSilt350/a73CzeFLb
DLRyVo2nZoplGr0TbfFeZzqInWCRy8KN7Pswu7W2FKVl0tewjxICIuiy/qRbeRySSURI1jMAn0GE
3oHlPiziDBRrz9vGBybWghSd08Qy7iqjxWRYgHwqpGm6X2ggXyHJVWPnsB+kb7lu4iYIAcMG7VqX
Q6qrWQCjQuv/iXR0+lXOvyVgBigNI4At9p2frBvQNAox4u25rZrGfLNqgCCB2qKcqUfyYIs1GVIF
SYwjC2Kr12Brc35z2QIvRS6mhcasx4nnxDuiCVCaIMxDGo9wNLvqVLMXclNqn63peMpwYdJntqo2
+6nMk3U6x89JNy/vq6oRk/WemsPrMbx8E1BsofHrixp+9k667snSNi7dhy4SmiEKyxSBWvnMXl3q
60guayOarmS8iW0m44hNR/E10fFCnXfC/DODsgMWunBrZU1xU36saXU2A69iI2vxGshtNDleFm6p
idtTD85Y7TdwQW5AvyJp9FM8CtnISVXCHzC8SiJnMIMXPV2N/r/PnySW1m8EoIynHTNzJLod3aPp
4FL926Gl+if7aNu66+BjRbJ0xgyhbfyrNjGujW5SnByVJWoQL8sd1s38AhoFmV7DflXWmP0kYBW2
+5kcc492Nh/RErNii/h9e6PWkySJ9G6g2Y4IJsQ7awTqqmFTtPNxrgwreznUT6NkAJ3teXkrT/dg
ylbFGM7ovEtLqQqYdBeYl3aY5QwoISm+2u6q2xJ9dZzkBP/vPEc10YKKlzty5ZqA+1Yi2qX+0u96
TZMQpaQ0tM+qCyZ3Kjd7/ZCA+ATgecyUKGiHv4xhKBSUfAubIYs9tcpeiuqxWc4V4l5a8cxxzTDE
HAbFMoFXAWFA+9Pf58i3E6pVm6U8lznV6dHMMTQOJ5lK3adUtk/pQ4Da8ngrJ5/IWNkoqHiUcmbJ
gqcOU8xK2PVzMBpKwlcKrlS5ZI62doCe5JFt/9FfmYNSmwwvLqqh432wi5goe8TQ34r9RmA4oBfX
QOzcKsJiZq+P9EdEcZZxcs4bhNCfPQtfa8sRC7YB+hZs0rhhPDUDHQX/7bDLeQKOB0U/nWNjq+de
vGXFWl7lO0XAIALe64Lm+PR/bhi1c2YyjCJGPFasxI2GCA312t3brWKIM03aXiho6u8XUSh/yQ0v
2Ua5cxEsKfEads2XC/AUKQDMOUvdNFYCM/66aotffCJvyZZ/Luj2TT0LmwnqQMMdU9Tym1yw1t7s
Ba4rEXc2Sk+EacNY3WNhygCKYDjZCB2quZ6zdPzbmSqqf+fBVB49PsbJmvls4Gv3DDK8V3UwPL58
l3aZGUOinjp9zfHRWfaQpr/wDvi8qOIk4PIYXjgZ1w5Yg6olQqOZQwxiYDnN7y54Kj2oeUpHhUEz
dqBFlpPa5Zp9N3SCDN0YQ+BuB/F5XhNI0znOxsGIYrzyKSMt3arUKT5M0952dFKYMgxa9bOM03we
O8jv36RzfBrxB15UKDblrHHITGvhg4MO+lMYCyDSKSM6PEBaKHwKBW7l3oco5BViJx6LdLfSrf0T
hDnBIBbVjiFIlk+O9i6wvtn7zYwaZUkBWDdzAm5ckhlsz91K/ILMndlFRBs802GuDw7Xyo74Sjbh
dsYFltrYvTCj2UK3hFqiiuBvhryZUGYepczZ2UapSBHE4qfeJmAq5UEDau4R872PmMCGDGUZg+/f
tkRld7CBI8K5+L/YBM6nolrnyxiA+NaWJRNnsPBM0hsoWwyW3YTpLRAVc4ilzLAOL9SlXxDJZ7wQ
Ma6p9JhkAedjMfwb59B3sioU6sX9LkLLfEAnloBAK/5W4yiuBEnIfqks5j4OAVvHrnq5BP6qBZvh
obSBi8RFOGRl/yEbPN0BfLKT1CmGje6DVcgYq/aPpsZb70/8fXNSJmHjlj3yDrzPjNlg8EUZuV+7
njwk6+6WeW1De1jIWL2El/JgmU+M1eja6xFNk9W9LR2Xp9qeiYF4lmjngXFBYGkJT0unGSCsHak8
UmsvZ6sfNwTb9+zNdFsHnKcxGUGuW0o/jtLXuMFfRjnxEGAI83bokuF5XJvP7gmEtyK1d8TS6ngn
dSbub6JuM+uqTRyi6tkE3IG/gChNSFARikMumkaGF46EWPSmgu13/1mwJLfr04F7hsAyJ4ubF0LJ
PNkDVnJzMZVsMY1GF6HHs/+N/vLZ9lmtlZvZo1pJcp48Ha1A56CMxewfHOPds8ZhD7N6C3TyeGiz
87opqLEqMY5v5FxgkSL0CHq18OGv+vC7w5Q2PSNUia/0VEHfQKxkDMgOvM/M5Xq+OZyawdKauozG
xWOEjG7Rf4c0Krl1xAegY7FxqwyzgmmS/QbDYd92O6a31rPBE19ADcBFIypUVwgBZvK8YA4cnqsA
Hc3Dbx1oXHiyiwWuijpL7dfHIZZy6yI8lloD+Ys3sJiQqrhHfUKspldqFkhlzIYlN0wRECWKPvxo
LRvVTTJYtBJywduVqrblY4Kw2TwamcOnprzm7DePpGiJ5uIoLpP4D6odHfQ5PbyoUly1USSCf8Rw
52No7VTBh7zD0iJTnHzB82qbkBsLGMjjKF1GVvonO8YoGF4PRZ9bW9c1vuMUnSnTlVJQMQP1AKpB
/WzJDunDRNkR81QO57shtaNKAGs5Jt/+9DzKddj/wFUU+LxJ0qu4o4J9UF7nGqDUlFoEQPJq2EJj
u186JZpc2ixEv7aafjMt8J3I/R6V2hVtuF1AWaBk/fLZNSwPmi6AKY368AzhA+LZNfRpzL/aRc5X
fddhib5PT0JIOHrX4TJoOR1vjkFNVf8fE1MDzuS4emWK0XQ0NaALio233WzKhSYZoMAgLycnGykA
mSeTiMKa3o4yTdNBU7hdj4pI1bJK7Glc8HNr2kLrVmebTHiW3aZN1/ocgDRXkU/p5XVm4nqJfU6W
H+9rieDyUd7wdWSEJ9baCZVlKjQllPTeSWKkxendttx1moAAHFYKTEfbKzjPmEdIHHnhuZtOnxOH
6y0k7J8+BattvB6fCMmUyy676ELCtWHlKaDNa05IN/szvHKAOUbyGOuNr5m1nZJ9K+YQbIHtu6g4
SCeiLM+m18wvfSUOHa+ziuXXbTDcn8poYn+9pvmo6S7PMZg4OtmTLSDCcz9HEo03Ed7PqIsm2r60
sbLwtnoEvYZhH6PS0phL/KL/AlF6wEtHoH+xpoQYGqiQnlzr3nDOzPWI6Iw1nID5qD9HvFcEzzOZ
2w3dd9qXU0dzRseakwgX9RhiSAcVGd9JxfLhhqVWeRrBEfIIeVF2yuQ+VIahjp5mw59yWmOYFLAC
Qm6mFHIB7Nvs5DUdRyl7nTDmfwjfFQFOfmu3zo7tsx6KdcBf/NFeHN5UJAvnUpcbEEuM9GNowzeS
1Of/UACOqGFBY4urZEP+a/jQYXlwe6a5YwW4vtFiKhLAk9HRvUPRxjF+UzI5Mtj6cgu6WJUOaLm2
AYH7s29TvXqFtOV5A9ATk7CQyntyh/9IxxOvHg3WWUFVLwm0rgvag3OOG337q0YTpAwFOQHa+FiE
S0gv2DQO3So1JwWCuzSdpAl/HZZ462fqn91NlcS2+2GCzh+Tmrpp+7jS07r8oR21aMUqIoOHRgXp
JoKA0r4upTEYUb2zBggtqx4tjP5JEKJkthmGQ709Y0/BfxzoBBD+bCDn3DWXIbIV/2PhaTQ7+XDU
Kgc+lPdXENM91FYufDDh3rJImz6OZp7jhFhfDCf6kQQ8qQiV9TKDmCYc5k6dL13IW3RcBf29Tvtl
QekMwYh7ZOQzEadFPgKLT1VvlNRGCFroEIwOyLHlmI4gYm4zibQKhubRngWQ91qrztuhBqthbRYq
gz1kCRDTrV6MZX3sgEPwPcvvgWR8Kq3yBT1qK7YoN3VorKedmAoqDU842Yw3PZUaJP0Pzz9Ncm3X
326L4OMq9VTLVNmmSq00+GH2tL0A6/Yy9Z/x5Ge6SZ7Q7n4cC84LMHqGN2g+om6RrrPb+XNJm+Bc
LxQ7x1XzB7Afhtd+Mvo1ERspHdZtnx8AUb1ytDj7xn2rEPOqTAn9jrZ5uvJxb0ya2g3iBx0KBwXk
3wfvoIxAW3dIhaV/3yDgrfXuCSB4IgSeXISD/d35nEBqbltRsz43NCkbfwYOR9Ow+6xrdcBSkTVt
kO671c6aMPQyLHTFRQ/iZFKnfhS6HCx/y4QD8ogm7QgRArBKXCWAdoQSk2xF1ExixJLRKX/wmTqg
MimVgQAtKHFau5+G33j1UgZsnTl8izjQvtg0U3wGGNLlvAY1zPbvZZtPC589HxV2NNq7vOjdL/sX
4vv6AA8571u9RzzishIelK5ATeKbAvXWNddWSAzE7sa6N3660R0ynqT0aXrgbiOMsLYWxx1OJHmT
Ki2pILKtj9CyE/ci7KRjyJ/ZFrX+SDUG0r2xvd/uD3du/8sg3IN0F0RFVsWONtOf/HM9IGs/9QYX
A/cVa9gx+Hwl94wTKRjmHJFbEBPF8ywvLU/pXRTCsCfFNpUMYmL+RXi2wQT8swsno4pfsFAR3WfT
qvaqJfWlRUSK/zXGyNGKD6Sy1/m5TgvQtnFOsijUSunBNH3zJYXP27Nb93uN8m7PaWB5DQdmeOaV
s++vHU2LGWeOCzGybB3fmBh2qr9GbnX8Pv0hviVyBZBt3iSi5NiJitn0WSDp6sz0lIPV12lZk20A
+QzisfF6t/Ch9MMNgkbARp/ciKTO0t9PyHLKiykAWz2o8d8frpwZ15gvKA+WpJaX2yjPp9GyHKJo
5MHyA/gu0EFMe5+yWFCrdJl52J7onWI1+5baDKpJFK6ibfRQHqU8TtQrKpjyfUXJP/rDLpNOHE06
3C3qWZOeVlI7KERc72FCX+8fq3jnfC1Rr//1LZ8ogSeckgDogcMZdSokgXXbQRvffpdFvldtaRB0
aK8kNQjE+fYl26czWFhz6DbTrAiIVS4Vh1+Pwv2Rd4tbGhCrdJDcuhtcmj2cGmmXANzUwMzxdYsK
OS57P8HhtYQNkJ0RlaOOin5jZl947u+M2l+l83We15rgtajdHYvcqBzEaGiEMTg1PzulrPejTKdK
1pKqNnHMHYcNYOlunK4wUYeMXJmfQ5Ac4fvzhkGTB7Ef88EAHtEWE6YyztoWoE4T8b5Am1GZyy63
y2Xkgo3JxLu+Uze2XlmhySU5XpAmOpQq0mJ8mPCLf/XietQmfavM+aEhJezhrDyCieRquQuwvnbX
JVjv24S/4hVD/4nqJetd/MiS1Xxe9hXBS8MVJuAox3F69OwM+EowkMFj7yUxJAjvB170/JV04UrH
logz4G5Iwn1rVjJxAwEgA3Cas2lo36+OUnRZE6BoPPvILqLicmQHo/ENwZ1TThL8Ge8XeDnLgh+U
P21WbGpKcQKJQHFYTw3qj6buyJzLex9rR161ijLrxIyQf3WZqoSwCOOSoH/VvBIcqsdRawP/ENcT
KqoVLUOUS7WhFivoXO6Niqco9+puGJifsx2bmAgoflgDCfkoZL3O76SHOKNcbccn/bcQj5Q8ZxqK
XS2oXfC+HxUVdkT+aXnOqNDGyIzLqXA6sHuKQ8DmZPVwJKP2mBi+dirMn8Zmw/ALVz2PHMsOjKrA
c/iPDMt0g6JwRKTwYIF9Qw5fJrUFtqXq+XVS74kDyUUK1t+9lUaAQP3jcb/4iWeczvz616H6o/JE
6S8007B8+Z/kIZwnXxTpEMqnaLWbXKTgwBbsRuSspr8muRwDfzWN1sGRF0SkusAXHMktWtX/EAfw
7fKRhLpT8ZWLvYwC5Nb4KZtSB+O04GKf2x/8PdgtvCphWp9w8215rkz2IjR6eGpAAdxKJz3V+dIt
KQI7LGiAOGvrwtbcxHD2Ox/Hn+pnF3CGd0wnH10+gVe5Sfx6ljEDP3y/rylJnlVc4SPmmPZimxRe
Ajhat+xXQoaRaIW0X/vr2O4bAm5ZMzsF/bktTJc3aFPhzO0huGOG9RZaG1Inxwx1XgyeEA1n8pKT
8hSPcOtTJmXiJhaiDP9F2EHDYLYesiXRRxIjzTD0SKAV9sQq5gSfBVfYuP/c9fX0fXPNWEtCTa4g
ZitdIqVE9062dvu6UGk2sqwka12nK8jWmfG9hEJL40Fx4C43v7zw/YqsjkwYh2kWHaXOaBWF7W6l
MkukDIXInTA6dJt2lXZnys3IAMmtmLU2jLA0uEknQVG7D4QatfOL+mK8Ib8qsYsIxBI30uqER41+
PMzwXjwLC8PV/ozHbmE2STnjxAnNZ04BFffW1PUV7DR21O1LyEAZg0gsqd/Y+wsoTPnBHKRvZo5+
Fl3+f7S3RN6yK85uljhjpRaPfK/GNAxRLMxwiMCS8tfgU/Bzb+R/+v5t8gExEX4KskuhvaqCGYjF
okkQl0HP3z+9XOkGKfjq6ASZZxTSt9FnY52G7fVYu+g6SL8j964rjRi5kiV+Ksg6cYhbd42g/Xxy
jqWHgq/VQsAVJ3Vwm7pGiAiT8AX0fxyITEziXI/68ZkcSRxFcPPL4ipAFTS4jQlRX8ffxbSafsnW
ez+1oL/QzAdWrQ1Srxbfahb5ECnVrxt+92vc23GY3If/JrDVvTwmQW1bqfBatmDG6XynxLgtXIoL
kio8gwJzBAFNvq0YnOpUV5GXm2Oyz+C2CQMZSBXg9Ab5/epZ74mq/i+yF/78PMdN5Y4MLVPV6FbK
urBODhtTkXIHv7GT3dSI0WqM9Pe4nzxhtfj+PXQDP0T3BnHAJdA1SAGmEO5DKyZGNiJx0xoB18Uz
z3KGLIGo4yorbRXmvzklsV8ChDTJQoZM7G+ituol82moDK4SvTPZKvsAY2SwdvvRoZ65eOr2awF7
ea9kb+6ARk3MVWmjKDUy06W/dPNRKQnQygkQkWNd59EwBJAnPTBsF7N5FgMz7Ho0RbVDicdQyCoN
B/N1uUxpTpefrle1s/inLg+A2xNekxve3rqR117/JMhYPPpLwXX6lhBEG1LYLQ0Z9KiaXRJSZyUv
5Y4TR5SDjInIHzVIp4Ivlqo5beKtv/WZZDtwhwKpMvb4TMzcxpqpAzMXefKI0qgBPaV3/g0ayeuH
iJNUEHep5iWfOD70NKFhq1NM/45youXNZddoVmjC55MK5qQ0ifoVI3z3AJlDhIHnkQ8DgiE75FYZ
VWg3JCSVJASzX3KgX40Yq6x12ZXYcleBz25W2fXWLsR85mC5wo4bKNYA66IGMuQlC+KNtOwBWv22
w2pGa2fWt9siTMvuzGHAl7AO66vcnnLzuwkF0XZOJtI+xHsFs4V75jUxJeXl9pgr1/fpUGEV5gLF
TiE7f5DjunGapfX0oHnxCBDiB26gbBXb0fk6nc02WCMSn7ZyWzH+ctzbkKtZ07FozwvIzLek1805
AkW12zpRGi3X+HmcCfZe2cXFh4YnShcjotEpB+NDOLchLYY59Jvjt65Wd/CZf4rRr57EEONxz7DA
p6N9lpBOsmKy+d74XE+CvT0GDY7ogMocwI2A6u+sZieK4lApUqSDd5B4E3GSCSuVkzDWhgjup1fW
ZkHenocrSxal6j8UOTJeMkx+C1jtWkHbAk8+/v+DnCd9D9EStPDxlXpsXTOLWJpDN1p+YYMJBdRr
uRJSkm/0vp5Dki+Uj28S9rFxC/ykb1EwcOJ+CDjQ7U0neWczvmDZUqqUWjcn9Vv6aNrUH+ngZmp+
XqaxmxzK8bVcbOhG4+H8b2RRThiCnUskpa4URjQuus8OHMNn9Yhs4cSBmPXT5crGC11lGoPimQUr
8BszeqL3FlWhzYKZjM9LtxmdfXQsUgFPMnjZ6WklNHxddLgj5XWyL0/kTuUAQBdjC1EBomVUzEjI
nvAQnFRc8syl8eEaML7fh+IgKl0EgBYprfX+2rLAyLttG9qUx4/0Lt2Yjf9UlGps2YqRz/WmRF0F
xIEAuGFUXyU/aFRQXZHdel6NWtA/+7M8OIKdxR0Z0GhSXlZxVL2PRm7JicqXdV8mAQJRj9B8LzY3
ukMbv26iUH62xe9qC9g1CS9sOSOLaomnRqTDViLj3cDBd9Av1WugpUTcvXYhXFcdEKCev914p38B
caRbkmjbue6dKPHD4TPUp5/9fhvkN8UiGBgL8zNXBH+jJaZOa/gZ4laAIBH0fC3VXfHVnbLpUkNT
xkFQFRYKapEz+UBkZBBQHCFLWsnaRn1nFmCjjV5n3q1McC0As5+r+k9ZD/9saGMICqOXi6y2Mhj0
vesPC20ujYbIwlUa9D4zxA0Jv19BJj2dXcD1cxv+65aNlPwZyd3QDt8wr4SInZkdlQQe8WHqsgmC
rc7BQKUWsBC7tZsjIO/ALSmJDCNaku9kvOzvy4nE/+To/L7E9N7tzP48MXwBwafPrB9GvPqoyKUS
abz+tVSrRQehLX8oxEu7FndtJ7yGQ4QjDyP/bTWQffMfFJFep+cvjbHMuPtKhhQ8mMLVuvudia0b
8IZ9nCkZDNSK9aiEiH+coA+VTyJNhp1PzB5VqaJW7kblRgL+VyZWmMvDEedbZHM+Ubz5musifNHU
R2RBfjUvoAEGyU18eW3RVoH0EkBPimpwg/vu+z0pD5yhc/4pYxoJeyUU+rjjzwqieq3A2IlNqxu0
Bi65Pam7Ep37b08tX2R4Nb1txPLzFb9ELRDVne9QTCXRxKCcuruDh/TaLB6FoxTIx8asqNhMk9TZ
YBbKrb7xdKWnhR5egBfZMydtRzwJkQI/DnHVUB9PXKNBOJ65ijlhx3k9RMACG4/iP+5BECVp4PjU
yJSCvh09TqwqiNlChvwR9N5JDIvBGqIvs63SThGzKHn0fUrExYrz2z7B8/ETGToqaD+7DpJtQhwz
aoxiKn/MluXuHRKw5nv55ZOxiUus1sis4J6izYZPwxvnQ7I3fUG+d3jMD/NnaSB09P0PbMBJsfUo
Lwqyekk7JK8H/Dn8HDcj29nhagCDY40zn2Yazcmq3CVqG2Ok7Z3gCQgMkei07TFUP82g+BQEp27P
LU7qwByFATZCr1KLPkLVL45b7fc5ERpSFkp76V/Fx1IOLVcUBMYK/nwSTTMZcKmEkOOu3YiJY1Iq
nj3GavcTJMr+ZXcrx+E00jCYW3CAwt2JoCc26xOIF0C+uQf8KalNcwoRWQ/ufyaMOvMzSZ4+3nCL
pLpNZERrJ2vwgEscaXhSkEak4ddp0U3AKKd4vA3rTdwnG+DMKKM4s9lcGx6uRCsdL/n/el66umly
ocU1LQyzp964uvev6MHXIOSY64htyM2V4d5ArpN9dJZU8dNgXId8knohdR05hJuCMm1N6Yh4Kz1r
B9YV4Qs/95kajErxjrw9f+fAFk/GNnPYqN0HCk/T7miEZD2h7fWlraaoOpHiPHuBKmLj9KldK8w+
40T6zyDevZ7mX6DW0rR9q6UiH+LLg0kTh/Zo9P+xAYYMz6pvGZYWvnHfyMESIJScd04z2btSnNht
pmk7O5i55/Pv8ARMIkuYoZ4UFrCspwsmNT/NG/VK0zDMYyoWX1YGsRv7rpSMaeZQdBpCfHgrpB1E
wCpW2v4uF6oBUGjQkbdcBnhfaD9lBK5MNy30Ndz+25xbys4D5sPowYZnrBfDKyaqtdX8T+9KUqGj
SykrLQzCaqMpzeeYliU8sOvhNRrlMJalQ4s6sNYNNTB7AIS7DxZpVN+EQEIKbVErp/zmeOhoA/oW
DV1sVtrqBSg854M2QizLtGJwwHYDl3SeELwFVNUahkN3pELcrt6Ch3EZa+yLty9MUeHlqVDGGuSA
FNM1qjnZiiLiZDFmD9BWYSMS1WKMdBMXIWRrcns/9+w1uHeNpxO4efrARWsFQx40P7zPX18sgVl/
ItcmLFsrgaQ9ahMkt8KV/bzNzBr0vakrRLTcrJOYi2deNPnPB57rOanHb58b7g/ITySosXWZ79aQ
P1DZ6EpY5+VKGZGllIx4ipZw4nrhZBlnyZTqFkZkamcRyfwyjUFka9t+JzS9mt+h5l5PPskBuTcC
BQ9EEinXzN0+ApKWQO7Pwvqngy1H5PHEb7x4dFkIrN/C6KgSAyoCyyi70eEAx+GeLRX1XWxbbDkQ
TtSrKulrA1viaeLP+CInqIaE7Ka+qUbF2l8W7riJhjzjt3qk+0x7T654PpgmIQ7R6dyaqLUego70
yAlK1YvxxWQ7jpJUnZP7pOcc8WngasjJ4q1OnOhRDiO8PfDOiYz1Hy/sEBKR2nk8llnZlqZbjIp4
2xQApwCnUrXdN7tL2le8p/4JWgWOZzQ3ZqgtVaHCysAQtjgcWlys7SDIXsq8HR4LarKkf/sRRD/M
AcrrJgdT/5NQsq2YArMYlEY1Qosk1oZbma22TCbacbnX8IWLH3I3GuX3Uv/yZs7k9dUlww5xLinY
HOSxrY+Jz5+bLyHmC9xFRs/VbD10DOCapPGMAEpmLenIcsbcNXp5rUhfep4QdrtLjummmhSxRmTH
94vTzMAY0JlG3gy/i1JTZN7X8GQZ+x8f+6lMGIbYQQgcT30j+wb+RJAeYapIeTfaOnY9ua7vYJKE
F2ELTp3dMIOeZuHiuWmyQ/8AahpbtUwmzOcSGSvQ+Fi1b4TEjwbZMG/AG7PpKalPniqHr/BzTsBe
nYJVS0Uw9D6T9qRXgDwQAPmURS37V8t0lmWfEQZoas2nDGlaM0oIphM/VxS8rBv7W+s4ZT3sI8Gw
PcaiO3LUp46Bz6q/HlCLSo+gIO1UonSDiW9C04BkjcHfh2eAW2sEgsq+LEYOPb2EgjkOjfCLVZ8A
B8+zg4qtIguQCqwNM5rd4Atj77Kh//tnxdtG35Oy2rxb+RUHVuNDHN5f2yZxKRsX3QlQdRvyr+Z1
RIbXmdMiYAY36ZQbOF3d4YAqlpBcG3qwC/qORP0Vc4Ya/Vzge+fwgl38NVwVCJan9y/8KdZQozgK
DwUXAnrDUE9ASELAEhta0p9/yzdCs8TsVrZQaUREse4z47475OH+fWFnKtuIL8c9zEtqKX8W3+5J
6Zg+Bx/ultuB3mknAGxExovw1MWp7R4YFJFscr1NnGYMO7BoaRjuVvPQa6PI9D/2Khq1t7eFclRe
6U9YxU2OK/sh0kQoBxbS7bcnQaZe18tTIoLQpCTXkFYGKbi82ryBwxXXFPU+1/4Q8Ct5QMVosn3w
JHRSX+zmJHBjaf8FA6dJWshi3MwfBY0daVd73LC4p4Pfw091ViXJOa+uvctPe7Y0rOPRsLHjyBlb
IWa27AVTd80WxmDYIZ76kUQzJTvWiF5CDsYpRC8gmEkKPvSpdwgZ7PMLmVDhj2C5jWiS24xVenNd
iT9DRr6qLICiJhFP1v4/DUcufJsIaZr19ndLpZVYuTr1x0ewnePPR1jINFbqHlPnagJIGo6AF8Vg
Cacs3XlFAOJyvaB0IinPAb0muidHZRVkr1ke/+dMLPg/bpLH8wgtQovHald4ylIWO7Q5CRhv/qQZ
kYsgO+Kufe9Ki7dZAocM31Sw7vOJiNK6BTsAhjjzNEjfkzl292nNzrX/r7U4Tf+haeSePd5g879u
mgKT5aAGAf7nJ3vgqwETPawiwYr5duwls9KFkP+JIL36B64WZkR+3p7mQjCgsnjKouST7x49B8DQ
9euWJci63TnT/EB/BjMDCCj/Bm4aupC0sgKAulXaWt8xaoM3L2+jv6HREXtVnIOnz6f9cjlDMPzE
u8c6pDH7qLPWHc7UD60CyM61cajbugCtnS94xW5z7pCf+cEr0lYIwi/K/OuitPEy8n5WkZsFGjhQ
nt4UsKHn3cesBZ/vGiLGGgmlw8KGbhnuIdtivWjjq4fYMqBO532NQmGgyXHZtAxOJ/jgEdcAAG0X
ybtxx1APXqSL3aW6nmJiV7vxI4Jayktvpn0JMo+A7Cc1yi4THKoDYaLTK3qd+ygHU4jG+CC4hJAX
lW9MQpCIqzK+8eKzpK4+ZlMTkOSyzBMHEsYkiPyAusb3dcv6AlymKnTskGgUq4Qa3FBNUQ/Eer00
i+hfLUf5PekWyzl/GSQaSQVx+uw26a4li9z6q4HKtKtpHY2KqQJFlK2/E+cu18seoWQO2KYCpQja
9QC3ULCTLmdlPt99E5SaJPbMw3bjayOgkcaMH6m+JK5ja9E4AkqZG9BTXRpR3Ldc0jO4c2aWdMmA
G2Tq6f0Kny6Kzr6f9OcUUtGWdyK0pMNjUiuV3yNItHF1ylR2gd3gNBHYMRMIXY/vcZeqxVL1Bm76
l8iYvqz6qk9hBCPO1B2/9fve5ZbWwIr4phBCt61csMe7k66FudC5klir93kG7XRPIrJS5Tt9lBV5
UCDxqzjD67ULcM/EKpGpC9YWtCNJ44HnHAXvI+LJa4DvR4nEat6jRdKkECKgf4WKF7KYI66voCby
QFTNPzDGsWqGn3VMu0yAOcSMco2sGfBlkVH0fXZ9uKjhUHUoR12wy12e8u0RJEW8VpiSTaBraQcn
P4nOkVrLga/AVP+oSUuS79ER2pSKqotvQ6Buj97jaJqetePZnJNKvGnhXgAeN4JhRcrCA1IM7JZb
v7auAmwN0eExae4TB+LUiWo+F1I+Gjb3vJ4MdCmkqOfVvdo9b7+WnWqWWlRDihwvrb/26oCB4Emh
/nhaqA0fEAVPDj3C2GgwpbLKuebTBVpEY59QStu2bo1SP6r6+mAZKKMmneiumen1+S0MnjjVLtSR
R+HTypXEmPaB6qsoIqmGQPOH3MC/dMHZZPuIlu1ddg8dbJuX4SDuklmYA/fHfQshOEIDWoxJu0WV
6qrOp+8T8Fre0yLCtWNzS88kc2rVSeJXyM5SEkpANLOoefyWlfZ0PNfMvclU/NHFTQHfSL2cCZ7Y
vVFYguU8M6AKw0NvzG4jmOFHL0gCKRrD9UsG/+LulOtuM8BvghRZPFA4GqWW+MvmSOon5iuQHMT+
cV1/GHhZ6LK6lbld8+Q/w6WNQxktfNXQfaxy+kF9wE/8e0wySvYIuag4Bc0ssWqEfkMYv3LnPN5/
R8OCWpGh7eYWd32wnERLjlr0CftUCcVLZhREjHgnQQo3urdvnLl1XX1DOmSzQWB0wa5BQ4/eu+9m
e4EhXMvt1mn48iATT8AXSxEQn60BFFBnpNcdjlqSRFZosFnDytu6pYJwDAPKkoNORgsCqUzIBOfY
BpUp+YJBRAe4EURE6AT7+GmoHFZM/t+1nBANv1rZ1UYd7wwBATvgLEfG3wq45zKp85W94CdG1O71
POi1gzaNKaSNVm60FsHEfvcUPaKjRv2zNgRLfa9OQ9TAn3X7hJVUiDMwkS+XQJl+GpJzxdCdsP/L
zVOQemDTcm11sFHDxDHTTxrPMrO+RxQGJWKiY5X1M0eqRkZp0fkI1kpvUFr4supjoJ+Pk5QZ4Tl0
uJiJ99I0+NVjpmgNjfD08nd1Ig4YtzaFKk+KXsPhm3FAzOsArsWEVPtmGogFLkmZ3iqBApc0lRth
s0288JzCuGj2Lqu5heaTyWHb50w0t9Ua+potU7Ow3NqG2gAbP3e3hNYkDjP0UWmswQ1sUgyL4a4R
uTDGcryWNH3/Zcuo8hQFB4ZpNatk6vhGfy3pdoChJcjo2v/K+d6SQq991oZYUzx0Aun2dvncwzuy
KK7jmcqUc+HjVZ6dXiBllo5u034og/drR8XBfG7PqFPdrarNzsPx6F9OiqevdZYuK8S8VdAZuauk
CNW1bmkSFMjpJ+cU5oMTfZNQiNkuDRz/hEFQUMU47t3zXvmzfbvQQ3MPhsrd2s6QLcu52OgD3jM5
nVm6cYwq4hWTTcYu+TTIwZgYgd1lXS2J1ggDSz/KlUsRwDq5Snl2Ae2AIyIk20dQulKhu0s7NquF
yHYegXj3LMpdPqE0ws6ZWvIQwuQQK6lLCyjuvEbyUXECtASTxeB5ni5v5DVnFiGwenNNBNCa2Os/
H3se4rdvU6tH4yYBiiGxUGbAk9c+vXZq2Mb0maPE+UnIOo+//jZSJOFlPFkWb4J3pjOM7Z6rlj/O
LAAvH7VPOQ3GPaGDCrQuiIUrjv2jt7LQ6Y/pfZyWO/hgKvsfMi94ummKHY9k5KpfJREgKuL1W06L
6bCfYhZo49MMH8i4O4kdmUjs86IWsU30RU5CDmsnnHZenv9DYUrwdMxG0MMRjwiuAM1Kw6vuO76S
8PSQdJM3yHRM9NhBxokazlKBMTpc4xoC1grAG2t7/oEeZOe4prCuYpMFOn8ShrmDfKYNL1zpCy7b
gH3z2MWRFHJNpSDTz1sw8grHucCzCUOowut+UEdKxPTqYWwuzEeM0JzghKl9lLRhZT9WfeK+0ACm
sSYKTMFQi4ewwK96b5S0UZa37+EGQHHOVfp/mfRe9Z/sewdIEp+FoSCSr5zVX4qR8Pe3mYFC4FAG
GdwsXTb4kvDhiMal4bouCj+SpKy2FYOgj6k4oldqxrf96n+7V39UYi8PL3RUGfKEYJWaAjzclbly
65FOWG937l/CpdsgfbBgZKHgeqP9+IfE6SHvCV8pImWw5kgl23zqcVFgaYIjbciaaZkBc5SFKrC9
+ohYhI4IRHIY8tWbM5qBIhCHtKRBQczU038PCp7XfE1Kl4PvW+Duw47pP63QGiLIlzQWoa4LCjfk
eB3gxsvI6zgBu9DvBNl6kdtQKrvRQG1D+aZKwCs+V9NbEOd9Ah51niDtnPUIAZjoZK7GVcfPqKH6
sbhh53FC0LbiI83LxnPia6unbYo/CPW7VD8dsLR8k0llyUUD7qDWiwMhjiIJhVW7i/ijayNzu9oh
AQmPnvJuBW4kJ3gW5giDe3wUGWPbNoV7MyOyoP8tQoHMRYlVmkewxZWu5qnAVzemyy7tHDvHgRN+
/eahNuuWP6igEiZCLBtYG7BEBX3IA4qlIWyB+joKlHIXcSYWJaes+WP264ejS2LV6j69Zo+6GCGQ
rG1HdYYuIzTX5+MsncqmqhfTpNkC/9A3XPlDU85zuWq9r0ZLqK/EGdXNXXAcn0J7fNkLi7LP+oNS
mfLxWaC19wCbGVUrcRQaOGZkE018otb3dHJEwua2fndzG19tU5nza0OcTpS/BuUUvIXs+oQFX52b
kheoWwcUI+FEMOfo7Ea/P2jRrs48JxhRRLNjTUCSLXHYSNIYKNqNOk/+z2xAjvch1Cm2PQnGyvBX
bas3nETgEsrNCFP3nYYFDE1aKG9RQC6Le1CQsw7gMk42MQELmiR76aaWAjj+iX0AimraE6y/6orh
Pic/f2Zzqye8lp7q7UUp8jIAsYfsWKyziufyhMwaDiGubtPTPn8an81767Ban7otSN8Cgr12s6WP
ARVQ1V0tLtJrsLGglYYnK/Ty3B8zbyI7ZclRoT0CnnNPKUUpYGgKT+cqa4Apfdnk4hFs4SaTu9gt
CwCuilXNnPIpzk+62864qGJ7VsWYY3brr/OBUvMuH3ZCrCESocdQHjuJwH5BBH+l4auciiv7d2kS
sonIUzQjn2xohX8OKr7hajNgmHjspr0k0yDAdq06P8UPC62zatgjuQMe6pwYkkOZwpRD8I/KvwP3
X/4tROHHprywnNz1QauWWa/nfBRcIduYad24RCqgLHgAMTM7c2aZqQbMWZubnMOt7vAy7+frEmDK
4aBeXadhI71H0rlxdxpw25xxZ/zO4EyJDVQYQe67yKJB9Vy+iR9Xlygf0VOIBKTFy5QBfChBd3Dt
mUEXNjMoMQL17r9fxaTqk0rxscRhG8ZnS8C7pktoCH63XpdqLL79EbJuz7qDzmwSVdG5T4ceEIpI
tk+8/z7JgkH1dIuzkKyjkjFOV1nfIofN1MfZ71sz+umzajCGE+xs/5aBfs8LboDvxwXTp0HV7etF
UI9G5uZzvD3dtXrnTiOPWdS7RtU6Hd/TUFfrXrmUAcFkpwabOJGHH7kAt4t0DclTHrwfYvwBibxY
IsAkmrCHJHQPwR2flixPPYT1ASDYvOScsfFalHuC+vITHn8M7Ei72jf+K4DTwMQOVxW7UkJL61Av
3gsj+78PzNl53h8a3JOpM2ekcq88H44qDKtNJXe70eixTb32QDF2R8nJG09tkzAso6CpHL4Mwm2p
Q71KUrOCY161LTsdhVQ7j5+zldwWE2T+MYgTA+I89Wuqgl0pMMqrWDXSY0WmZ2Ujp6OvyM2ub57a
sXIlYDsKmPlFrGv+mSjCIpPT8ufXHDZmfCTbcslc3EK9DFlTtQZPGTqOYP4+nJqGSbFrq1JqkoOD
2bj+gqbDYoMkhdrcOkSBJh5L7DqhSQego8TzFE6TqqprAy/ZmxXXIlBVMRrGxlcTOO3jsEm4KfiA
4E8lbYkF91ZkeojKI6UssKJZ3MTrR927j4GflxKnkuftAp7J5pJpbJ1PL91RNsxWctPDvQ2zaaNb
1Q+Ir6JzELMJboKEySkcTUjSgvzvUJiX+VUmNdMhSSZhu+j5igGiqdb27gu7y5qJShNWVpfq+JX8
eXjKuiUQl6mD6sH3gdgk0LPZzvTqDLL98liZQD2aQT/umlttiT8ggXRI32reE9FKRS20o6I9QkAz
AatkDpkscZGqLT7sRs1GLpYW0app7B2I0o4Lri/C0JkmbafsZMmXp2aBKwXqh9mFw9CurNZ5itSP
f4qsO637zNJ065HLmmVeKDg6F3I+7JcO3QI7p/QsCnEO9h90B+Xlet2n+RYG1oUdEBLYLJgLkpOo
jgJdlEaliOc153mIT9JSu4g5qClyA4HolXoiCLrChGdwEgcXCtWQ5pC85+X3HoH0ht/XC+oG08AR
5SXS+umrOHmfEmYgnv0gS2r2WfZu/WFHY9MaqO1LPfOR5Xlo6EDR/eeHQmA1i65S1y8KCrGBibbW
JsDUvRoZIKpzyxxtLbfCZWwn0kkns6sPHsJ/8Hl5ioLgWiKCAcy78j5ZNEaB+yNJz465RhlAehUJ
XdDx5GZO+ADf9dezDltZ/i+7UK1luJ23PzKZZby6JNwKTjkGiTWoSMBGpY10dL2Bs2NofakYxNFf
OqLxVNB+bbgYoUpgrFTDyksCdZgiGWqyMmhLZLmhriHWcNqbavOe5dQvsElo0HFRnAOOko6Nq47X
NUuxg7kLhDQ7gDWS70sFqSPU6ho12/8UUwXZ112CiP1DNh7yn48FSU95dPsI6NpetkccMO29vtNN
up9lki0s0ip91qILVp/6AakJ2a+HNJx3wp0U+YGKGrse4w3eaYzKk024Cd/0JPz+duK9mcqcnsQo
xxBStub+7u24sFz4zeWstmMmmMzAfJ4DNUXn4gXkjIgRNfAbzwfWegVMqk0cgv4RtOM4ifVCI4x3
7jcKSWrdARdlUwBxyTOMvGrHzttiq5JJBz1ceDov+ZQVgDz3CDDQme1oIicM02K3UHUMNA2PwFqZ
4cXmC9dBOd1No4/f6/EmNpob95R23m9vm4P3Fw8EgCGrLx2VKEQv5wlfGkOaNZ4tjNJXNuVStoTV
lqeG4RB/xGEkWYp5DrVh6fPIzh8FMGt+TKHYB9S/CkTguGIeyvWT0FqucS2cCiRf1hdZ3geRS5gM
yZSL99nnzeF0hwrC6pXJaDG/HabGhWw0YPc8DeOaBTbtbXJGZD/a0Sh6pNo7gNFYq3zOMinh7FOX
yVu+n0HbUwwcGle3abRRf7ZiodlEg/ZDn0DBIwa+/OMablM948a6AVtdJFZKMoeHopLtuVvRnhHC
Gm+PenH2zeScvoJz9U68RdgFuykYFNx7ZCdHWRxB/sMZS7ggfXWOahqt1VcWmp5ElYIJ82G91+KO
5lfNcmWNMKXTEJVIDRF0R6jvcf0DiGvxD8KsGnMbRiWtkDSehELkaGBgMYcwI5Bml84l2C3XXXmi
POSZg9YF5UhT+nao444/m+//lxj62EcpsNpUXrXAWVxzesWCBjDnFxr7tQbFOVpdeBF0oW7EeKda
oquHZr8LIySJJb0yANNSM1WtwkqOEmTCZ+NIOKg2s++eBidtEHJ0PwlVKLwjbetR3ByRkc9V9Paz
eSy+uJ/jtfaGXzhdxk3ulUVGgBfMddeIPo8s2RukV+YWZKdadP+Ff06yu1O57Kam1QVwGsJEryD8
ll5YPJdnsGn7hYp2w6Cd7kxVinrHt/xmCxSKVVDkL8443NkiLMgkg/f5DLaJHoxqSqqJStc2x/SH
dtHuNYY3VzLB6VX6AR9YAfUvv0E6wLZYZX8rnEU3HPVYHm3TNGwA7gvit6ZS6L/lU5GUUbsrkFPF
5YphaXrdd0lpJpelIbEXoEfZCB5zIy0OfnWqjDdmWmBNQ3CU7eMcBH2K/MzSDEVZf/DR/IMAPeP/
IPtcsnQ7gcfMBj70DszWTzNll7q/S+savVHUzutxWynrDoZWlkicXhMGWXIL27ToWAEf7MmiBx0A
0X5O/S6fBTvqvHQB1I89aeIshd+KuBCvRdRfzoAGmrrtTEWptG5iVGjzqEKxjVe/lAFnrdCxwaiS
ZuvXO67tL0quKlFQvxdHm+qldGjth2nvdVFndCoBjyl1C7qEm5p1uSAyk4DRz2NaVdCb1P/iDMsX
lwuAzMaalvs5TeYohHWJycKesHA1lH5GFDwQAGfNyBrP/06vIzXMxP/bkHWfh96EnlQPTrx1M3FR
cF80wScfIT10AajvyHatdvMi9zmisKwpAbhGg7hfCfREYy5SzKXhH031N4Avc+kx7XL/DPqAu/gP
t3oSxULGg/Z3C6aPg3AGXO196mg2XDWxvt57v3En2lVdYzvKK2KTT8avNDfT6OX4qy6zHWzq3+et
zc9cp3O5Q2uqfcbUjUiZ0VcXfms+h8ehipBHYdpxRPEwQOI/XlOqB6k1A6jsf6OMFajvmgc/efaP
LQ+oY/GMcZuAbCMhNUeZhUAk9ellOSuFgdahihugiV4bxc4tu9xS/1r6V2zFBmKgdWqLdlY2TRA2
KcdOAQdWw3IDm2t2eQnXrL5CXvaTvY/z2Stz5AXHZcOxjSJ07XKLwn17taeh67PBXBZuSW+FLk3G
I6+mth8QbSq7wIx1fERy+I1K4VYpQaZJlNFY3Wb3FMVjS7qRg6WWHlMCNH+HYwTj1VQ3ZPZ/2cnt
Ft0xXTWDOxKaYVvvgZU+OumzniQkZidXCsNnz4749TTNPeNr97OSvk+fwreQslIFFp4zlnf7B7WD
FleAwYrPbmN8+EaVSJlMLXaqnsUH4tjrUCYUJ0oXcc2MuxJoZVvUmbhejcuymWRKhRzyKuYQL8Y0
o7W+8nC+yai5994QtePstrKbhEYjR0mv+sfS9h4zxSEHRFdQLOGVLxIgDFcAlJs5naLC542u7Gix
zDpgiXijYe0wUu+IiIrV/c5g+yantJNbw7obH+cuPeaeU0/uZvMBV7VrKtKqnkmiO7ZhxYHCMyQT
3BxoFbKsnMUNO1LntYJl4TW0GPl/BhhhAm7Vfn9XtFJ1GHexKeJWhps4uowBAAxw/WmZplOC3h/x
IpYaCL2gxTkt6NMsRIHn6cfpFJOik/5YMAwvmI/2OExBB7UHq8C8AtjdI8ALbFHSARtM/a3FNlQe
JSMrvA8CPxmfFG+DIt42xENlNL36MnkkGI8ZB+S5DnJDujbfFIXvnEA1mNiYcfQ0l/1SRRX6BHef
KtYt+v8YccLcZO8ULEyjwvXegqLzkVZLVMfRqZl+S2SlHx5AhzOzmMxe1jJV3CbnDzGNEtqtTZFa
iW9NshLYPhZRN7vQ5AaCVSaMov9T4eogD7n7greZ8EanVJLTTVnJIL2lPbZPuoPQOTrjvYXXn9kf
FgBHhnW7BbMM6Imw3lajWRroNL0VRdztl9RzPmjHvJ4syapL7tV9w5V/hBfrkiMt76z4CUeWMONy
AnTR39B/adqYktHiHdN2c6OmimUgmn4A4HcJg3xP2vQDjprHtAn87qnpS8J4VF1CE6F3ffk9sl+8
bZKDFHGypjSWa4c8gpFXbmopkPpeA59+Y4mOqbmHS4p6HksVsIYxP0AU9tZ0zXLVwdPl93hMLjCS
cBGhLxW0okLg9R2Jr9YhOX27k5B8C+Z+I/2lwRyRanzu8a/HiYSfcaA7ZYFzTlRiww0ds2b4s4mX
H1VqEKslqkYRUCNNKibY4T7TC/iUQNBtvNDgGSqzViRY38XL/X0Ovt/SuCZHxwj4918J0vLbd8Ub
RsQkOGSMrEDTDudEfL+lkoFpgl1Y/zQCiMlM1HdKzz2Fux2oM9nB4IBWPQYQdoYEqDlP4TnDAMx3
aSkHP7oi2sZ4tS4ZVcaFlSP7ddPQKZg4GCv4Zri/eaJbGFsB47Mky7iPgBXVBk24NZQuFLMr93rW
czVnX6ch+OPpchuHFeLZciZdA/PUplwmRaLbVOF/iuEf/GQDfBanEN2NPqbdHB+R1dUm0adRZVOk
oPXp7LeHu8/9hGMzLfekQYjwV0Aj2szgqdWx7w5+ILtRHd+TSQp1t9BJNgpLUSRHMD0SF0htEdZd
JwiIXFUyyxamuKEu2j28aTdzHfhhMWzvOrHFc4HNNOvmI8OQs3mP3VmphJavvi5zeSLAGJH7aOyL
yrVABSLbhvT69qFDIYUs4O7Y+9MYC3tlUAGzZd60x6viWyA5U923vptL5s6HcoFhTbCsmxUGtZs1
dQpX4HUBF9rnAAUQD5jRIoxWQC8ciw21xTrneo5rXpOCxqj+8LVb+E8wOcH6NAkWWCzoWYZWOgB2
jZw8sPZlye6iBBsCBkcDdlBblPu/wZCyL6YTeaOWSpUtAxIPEVEmWBJ285+/QrcEFKVFAkm4e50U
/fIBIml01zSNSh/4CCdw4r+xUWo3Z2D1SgyQxtUam0XhROi/LbFpHK5QPAbcpG0PwZFNiXuVRHWt
OQXW1kbVMuwmzXXUxiY6hIQpYy5JSS+vIHO2ZHYhXxfPvuqw46Hje8YdJ69Ygw7N9GaegIlJ2pzf
DB18LrqXamDyMJjeHnkeXJUo8YWxe/O00onYcPfvKsp2DsReBWf/Qz49y9rTSl6gcm/QFSdBFLba
dLqrEtkU3EJV0Avd1x5MVYLfovIUlYg++Uv/D5a9Jguu32s7p+hI9Rfn8eeCbF10fh2Ty4RMVW+F
vSflrlsOC1RkKucIFeZ/qSK1Js9bamQ2o1aROy5r37fwfIbkoALNYhnMfpO6gQZ3WoVAs/9N1X7x
AtG8RiJfEdBQ2iLAgCq6P4jlrgWIZVGLFk3dzaScvf7iGAt2kQzar3917L7qq8GXMD56IHgjChHo
JPqVdQufvQnj2MVn4+lqbqVLg6+y6N53qFupNTFwm1LCx+KsKjhGF0SAYcnDpOC8m5swcSTLDb0R
CQepE3NcsYt+19KGbKVsrjHhhDW40zZx3B39ib36nK//3rFI4T62fHbaQSZbGUorXcpg0zoP68ti
5ySgXQmkJ+2FmpUz/jey48f/HqYGZpDnb2cRYxEDLstVX5g7HDH+TvFwbSXetJt4owVcgIIPhI5o
EgsAB/fW4cGatDsmE+0jkoWIQOVPaOi3EExAtQ+moHfxTDek5kYObQw9ELZG3Q6YQxmKLy4kRzci
TZ0I1kl3dZ+l+WDxhbH6JimCFB9W82OlgA1GExpevfnflJSqVz9otJKpmsuALiMcFt8R8VRlGFml
10Lxnivq1/oSq9CaFZY+AvvdKxvNNYnJAeO6hZMblNT9JTE8aZaUQK0KcbhOs4a5swWgue5lUxLQ
bw+3fZNsgioo2IdyEPx51cDV9zGKafBryVKH9kqcvm666fgKCFikF9hZN3FnCF/bt2T01Z8tSfb/
l8AakHyxwLzm1t8H3yoqVWtdSAlANbC2LT5WEXEPiY22Uyy0HdP1K+fHysM7OIR9Zs+LsJqKwwtN
ytFmvQpxcxvZMYXCxjifdkbiI+BrX3qCM07d0B4wLl2Yu92CSLJs5cx7mI3xYXcs+s8jHkpJEBZ2
nRcoFqxJHdFKGhGkeLDtzxEPGi6ykIAMvGqXF5IslbyNp/twNEClRBmFo8eJ95Yz9lubfYK4lTCF
cW9P4cs4cV1MBm04bzP7KmtnpYpPzH5emes0h5bkNAfPL+g5lQvQpy+XiBMrfBmO5WNGvXZu8HNb
j4sAdaNDZLMEyZHJlDskFlAEz1b/WMFICmWe/lEwJnt5szUgPgEjSZ3blYw5q2C6vahTVLQ5fhzc
wD6Sx+C7klbctVsOdWsO93zdV/o7zkZyUqRngsHgfnVeXC9khwJHfajwObc0fZiSmLZH7NKIkoY/
FpepXwUD9F/L+5AA4eg/OJTRhSYJpmnpiJ+w0pRXeAXyS2vh4nh1Aql9pE3YkL4HzSC9+QkiYwS+
PbtsFvll6kzo/8pBCe+22Yb5ho5uHhe0xfQsBijvhWKajQl0tcJHw7hrjQnIpRbw4djYPYy4mOp+
nKR1v7EXwUio+NfI/2Mv4VvSgXexwwwKI3IImCGKQTGOC1940NkA87kDue5uzIPDA0D/yp2osGI3
+vIFvyf32uG9qfWKkwIJaZNQzyjbKyOII2kejb7Hp4fi2LMwH132c+Ov6bjLtiGVNtlg0DgRhyoJ
d8BLWqmSEKswP/2r5j+Hd14qbgXPjMuEvnyq++ZeIX1slpWK/q02ow9jUct33JrxbN2MHqaerlwD
QBKPV0jpsJj/ckDTiMy7A8vZBU9SWFOzxvy/QoWPP2VIH77h+B+eD9gY87PLaVW7Co9QA9bXLDj3
kTHQD8C2qJMeOuE7SPbtxn1MC5zariAxsxuOezeqKkdtAqCT4pA4df8HX80IY6/7tOsVuSXokKkO
mpxjHGuxKF8DVGStliQ76wwzmN2b7WCwtD6IPvp3st6dyKXCm+ALWwTnGgpVeL+FXtzUxLOO+6eq
hW6vTslEOq+jI06Zy4ALbb7DXjYApRd301ciGz+zzgzSBGTY7hw7A4SmuLyH1IG1xucdmdFrerWS
ZfWyfSlXy6RZDgyLlYzE453HtZJeq0BF9lHDu3bBtjmreGeJJlpQ0Nd9kMVXQ87RhgQ99rFsk3ce
aQOjYtQwiqRsgG10mr885wg3ZGncjEQHHoJxfc/tCDqzQOAQZDwGmiy746wLkUXrujw9ZRfpOlzY
YqhKGGyBPWcc8SYztTw4H81bj0ypvFNgkhT8ySvikD3xjKaMtJwMBb/Qk8dzkt8gGQC1j1EQWTSE
icXSmF94DZ3ReGwSQJ4LLCtFsBkrPNIHG60Z+bVKMG+I7PAccmQ37ZFIN3WcRoXLXQxqKHPJTHrP
mAk7/XYROXCPEidER+Vcdv9YuIcaqXBnpmfWTeCQ9UBhhSEuuG+cCyaJy+WH97bTiNfggUDSG9oM
DmKIcSyldJtZVE4ROD9g3aIqWLCkhyhFojDx2KwVDXJ0piGdqp4/bOZM5lJdh7f2+ktq+lU5gXrL
fMaVu5VtSZDbCF6UrZnZtXAXaV/DDgiA8F+A2xzJRAmiFV8iQBtx177/oj1hctGheTJPHSd/iGYV
FnoMTPM+zEGHVHulYLqY4+hAqWGnlrSnoEZg1qQ80t8eN8qm6XA5EArMhBCu9KAkWZShPfHtjDAK
cGZJ74jJPPawvtxR883qXz2ZtQ5z5GMDzxLp2ZJ4TPMlm9G5zZHs2rj/Un8eXGI5IwROU/nGSyqz
ufdztCvdO2uD3aZJ2+goI2McwUMYi1Dy2++Luw0WoqVot6jSqATRb9tt87ZRSuPT0GrAGumy515l
PIJsjF06uptmzuuak7e8ro7lWsYUlZn9362DhI367DhP212xhinUziQfTh+txvCFNSaIfZveqyME
WdpzppZ7uXuA/c5nCsQGE/6xuArGcvKZ5ZLmmOVKYHnSl/OWpBIJdurLnbFqa9/22XAvBGSKaX1r
R6OZdkJgc8FFOdWXUdUMDvwgNTIYKGiER/0//MSvyfX31AF0DLl9+CNL7Uk+l43RoL8kh+Pz/PDS
6uG+sTKs60aAYf0KrEGHVV2/FABo4MhnvcivSze4SQbIzGwMVl2dtb8+E4CQVFr8j6ChNXWjWASG
o1hXQoIzCLyLM6MSkzKivBwkKUl3K4AcCezDoS9Iiy0JZDY7h0kUKGbpT8cD+uVjKmBfhyg2NcDO
E3x8ng+WtFWD7t6uAZ7alkufnSqB8C6irttZ5RD6LymSOIZtK7p0JHGA72cMOOIK9JrjDW6HFsCS
n88/64dhM1ZhVQE7MxgEU3VVkY4M3wwN1RBjLITvez2cLJWrt2pMHKplN2hpyZ6AzR055RXGQDPe
Ird6KllFKESq4Jz/JZMRBVnfOtAd8Waz/3N5vA6Coe/EsYByNnKnWuFL3wdyGBg4c6VWLSe6wvJn
onjuUs1x3rWbZorT+NP4xrrPBSLywLBxAjqI9/lB+k2dfztHe4Fj6uA60pZqroDY4hcbx5O29HNa
VnssnLCRBmiwL73mMpgnSXgBihur6DjNxZ7ZVLx5ey/EO31yhPxef31xRBMnRflYeX3YoNDdOS2X
4vHWHLAJ8uENa6b+vz04lzokFY10a8FRkefA26eGZh7q7PFqtXBhVEUiKz8RD4/HXVRpqyBRBbMU
kjX3sL1iaqKeezMm+e1ICVdujPQJ1PdO9HdMHkz3ci3BYS9vnCBZJBKEdTCIuhuasjgzgeDrY0pc
pd8nRmpFSAqcvw8B+/lhmhDvbYV8wSQztLhfTVxLCJl464SGOIK65C/SUeV767mkZsiuggW1HT1p
Nn7WIgOToDY8VCXE93rMuX2vlkmRGb9a8fW4O3jHytt7B6OMmn0VbbJ5ZNcAILSzc383Syo4YkVp
fIzx32xNXl3Wt2UltxAjpbrNIo/RrEqVcbOkR04TWP7kNrokeagwmTR3TEpmVJsDppExr/RDIj3G
cP67GzbnPvTcD8e0uIM6xcUDdIinzZg2lFAMHXBcz+zLg0YXWaVmjTuAOgJK7JIxKX2vj7/bS8lw
v5e+3jZqO1qdrrjbvlY+AyO5IzfPAGgqyZ7zXi0pBHkMXnwRhcAjfMYMPJIzds5zfUMdH6N4Tg8m
O7dUmKvwj9Na9ph3jbyMFXuovJT3xkGtyOxcPC6ekmvWEY0LpNLWdqxgUcFk5NNLxIGG2xqdohZ2
8wED+XSJ7GmeLb8hR0wwesZ8R8bGW7qTO3cshQ6+SAaK5AYd1LrTT30BrRrlc408nT6SFRVJcWqQ
jC0uQtSoTMYy0cdCn18+WAx7pJIOVvplWnyVI7gcvp6N9up3Be3H26V/dKkR6TGmAYncMrAvhs+T
OJw/KPQmXgZpEO7Px4FC6ZAXKSvEVLjSokofWLVhJ9vBoPQuG4q1yLmcc6LDDbIA+OgCSxlUYuF4
JQ75xvvnhs31S9x+4WqW415lfwyetCo3k7/IUWdiHhISyH8Zh6R+8g9G/bT6v0yFawY7fxm/+x03
GlxtJLQIfVka0g5S7fgUbPSIk34/IyNLP+HQ7dO4iv3msbQPJH/UC21KGb2TdHjIGHjkCLyblCBK
q2KRjx1PwSO2FmC9edPQw1Qtor1O7nLKzv9mq1jCyBZz/t1pAtKS5bFOnW03pdZxXAfrsGxvb/kJ
Oa1+QTyo5L2Ofpk1uZeIIPTK+AzEWcQlPKZUBopOzU7yLgiZTi0JAGEFCXKCHf/k5QDdU/u3FtMs
SZxn2kSlD/tvWCvw2L/Wh3n0kP3q2hVT82i1T8N3GtyCapB58XlndrxKEoTcs0Qy/Q9xjKAb3FHO
CtYmw7gh/rvuJgK2YkRpSHtbzQ1o8AWyhg5drNotP3KfCmjv12ceiOPlmGUUWGDZGSw240Z/BXCo
H1u+/sXQHUheMaIe7LfPJpmKnbk7s8VhKoEfRLUdoe98NQa8Hzxbha9B9b1IsV0TvxhdtJZp/P8a
MLVSSkmY13oRYnClx0+KuaDAQlQiKZxXhNJ4JpH8/1gg5UtiUHTfbz54jNcs+EaYmMZg1NoJIe46
7/xaWA9GtzBzS2phXHdAdLGyuszDEEsQm5rYZAH9nYFKVzvyrWBeRiKWuJ4SD78qh7j3Miq6D/xJ
fx8R8b0C4zyWgKNEi5LAoY0lmcdT4NseaA2IdTRWZsLoMDYFYxowRvJTslRE4wlsmeOcapveBEk0
1Afomw3cWLAsHKVtiAH5vM9Ibm0YBaICX7i7/TRIC3qy6qRhG9P3YD9c7XjlfY/IcADIaZrdui+j
3UqhSX7LlaKNK1BGVXTzhC7XYLTlNaumW0Vj548M6epQxe08f1Bv9BhVZIMLO5u+pzVITBhqrDE/
SyiMHJdif8ybv9ZQWwKtMs+ZFMFlVgv01mK1hqm+wWx/y0cyPPOMZxHB8W2+2SsQY1n2v/1r/Umw
+jWY7NoMJ81RWw2aOpxCyHpzC/UQR4SeHKZC1gSceIUYP9OW1OX/tigVfgFPAMP+MjeKbmM2Jhhc
UGJ41LHPz+uoWGk8xnm5OI1V7OCOYNLFEYzZWRC90mvnmNz1z9PDLqH51DpQcNGvY8oUzR1rq8FB
lZUVYWJQpPo+r7Ah1uccOgGOX2CHCd/ti661creY1YMb6TY4xUMQcKiPJ1BhMZaiBaZdVF/GhwQm
tVSOqLGP3//U4KL4CKtQ+0OW7/3fGgiToyPc6YQrw6US6SQsNyMHRhSemnPR2pb23XlpLxhQGL0T
4iuBjbVhBQaqa9AdiJBakhTzPg4O+BAwHH6VJqgnpVKPSGTqiSi9f/Cv5At3NchungXGIDYV+RW7
FVUXA/xM8SZn3L9y5wIH2gfRX0DQ1Itmc9ym6EA2jiiUw4vZUhCxPnPtXudq5GJ875EpuxBlqG36
hPUxPTh4/Mc2hpImVAfBf6okgTGFXDPYuxQW2uAPkRNPFPEHa4CfMBy+rupzo8LhEcJtqRp/gMec
0dltJpDESkQLDCvMG3Z88WMMCmhsen4lBoRR9FFEjsiSeQ/KO8iee/yYAe0QsGcxYcxvJvk6xsPQ
fpYkI4UmI0oZz0FoY9MHyqxx49xUIo5Ek3avId6fTDCsRFWHsMKSdF5Tcz6YbbKPdkbme2L9XDQX
qGyOAG+ZHyEe5j/csvS1ZlJ9n4Gs7ULftrTkaqOwkjzP0zMmeR4qGAmo1YwYQGbtBE1xg/qwpOV1
enACXDX3zZn5KR39JPydxXQC16pxrFrWM2qZUS4memjdB3j0NZYeTleIAhboJ9CQOrW6u3YHffSe
A5qb9UZLgS0VtRR4WhFYrShWAAbDwVzjv58S4Rfn1ytGPM/PuRZpkW3WGbSVpwW+gDiAkizJNrH6
okJn2tE9I7EREPIHgMS5ZZfTZOQtizDHQaJTSpew+kJf4gDOTUYMRdiue6xxi4ovNi/KNEV1icsx
+x1zKvt6V11hYDttGvtX6cDIIj99mPX6o9kqkyFJ7vV45izydL+ooW2pmLey54zasebf11Wgll9W
R1RMlwKxreJDiEUFGIzwx9WZcj9xhLKVwiNG4tiU2NG9YL/VR0ZDdqhWaW+gpHoqWzv0+rAu+sxV
axN/m3XqgZNKx198XhARbVk2h0wm4XdEE0D0aA81Ju6lVC+xNyBCCjVRNNNaAvZnlN44kY5EDNFg
ZG0qh8BhyNj90HCBxhm0CfF+bG6ClRd2vsd+S3jlqjWLjqfrMXZ8vxHUkZwPcJlwunFbgGf5qP6b
nsWR8FKanXYlkGJROEZBcQngiM5tF4A2p70ZBx903ZzvK0gnhvK4PNcJkIgaAyHQxDORSBThutns
yLWxThgVnADO0HvmjF+itbMpnOEgnWKREXY29jiN1oJvRmB/fiwA2+XLL1WH63/TGs4fd9RIgBBA
z9W10UCe3nrAMOw00s4UQVwXrfgcB2eJGfZ6Ujo/KYCq4YQaRoPnHAukE21EazN9joats5QojcB/
0u3DZest9wz9sB4TFfWrbYKOZ3N/1Uf5vDagvU9bJMfw7WLz4pi5lWVEEEsbmawBQkCyyCIPFczk
3YWdfyL5UIJRZo4a5ABPmGVx69Ml1nw4gTeUxrfSlfYYQ3hgiEqusbSz1imVS5spj+UMXhqlOi2Y
t+LCoA2EBbGweQCkDo2Avny9hEW5q9xxPGvfJMEFAA2P8IYbZoA1oVi1dOGNreepODEgJRnqPHeE
EnofxSwn2TmxV9pPvdDNcwLuNzjja3mnvAybV1TzjoS8aWMKmv1ww0aXo1VUg+mV7Lp4/YtdHEVh
J+vvJSVQHUGZvo3N4oe7s9OYO8FU75HTP7hYwE7DIwiOcuDOddewVcvHzrk01iq1jxj0+kl0hWvc
6SABXaJCT1cCu4jg+U6j1uoviW1TT0qaiIPkxWmeD5sVt7Y1HtwtZveLPVR2DMfXH9w6OYLdkCUe
T7lScDDdBgBNsGFhfkRG2GkpKOS8G1jHDcTjB9p2C3h4Exh7Xl4mLcNl5rin3cKke5m7xuTSKhUa
9I0dlrStSzHC4MITOrsDjUDag8tsCLrIuhLNux6yD8lSuw8DZPSIAZDHHFnUSEADJaNaQU5j+Brh
jyAcj1UIQjJjxFAs38xy2/6NWE/fAtxFh3c4yI+uToP2PvEuMcruPj31SGgPOqahnD7eT/R5mg5o
w17bwE66R1hulklKZGztRIe0nXO2zWiCnDEIZi/SGBZdZ/y9kdVrp2OU1N9JRRDLJ4uJOvvft+i3
HwrhDLZkv911zMnS5rKgW7KCL2oAb5BDPCcdxqJ+ELsHtTwFhGQ9rAzlbGA7f5M4FXKhUOakftnn
Xk/xCBmojKOXBHYsbpKj+ZAO9GamnqaklELOpp8qrz9e9iXauINXZ6tBjWAUjGEhaYR2TPsvyF5+
FtTsyrENtSkXFjeASgbfrq38LkgGCfi4VXLMHEJ4rA7XCXHyYBWTfW827XEKAmRQDXHGPIg6Isnv
WGof5r4R+1OgOhZVi3wLIyBjKHe6wHwlNK5Zlj/E34XUvtvDJCkozPhVpjoHLwkK5yQbI3UQHDdR
chO7J8et5H8rZ6K9JOlLIsV7zAxgYTjOH3Rn1PqZEssWMz80k35q9ryRH1hDt4cETWn7iACioD0e
j1WoW0RtBY1wkxcea2nET/57sGmMRRR5uohRu7/1FU4hDMtTChB/aUm6Uawlc5cAwCDaiDmFt/KG
WdDG/fZL231Yvoe1EtVeCRJJfB/2AquU3LhJsj306bXgQbt4rRhmRWRdaxCILntjKBwJBuViFhsi
61H+VoC0aDCCam0mHgVXZV0lOg9Agm8v0+HsHuvwZV2F00wrRZJDcHtThGDqblT2SQBThWUi2oYd
lyt7i+o1dE9u03KyD4ZJe6N9qVtNhrQVKvWtc95Rx1yVV2OT7OUpi3/Q+2JSUY+QR7+TV7KVzkcX
kmpDi5qDLXsGBptK4vDT9YwH4uJ+x2a+HXw7qDcc7Bo7VHry9b3A3PG9gIw892ZbXWtB+FWC4JRl
T/koxiHtHdYMLN59xMbXFWN7M4U/a9UYAwOIf7Mer3DZqOak1W+BEuUOm11dm3ZRzBZOiSmEluK5
d6gDSUDv816Z6Ptjptfb6V40ssy/wFHQ7NJ1tiyh5w1jV0b5WUjfG1IteT2IIdge3xZZpX9SCOFj
c0CDl6c1xZQgxkvURv/dnnJr8erYFvyRYC/ikNr/C/jaKS/Txo8QX06smeVhzal/Dl6sSzMffMxS
o4Rn2mwextJXusjap1UISztMjAnFNcl6ZxpgQWrPgQEYzDjBnnh0M50mRLwnAkxR+MBlnuLbeH8V
MxGQsNp7cow4qcQJyYlLeacA6Wia8JkRNiWQLgKxMcYC2695Hj5Di/FpqrUf252XHYOSBHQA9Vt/
2Q7K2tQE5T4OSaHvCQDt/LUrVWQ5Qz7jbOeqljMjjODg6tCUnYe5Vv6pSzGaxXoeryJbtDg+DfiD
ue52dbjpweJmURqnUkLJ6TTnQv5k31pCmFZ/eiNQXqirIJ9d1E1emASkZ2jthGPiZGG/NzNjq+8C
rHiD4i84eTVT+FbcMrs/0KM1kPz0NKPBgYxKo2+qzu65mfvJmnO7SkENT+8HlehoppadyzTJDhHY
dyQ7I0D8guesj7kpBo8qUvbSiCMpcfqjyBwjeCso/+V0hbCIIjSrRMr4ltbl8BwP3aJVbb350qu7
p47UtBTb3F+z81RPzVRMyzisY6RHJl3Vvq47E0OE5CFvwKiRTHodR7q1zl22ZePme0PG4IT4K1SS
FFPVZJ1bBKHnpvOs9tOitI504MP/PuSfkXd1vFTTQ5lBtmbeHwClSyu++V01fmB7KMnsStlLPp+F
WfLWH0mlClb//voEKnnSsmY0i0Z5u7v+nbWaU4+zMN0v6LB4m1Ri7ryt/6EswiH5Wy+lWVnlkW5p
tifCPu4AH3/8D40j1ymShvhrr8toNZ7+O3+g27i7BY7cSf4De84JWCrm2AUkQMoLRuuZq5tX03zH
c0biNHuDmokCUe+vihCUDAbYpKDN+awgaLAkVb0sBpSwKJwxFSlHD3boaVGNiLgLetwkHXBw+KAV
K96ArgjiluuTUzlB4ZxNqn/SzxFJUKGnJqlilvgTmCEyBaDTbNXyg+BTPgU+fyijvw9CGXGAlZ/V
k8bsrUCj6fAROjAHX7pkjFWgba71Z25SQ0eh0l5AQX7Wr2ypnRxVG27J9B/QMUzHyjJymg7lS+NF
Puhzbec2Q0MX4yQoq3kYssX/n2rmFsXEyAjyIjfdhe+NYHdrG6SkN61FlPdsXaUjQ8dg7uy1YWkI
YzEk2tbhMzYPtdP+l7RIYK4/Q2PCZCGpKLXRLRWjb9goifJa4n4WWLmohTkPCdBfeL8/6yoFXL0P
kvsKOqvpz220xWR6XZgvtFXHdZtejr0VOBBLPFln2ptYO3jNqw/wLuzdCCvBZZpSV3D5lNwXhkJ5
4NhfQO8Cx0i8zr7pVTigmNMCZe8KkIGUNmVSXeg9fHk0qQGCUL+9PLTc1x5/zsir8zcWD+0JZvXg
Sr7ozegynFUOq5dVPdGq4Mr4vbHJILM/cFtqZmP8WA2wE8gXHGBbx4CuM+i/O4kHIrpZUyKzKzjP
bJloqj6m4g9m3Su6cgCUOWDaREk+Hoj3OLNJ7Ujw0HJJFLkHfDnRMGCyISaTezQ6AywyXaHTsQza
QvGrpY+PTJD7bGclPUoxY9EIBOfImlGYVlbzjL9TQg9q5qF2GiTQS7tuZx7XXF7HAXXHvwCYFiAh
tBG4CdUtiXuVRNL92cq9RcBA6ZP7hEc08Z2wDUpDKum/j+veueP6vEZ1UQnWM7UFN3Q1OAKsiGmx
SQVuhRYwaPfcwdfuGW/9WoRiFC07u4Npzpi4rdT+qkKiP5B2ObWj6ubRD1Z9AypLkg5Y0RHDjasQ
qK6GoK/kbrFrOst5CrGnK6A3xJA2Kb/IGb/5yczCmTNlJidetvvc+IqRlUFbFqX1nCXc7WdU0hUc
DvbU+aSkuJp3CTiBJmuSyX4jh3nsf/rnZHU3KXhkzLlwC9qdsBvBA6FvtYrvyhAD9Dzx69Gcrw/V
Qlbhx//yub3zSM7oW+f/P1X82Hr4HPeCCmxbE2juMkXVxsxgIcRIPc0iax9Y7eFe+27RtpSe6MnQ
sU5SIbrG1xO9xFnG5GfxZ4pokUAIpwBFonWFUGWnrEc8AVvQ83MM23Z3FN/IrkIni+qQ2Dg3cI6y
7e+45VCVvJpvzu3woZimh6Du4po1IuZuulP4+ufNjDnGgqvP4p2IuOxJFF75/0AYafL0aKYqC5Fd
jbwY+t/aIFZfIJPmhfHhEzNkIxR0QKGpdeEXxAgi1HTzk3Ij0meppXirVTBwu3Tbp8zsUYb2ZmQi
L0EZwtpw6as5ScedZhpQEbuPPO9rLbOThAxb1aXAVunmBf61njkttynaf3sblwb8n52xHsQumM+B
gaYhHKJCF11GV04T7gA6Axqh4Yrj7Q0VcyyFHPyCtIS/LrhWSVgsd7SFXkDzy3ghAEGNUgRzG1q9
F1bdS60wtvZKzo5Qh86V5BveoOoUucSNO87rsoqmDC1bV+LEga/0I95ndSgTtueeQQeAWVFuwPqn
i1gtLTmFEk96f7Ig1FWKpLBLq4FiisFFKkzJTY4kP3UKXmGNpZ15NeOGc8/iyrNIyJbYGXpvJHUa
KHGWO8xgADzAp+IhAbgmFlQ6nXR+l4XkKTW619ti/2qGF27yM/p6WcJ3gAU+16GgNLk/BhsIMUZ9
SkLdcV5UbG2UuYZoyFIejb87wvxg1c8RhzvliIv+J4m8KIeI+JB7FB2+LU//nLGr5sJxVIqaf/xZ
pNc1Tjw8TZr2c94d40WVQvi5st6/HPduXRyebYb2ygCvgue/xxotCR0A7DJeEmGyRKQO3f8iHxal
4/Yh+K3sW2i2HfXl264Jypzst56R5u8aaPosG9+HOENxYXqug2FmJhQxKtgPCyMw4+PWZMEUlhGt
n+uwRzX+w5m+Tw8Io4tFURiwzyDFYDy6DBFedCeas+F/AfEY/IhT4UNPx1V1GtT7vo67Gai1n/cE
5fa5OJ1A4PSbDx1O0MqdEdNDy7V3U2z0pO0ia73WUSb3naBWXnszXxUF94EiZLmwQ4VKA1Pu80u+
MKRP7HH40Brtx8Hen9I8OfG7tu2U31WNZWb8dvTDNntnURlKQCO1RR4o5mSMU6eAq/HbntWWafcO
ct2S9lZvelmGd1+QT3PUWOf3GIW1Aj1tR/LrP+NZNmKxQwEKYSqN1lhjy3UxkRAit6iOIzkk9t5j
jt9e7cizZBD4Z/zaE41esPHUqLYvm/UZQWnvtgZr7rQA/OltUavI80FOSs+YqVYsJqmxVVhTBsgA
oC178O6Fx9WZ4K6tcGGMVpfa0b+N9QPBGuIrZzpNPW52kdeSLcz6qSpknj2URxDYd3noKIXQ0cRP
I6es0/suMX22DNPIfBkXRZTyOL7OAeCvIeK/BU4BXenfsHGErxQv4ldJOP6nwIHvZePGar2dUCto
w82gJRGnhsQKiYii/OyqrepyMXqoUNXBV5lw3bOenppGS3lOuuvJABx7Ws8rF1BAWYgYf0Oo26vs
iAuNPO+06Fxqp/kjr8UmZTLs2RXif6q6ovC7JMEDz1k3ukYwyextAhKUbFDilSwGZFLjhTAXl1aZ
wmWmhuulaFVlzTUaOOyEZXDXWmNq9CY9UAzMvCDAa3NwGpTiYCJ2xlhcehSYDlZbpamSgwaA2Y8G
TZKf3WcbM0d7SOJ1fbonO9LAAhfVVfXoadFic9FWlxKdzoLDKbi0dmV9r0e78hGMZ0nxV08zsoUi
xXMuCGrjqzQohsYj25CzHJCask0Bzzx5ieEETxnJ9VbnI0sUQz390rTzxhIe3qcv/PYLKRXF7RyH
Gzo4jsLrlXqzjTiNTI4ghIzgMOo9aSXMXC/IDOgA66nPMI8V/rGF5Hwul1kQSWYf70B6kTjkglJG
laJMlqUEXRBJm1y3W+PINuNWh9QphBUFgC21L+rsyL0JUBq6FADi000L8uMLfQ8ADWzPf070sjmI
cPmvRRBdq3B4XT3ZeUBcrBQR5IqvK0Cm8ZNmTe9+DEW/YwtZW8DMPo1Lte3P0nmj61Rva6eY1OBE
R3S3ln2yKwD9qPEOvzZZ6oWqVWVwVpub+J5dsSYaOzrO8r8EaEgXz5XA/pzZMDFm2Tefn236G4yr
MwXWmn0eTdek8PV/EU8hUEkmdJE0zOhph8kgfk/OcikyR2B9S5VzQFpAhfmxWPnJUdUW442Wipq+
trhIXUdzmhNozRngMOWJkLsTXfHx5khg8UFQVgRgLf8mVw4Ct/RsMyXByp8EEf8NXsoK9+GqxP0t
k1/ufB7HLC/qp2peI68x1V0xO+djkNVW+hPrL4jVUB4RIChYVD1ngNasIOi+yEyAPg3A3oMsuVJV
UHqQ7jFEI0LvcMRtheRuouODR6ETlcK9QIJ6r5ojNu9LLc9XC9Nti+CzSKDBslgiS0MaXRMZMehg
zLtj4Mf7zadRm8WkDS+SOfxbzHicwg0jKQZuwjphAuUkTOX6gJmGxCTi1tkFCJTc4J59fUNDbE4y
hHLi06EQ3OJ9R6x2MXMf3xO2jDMueusAJLp7pRdvSTRXcA3Pmyjue8y3/aYFMhnImrTuEm9YxgZ9
J0l7ObwcW5jlGCcBJiYf5mltd9HPMp1fypsMR/8pEJ548JEvD+01poqBoqLYyStMgJj5YKD16ai5
SqZ+U/ua8XSkIfY3OhlQgHEHQnHp72pA5c5c1keHJbc0mpMlGy/FY1DEXWqQ9bso3P8AYdkgRimg
FMICKCZRbBGrWBoo1uYndb9mC6YQATH++wgO0l9fW++20PDD9RVQ/7JzTCOTUp4CJm4mLEj924Pp
bbtdngIr3JSuherF3Aq2ghDEwxnFOmfjSIkAElfz7WJoTUTs69t+6VeXzOoJFE2AqnDo/iQs/1wC
aAHIn9kWMIXMqzkAO1WegA2INx6Boj5SSgjxIeEBKfSllOmfGon78cq0lpm42zkDH9imRppdED6x
sEuShDW/EIB+GJgUifbop7O7Nii1KLe0VvYEO3owH+0ynn+zWku47rkgIRYR7WoEM9Hek1GMAwaQ
kTjUUqVnffvKK4hDpoj8nUlGEQlK2ZYS8X7SKjxTsKlZTQIyNShP9FEND4jaTlTflM54SNNieH1v
6bGhxZxi9IsIrZooTpoirXPY4x5rJm7stHzxuE/QFrcdO9eMyMWqYJtsxaukPqe5BDg6SuczRTYz
Wm52rHmTsC6q7FbS7gbdtmFPkp4mYjXE2L6okGy2/JvYitZAceK6F2C8SY/M5tPF3k/x6ICd0v+c
CJkKU6mLYPuRBNOGaPAEr0PMp/morCUM7aV1WyV4Hvzg6loA0Xx5Gau7Y+9AOZ5yQFBBd3zxG4qt
GKf4FRxtkF/jcrVUUamEf7YlcbFJ3DpKY0wGFEp61NQo3+B5DDFZGOa7rU4Z/xBtFcZ0dsHTjmBd
0YNGU1jLNQp2PvSX4g8ec30K4NpbX84t71HfAw5WFvfJiO3xFBDEBzacpnfFXC8ObUZyZgsPK3QH
tkGDlnQqY+ztpn4EAKmKXwXKQwRT75Ti9S37Bx68Hi9cv3hyADZNIxStiAcG1G0hzkn8BZZ0Pbhe
piWYVYxBY9vBDQTgDX3vMpWBaBtck9x6SQtwhc56EyZPfImjfUzbH3UzNo8xWD4GBqx2WiK7vNEd
YEzs49r2S9l5HDw7NVu++jBEnMGpCHnpxx27T7ayo15VWd+/3veb6dq7ZR0NwY9s7WMIaE0abSku
Ryqeym1sNHq1ado3fP3fw8MrFQy0BVrDQWCgTVJsYeI+CRWTeOcIW5uD5FXdvA3N0eBAEW4Uh99e
VnrbFK1lKTtzJop7hyTC6E1Ba9JDrRCjE7r42YTBtUly0PyfjIh8tY8G8sy2B4aDdEBfXwtVl+bC
pS25Tbd+VOp8eAx2P8IKKJ6VpUIMZ2IT447F3mFOPHdYooqCOM0YSS6BSBUnAoDvFMAaR1C5qRAW
JH2ltTeOvCLjjY61ThO1GSJ3koaRIQA3OEadLdB62SxHz7TMTiuRwOop4mLNSDvzY2JRrIoiDSJF
dOfpjrBMQjgvNipI5B9/K2JT2O4em3GoftemyHWftWNbcV29062e2DFcRo2oAsqYBe4QWjm5Ktub
XoVc/E+YexJvUcNdAM0WcRiBY2gEFw/ur0dcjlgRV679g39opKRwkrcxB11b7fUWVrgZ3Vkr3+W6
YKZU8KjzUvil39O3wlMX4+dA5B8rbbX9l8E6f1SZIggBRAKiRlYMO4PxDmxSBsW2caFZ9jjISGEp
dZfRChoUBkmuspH70SNJu5BewMXIXVwkgFthd3RKesU+NQeSGVx78B0Q7a/54AHTu7I8odiwMy7e
S+wFnS9z9obwGO4yQkid8T0Zzbx6YcSMzx2mhG9RcQrYX44WXyoeJJ06XrNs+YXJSTsrkCEc0dFU
Ni6e18B6/eweuEOmK1K+G/Zf/O7VfzQwes9rTEx8pnKKZzGZip0UYs4A+SoiJx0GmGZVK+dPJBuf
fwTp4uQ3AUAFy2CvLJXKcQ3IdfGBlNuNPALoByve1DfZEnXgGnOU8XejodBAVkKgAPpNkYiN2rQ+
l9OsSQVgyXtuZ+gc9nCx/d0hHqiWbAcK+I7I1nM3L2reOlwT7sRkveDBTTre89fpIR1kYHAVyYAn
jElK9g7ew5Zd2DZiak7ncpuzriVg8PUuHS2kd19fYy1gPRMiWHRNt2yG0CQGZqal146yac1HdJuo
H9u3oRXBtgW5yer0+9IQIx4tKsdJKeFi46K9cdMWm0qjgiqK5Y2pVm2kfpTmkNhwK0hLim/Az3T9
MVUISMD5LXhK906Fdm6waDyEs5JlQ3Ihp5/yfB1yn3NFo8fgtwb2p0af3fgNFEN+V9qdGfllAT3W
v/bXCVu21VydjF24sOVZMK1Bef6tPFt6SqF/WT17/mlLGcN5PnQgHzAOQ5qpqI/nvGb5Sf0zT35D
W6cY2Ic/ordF+gAB3j0bOZRbOxAXFDlSXTV7DgPL8PMNVRqMqW+yh6/OpIhpjhmOuVta3tLFscvS
8yRA11B8baQunTuDXNBWLsBxLceFqft9Y9X7cXfEsbeolRcm+BBjGRngc6sqKrVXIcyENzV4fq4n
GOLATL+HGkOsVuqi/eiqHJo+yFMUzQ/EF+VcH94dKsWf59gg1ea4Ta4HZHYhC5sK/yTGD5DDZWsn
DJCpwSl1ZTVEAoyDKO8ghRpBWVfaYBy0eX8B3SwAcNkPuGW+ygo2hHs2ObY1yAy68sMlYYsTXjNt
VQm6ZgmbC1g9b6ar+nPMRefyxtIHWD4O/cLhI5Suex8WwzijFDV86Z8wdRPeBxDeEQcLr6N0u/6n
P7mFpngigWldLTH/FOWQa/27Rj9W87s/lQdY1i2T9WUNl4gzP6GUX/+QlGtvCt94fjDjVjzTNTSG
kg61LK9jJ2Ma0v9c34XRZRgoklgBVXsVkmOE8xdd2YTT9OiiOUYgmomtBrPDT7o5frRazj4df0Qp
byXvdCYUphgLIi3KNKjEs/2gCnaL21tllfSdx20IaWi0PylOsPSwCmNhe/cvefcrq8bceV6LdMjL
t+cV4oNoG5aMv8DAGvgZLVZBwQHnNynJnT+5HnPOhLTrBYZzDx9j9u5Zey/UuHk47C092UE/YMOu
pULWhvzyXObhDz7VfxnOI1C4mPX8zfOKttpW1IU6fwZHT1cGDNFZt/Fd+Vyn1bGgjyz7T6e4l1pu
hKiX4Ba9h6vG8WhaeyoqbsyRnYDWtAwgFgCG1M2SYCWciSMP1el2O444C1SAsFGTyIu9k7OWOGJ7
fzXNapd/gwTnGvapvtQ7mYP4YpjGe6pl6pM+Kap3wHodCG27s2EJVbzunPKuk5+5phlfLUj0lIGO
WRuP7W4q9Bj2jN7YpUbUnEst4t2OaT8qwfzhUlgraPPscMVvsHTVRhr1aTg92eHajPYT2hziTr0X
cCpTZ4gOlZWa+glGJV5konvwgelL+Cxul9VBTbw2Qm1rZ6OW0QCnjkiWaSF9M+sKsQ76vPuM4My9
fWI5TGl3ejBkvZ04ofILr8qwL4apev4C1bJLQ1DrPpi5UhHIiSmBRqMPZfYwXwKc9JF06VVfPSj5
OPw3Lw4s/unG8mhxCkET/Z5MhQXE33ZsW+D50OfSDM7Rc1x9AOOnfmT6CwEX39uBPCQiCcSv6GjO
jlETMczhlH+CK7iAfxfcaXo25h3nPhJuVIrsRrtnatLXQR0YTMUGLczLN1ITrxJ/VQrPF4wHhJvw
McrTZClL6mhaNbtFCO3fPZFtbI9+N0H2A9mOina3TrhH3cIxEZF2tN1ii9NLrfd3dB+5eIfsqOh3
UgIAqBT2TNgOCbFck5Am3XCVYjubjL7V0rCtcAvt4OhR4Rl79QTWU/KMktGZAOu2ApuLcrEGo7tp
II52GPddJs6rHaqHYccIxJyvsrtfxl63gRxX5tdW3KL/g1ewzMcI6cYWVMp9/gfN5+KYnFVrOnh/
Vcjg6MsVmxjeMPbn64bWHMlr1qd2Yimw04JfLTyh1YKRFLV4YdKnuCTaDTvxi7NvYRzptDW2syhl
LbqCtE9L3Qeq6nLyfCCGDBU5jfHWcC8e62w4ZjzoYunP6z9mEOhYTN3E2xTBoi9KztZHuqTe4Vv/
6Os2K+603ya28woq5nbFQV+7ggPJJQ9x6K91Xj/pFXQR31fYXvfjH3+4Bz5g2cvw2Lvxe3S9F4PM
pvtcetO+xv7TzOiXzAEjmcgkTh7pZo6hsmxYcXyl3x1240FxgKUVr5SIjn+/BHTR6FjbJN+G6Pc/
lWqb37MPD04imQqMzdTohtBM0+CDaUp4ckOYp3Zp0xQJahVMPyA3+BNFTNYim83AswwFNktfasi8
nZD5ouCmyO4tpzOERJ3KxromyZ9ROfKmiPN64eyktDbfmEgoXYbQ9mXz03Qf9VaZ5neQmLfmBXLW
ehwgZHZlfY6pY6N6wXa4XEx6t/bl81A9fclZhMVegldsWlyazzaiIhYBLg5pcLD811jOtx5SNh/2
s72BDbpygsjzoghJ7KN/J+S/ncC5alMHMqrYbFQe5Q8tqYDi5oMjWj7bqCzzGdIiHCWZfMeUEQJ4
OjT2DxDO9BW41VN1y3stGvcBjBkq38Yb23vznBf/DuSFLyR+5VhWyHfqxoc3amE5/5O0TSbHcFLw
+FSXHxeHlvKAQ2L52e2mUBC1Pk/ggvTgF2594gqrh8f6HbJEURhvrD1sm4RhSb4j4hLJDFi75SzK
YUqXo/uBw54zRh0QfnuAZcga6Iz3N7Oj2tGb1HVzo9iwB1W3/wo1NI6/1rn5QLXVydSx6o6nYtz9
X3NW6c1AQj4EvJyXMs83vImipTxuosB+LJ+zPb0OXZABoWMpgcI+U/H1W6ghM41jYVi14C+koDPJ
gLLZfS4Mq3/JlqosIVw7ARhNr7QraPSakVnWOE958AEyHh2BxALIGrqYNlwjqXEiFSWuY12KPJmQ
QdtV6+wPbJb5ZAhCtJj80mjL373FLN8EjpjJE0fkwpPe7e3bRqUQz8C+nV/994lzFc9qeJCOfAOi
U/sZGa7A1CLePdRAxIZ+s+F3WOUB3siJ2Z3iu71mnedqIq3gy5b2hidm7rctWccxY7lbWqxE9xJi
5WWSnKi3u1y3K7xHssJdTMbUBbIcyqOIoo8xbRw6AuwBreMijwdmy19/DbIWb0PNnjA8S0sDcppN
Jfb3QbVpu1MXGgTQPf2sEYWFhr86k2z+91oqkw18DOVHl6Ls4LkKdiGtSF6EvwHES9e01/Px/5vh
LxJ7A2Xyph0X4fi2tXJZSQpFpzhw/ifqkvMXq2Uv2SRjoZT5kJbKrHDS8YQTOZiUQyj41EgWdhBr
bRodd5CtlE5rFzmOstFM2+ZR1sCf6N+Jzjmn/99x/Qd/mJGR8xehIKKCrBW2ul1kmADmkRm8gG0K
ibgR/EGYuwlVpxfRRThvKMib9nwCfNu0QPEPQd+NrtZw0i/kt/kf+giogi3KfuGgKJ6YIDS13Fl+
kDHfnj9LPkJunMZf2FvndLxBFyW3/h5iRjc0A8HytnwvcKD4AYHfBwyiqVkOOUPIaGFrn3nc+kvr
t19rViEQFGKgBbcA1T0a9Pm7O3fhfctQ9YvHTrwGsZJ0n2gsq1jTW+ylfj4u+LZ7SO1PxvNV3Jaw
2eIFBG5hJMK3mBPgVRIC4QJxYDm6I8QH6kpFNU/mn6JymaJUXyEAWv3axPXmZW2trrS98YiPVmpy
pyoeIffRK/ifN7Vpywh78sgtNcI/3Q2gYZF0TjGKHLyyECcsjh4fG9pCK3c7EeAU4oLK2NJTIfGA
BxH01E8OIb1jlrc+G0lDFEBNUis+GOGycqxln+hvB8dV3Rp1yKP5A/Tp8rQdtZbZfLOMl4QvkCh2
iAl+5ds9tcHkw7br15PBko8Q4Rp8k6iohblMPU5rOZcGU/EWFdzKGdLm0yz2uYQyEkoMnxKShqio
kKHZOOxDA2GycVWRL93l/GLfSOw1tEKKrhuNuGdu4J1A8Of8tZX9nocOYRdhp4CTedQUl2MjVTBG
h8rInoUyW5ZGDRAv30FmXTg+fB1tlKfg350I0/6AUbpMQ5Iq8Y8BSN5zVfIxZqcN4M6tGbl5ZWKm
jhB0hGi29iHNwy2gg0DFkrWLkyowalSJMCXRDIqYM4SXwmZk0rLQuYwZR9lxDLIcJEE5QqhKJfpY
6oOJzPG39otKW1eEZijVPrUws2vNKLi0DGV1ge1CEhdvkIZNxgAoCb/pcrBqEDOO4j8sht6uaf2e
2vd4k4X1UMJOHloG7ht/slY5+I5BCJ1+kmGuvmtmLndjP/lfbxNhDGUNqr03Ktc/YqyObv+foFWz
BZQ3U8J4Rhdf/AKYEgfzoq4HDoVxGxVGTucSUUcuquCbYOAijwShAdMsdd/J9/HAjxtLTg+lCBDQ
Q3pdSc09ATHxJyeVekw2w0vd6k/pg/+bepKzSGp+iPjR/494ewZ/Ix9Duy130UY3pFXa3KJ+lAS7
6CxR/YgzGj4dYTNnZoBU0vyNFAhDw2H1wtcj9bAxWUFPUQAN/cvDmS4newnUxsQ25xhqRzOhJQjW
oF7Xs1dIwneDon8m0UpoiCyXy5evB7nJMKShZKfvrNM+3E2mAud0BKa+r+89Q1qzEJhAKK4ye0h1
g8ZzwYeP77b5rGzfF0klZajgoY70iTScd4eF346UZKk4a1psyxNvAO917Ccxr9BZtc9QdrngxxoZ
h2QxkorA8HdkgKdmV2lKUbUU+McC5XhDAeHioXEi4thREOvpf2E538hLpYu5egHyN1ShyVNAYKBC
vOt5mQIXIr6JpuibAfPQ9dYbtzr0HzYyKuLPfrYGW7fbAz+qemM9eKCjSpmZwh2ZzybEDh4vzB3u
/fnzDuETGJ1QvbchM2N8MvGnztPkLcVW4fGA/k6pEJY7++tNOezl3OT2jxjqfEs9HQY6nK8Bo6qT
wESHXntYh5lqiIVaUhBnBe77EtcvRE/v6xJADP3wi65DDej2tPtCsIvmB+RrP7SvwXPHFc5u8Rwf
bzJOZjY6OJbY5P5VltWNZtMN6+t4H7BFNZthyk05X2+ahZUrqI36a5HiB7tx+DalV02OB63XxGOV
g8PnjwXAm0B0lNJVlIpPv7YvD/JbS5iv3SITR2MVTlr2aPdGIX7jHPYwGrbpQ/HFTR0sBHTERpEv
Mj2pBMky3RegFG9rzDjnd+LueSvYHoldmt6MrThOGQFgrI4iXBh4XChG+YyFLXBR0/bDAOn0DU3a
0aHJxDuxdhDrbirv3sL6WO3cHcwV+oFimandaLkvypSihdED/fpwsqNmNn1DgcqHspkhnXmiScUl
m5wbYmnanJGn6w2rKhQrJbQciJp2f3Qz69vo+D0Eh69snbQFTVLW79iZ8mykR3rN0YWp3OoGnPbH
wnb5AGiu3xtXlXPiZB0+6rUnEtrWN3oWTDXCckYw5xfUfCOl4O4P62OG0GPpA2p9aRFDxo5guVxZ
1LvdcQwmnr2zl3TQz2x7DgS4rqMDiMenzuO/tr9RiG8lBO99tusDxQpiEL0ogsUdD4s+F49xF8Ub
l+Ex6tkAV9/wtGUSh1i4B3KYl9UVKCkwE1qMdcm4apcyD9swEnl5R1zp7W7qvWjS8tUvdgn4BeJd
Cxwit+7MG41/ZfwpoJ0E+YRUZiy1Bn2xp6bO4wZPOGfcHkovbVakcjY6CmN/B8sqs6enJM3SnmmN
KGAh8b58qLzQ/idHK8LIwLgd34udn4Q3APMbKWVG5gHwj1BPee7zmYc7b7Go5//MSJJM+hcGZsqV
ojqVH9VZkqDo5RiR9u1++vz5Z56RqVeWg8jY/GuwaVU/IZ+b99n2dpuhIlbv8LzPb6jcCSScoxoP
rvBT528dEE6Bvy+N/5Ve9x7HLm+7Dzj6Ars44qK5p6ks4U1+sXtq1fHTCITPnexWutlZS4z/zKj5
f46VbGpH8yFTHAhJH5fKgduNTnzOrOfnUAu/T+RQzVk7yCC3cggJXYpckFSq6ZQG6yQb67eCRTtK
FGmApDLDSF+hrKPO5nz63g6U9A4sjOEJG3KNy00HmWa8C8qSoHQ9Zcor9Gs5j6BeB4ppSQ17j5FC
a2lhp6k0uezDim8hQKChro1+MMSYANICMbnQAT7ZVfP4UUAMSvrgcxYPZvAtAFf4JjwB+6fU7oSa
nfy8oYLoAilfUXIb20+rNoYduGqCUoEu6X2IagvI9l1ZHBJOkALxhzI9W8Wk7BAxcD+oUcWNp0uQ
dZ9TRIMzayp0IXuMzPRHt/KrjEOgGG/0JGPAoVT34/7nKEHuAHuIkgLY/V4Wp4fKM03PGj7c/EN7
8EGfSfjUSyVaIObKrFXW19M6ZYAnkHFy8Y1p23Osy6vCjJGP3RhNSts85yY9kysX5apdUBavhmJm
Ycrx92qjSGWj5uPMa5qswvcBpbNQ8ULzpV7x0OqHvyrmkZoW9k1o9muzn1/oIAR5+jGuSDcNulyV
RCrZzgS6a4+YGFWJgOU4sF9oCPcWCPdatHDFlwr2A7hQ8BDWXNYwOrtKnRR8VIoScV8Cw/BUy4cM
aWgEaJXkoH1bo2NBOjPMhOzNJMwtKtVIZN3Fo6PK4w69D8p3MBNxzIDhj+6JdP4R0c/4bsflpsjE
AFF9DxxW6yGs9qnSaF2j5HI8KWWqb73Cg2MCVctA3S940QA2S3oKgS4KZCkOOiEW/KUrlcN26tSH
i4yOth4VSPeHDVo9yZ7l2NVp8x6mUAj3zFiHE01xJYnEmhGrUj/YwYxl45/0n1YDzWEongNIg/k1
NEjh/34DaTuxiW+M2h16AosLa6U+X5+JQS0rtR88HWzSG3RJZO8WcqYErQYT1GVzMnL+QQ8oLarT
al0YtH/Ll5Ksgvk02WQLXX8+HcySgzeB8opHtu0Hg03VRaY0mZ+yRereJGtpvZ3hjRXz4rShj16H
rpyAmd8w6Z8UQhdkNe0gjztvWMMQQPJ94XMMd7WAvo1c7wFyhBBzoNnIu7iaQpcIWdlcymrMaaAn
i3Yy7pIUJGIiWGMIux/7z4sGN0Ue5lul30m/gv13R5kNSMbmWyVwKjt9uDQRHkX42eJ4ft/O30Mo
aojWE+FJ9J5iIKfb3glrqCPPncUJMnJf4MRsoGfncGtll5atBQdGKbOADU4quIW4tpBXL3SxGGQA
auDbjUfZo1WrsgIG2IUv+Sm7MwcXcz1v85b728JX4VoHOAGIdfXBdoVds1xq/1WCpuDwf6q5ngYv
Tm1JVjYpDEcIXgm9DS8Z40w5RYlvO+XEJ/EZNCqXPRJTqRMkYHaShICWWFyrgkMMub3NQu9ngyoO
rX/KZkkBN8GBsClXQTapTqYc9IBf75MXKNyhlp1nIsPoDn2vvFnMOE4yB7/TKh+5u/0KQjEkGMHm
fCE6P8crsoGvUXCUsjltD9jGDQ3WdawRdUYDWm/Ie9bNzXitcpFSq19Zur24puhKtpHMwI34JEcK
j4LARpocdDjVHhVTFbBPkkVm/NffWVq49NsL9n9JvrUeqGmE3SJLKD3mVXj2ynd9nChxcXh48bkz
qyZJ25Kn//hLlA+e/NJJ9ngRogL5tbpICiQ3UPYbChQcOjGVvU0KHLPwoDaXLLD+ZqAhkvmUu1Hq
JG+INCq/whvWU9cJ0j+Br78d99oXFgIAu5eZx2IVfFiABWryNvMKIfb1jwVR6DT3YofKVQshykgQ
voa5R+5HJWWKM7w3/RUtJz3OKDSBMXRbefAdrUtFsZLN5eTynJLkchdj6tf6qn9/UpTj4D5N7WuZ
JmGLtHaNY9UJusTpMbVWHgat5tZqOreeXOTXTHAjrLHzZYXfYzrh1pbfYhX/re810eteUdzqmwIO
eUs7A6WzK4xgtxDHE/ktfn/X3Oup0Q5pkPsQs550IITU9aEwKxk+99c2aeZJA2n7oW6r8gelbnKS
jGlcP4NeqNGcHZTG861YtCnWMSkB7aJM3BzVQ4/fKH6C0xDKLJwtyhe4cXy/YVbbKS47hARiwnPJ
ybFOmfVr4QPCFrI+sgTZYLsv7ZrqSS0XR4k6KWNqSMu3SVJyTp/g5KBtLn7xLanIBxKF4vKX5d5H
zDkKIkFqlu5oM01Vrj3LblCK4/bFhgqOtJyF1wjc96PzsezzXQpw1+txNg+vZCHsD0RARIDoL4Vp
DKt8IoRsTSImQUbfsrSn4+Ec7U7l7TW4/adBMMWJDDPlb6QjjtgXygKZe9R55eM3HUmjikd5dHjt
wVtFjYtkS/xLRaip8w65gjwJqvLLW0o9L3H/RnReIZx2u7DC64FNCLGLSWiXbU3EoNBcWkWn56G3
Rtkr+NUeT+FNchiCYJvOu1O56bGwxHRpydx22Xi8ictEosV+4VN/xCeNgWkns5zbKjYys+rKiton
ZFhi4ZRCEMppz1lLPe5QGSNChSkedu6ujq6TAyUi25jzvPkvVm3Gx/OMYyMlZ0eAQi7IOsMqJwl4
Uh9jNPqYWj9oI9fBptC/DXmTWVq7VxplFKikRj9WhGMU5MYVojteq1oZzHQFRjsAdNGlDCB6iCXa
s/BM3tRDE2zP5HpUXe4p8AMA4ODRpupILzeLHajF65j73IlU7FO8G8Dt6PBMOn3WzQMvy3mey3/+
Aw5acAIpCE4/EjFDaiF2/cKqovoOakbe/q1C/i/qwzWlJcBSHTkVEd4WGqBgH3MHqved0WuRMz4z
na0yvffl77qU16BLGAirFpE+avAiMJGlRA8+SyQdN54LmPCfR4XVmYb8KcSx0QZCv6d3yL/zziyp
m+myBtFwgcaABQ42H23o2lfmes6iCJKEcJf4F81KCqbwRN5ggCrT3wInpa8GSGZ7/wGVlvG2zwn0
QUms+zVWhjfGAo/I2ogKDEVFbv+tHjNYEoWNgmX31KNp3wuvWEEjsiwBJ/25CWFSF2STA7XySKtH
SdeCTFctUopKWW1ij5/H3PU2SGPPp75vHmz4jXujm9thHoLqn4r9CBns7Aa5obEmryN5UsILneiB
Du+EZ6LkGd3+mXsKopu1CYcH2bpMmum9yztkaMDUqVZ/wHTOZy/LN18fkTDZpGU7zKAdWRfSXHis
U+Y8EeRDY2mryB7ZhLImkTAJcPWYL4i/sOT6RDBtWfSM44tYZmO8fp/mr3dYs8zkpKw3MI8OPsU7
GNVD5Ds/wIG1AC26ARBqHm71x7ubpORnTv+FN9R8AGvDCAmzv7BQSTw3JjoqxPMYbxRqsj7sfepC
8nILKCnwRzvaZwQSTBIYWo0LT1Jcu2zHgYbv9mmtMOI69O2qwcPrSnuXzKgbwvXijY5SHCBHMKne
Axma1Grnb+jU40n0BIXJCFzIiknConkGvb0N63tYPbpPL8Z6M67grNrYU7lunF5UYFwhiH2cUd5/
n4IhPbt/hVSZQM4s0m7PlxrrcTdE62G6Kk2BXXPjg4ZYqizbYmcNhSNrLqLU5EX5Ow7zypmah+7+
ve3byxnTXSqTPE1mrDSPiIPZ6PpANLi39pP+6CkS9EmkXP07zBAergUdXJiPnhj4glvltKUu0hGm
fbPmB5mVvmIG07vns8dcK+TgLSosu3t33lF58p0VvNVgRhttPKsY0Uw76bo9Zd5Nwry1P8Vq7CUE
Zxs/Tp8+mxDVPIj0P7Z3hFJdg6gvNLfPAxaO4S4VStwp5tp1kAdv/svqa4D2mvzDjIFWn6BWl5q6
x34KnH6Ya65bcBRmf4/TMxv202JrF3Gjti26l/f3goR1ddol1a3zuiIVoIhdGahddFWmRQT/1q5l
I/LgLRY52chGTio4LYbOQE+Av8bDsX3/wJAxDHhhhnN4mJ8lgK7C/XwTz8NneVmqCiPCCqkBZP74
XDBgWestKlIKkNwhHClss/7/908d4RrVubqaX8SEvV0Knz2Gyr5hiHIMT+v0nB9HvbN/o09TH0+u
cDGslPdG2f0a/+C6uwDI9Q0SMxwdq+2pVfw8ivIGuqLIxWhnz1lJiCne8lM0yQpT0f975WsSm2RZ
yk3fnNXoF6NwMLZoZOZML3uoAtqVeSGoItTBx4zwOuvMJmRKmCXtAC5DnK9ENXxW5iAgjc8vXG6p
Gh5tr6E/o2ODNmxfkE0Rf/Q/+7vevFEAdU6GAxBTPMjjxZvATAdZpQjprxyCzjxwOA9Np56UeQpC
FgYrDxi1qvFS61Ki4C92jmeZs7wbSuhFGcMmiLC+sv/lOs9vP957AT/LFHg386Nz2z8HJ0bwb/vR
XOxZzF3kDKVTA7j2i0dECYx3ek6y+DEt5XNmwpH4i8AMbTIHaq4GVUlZ+c98QW0qQmW6FqtrKgG5
2h2o2xTlyw51gSNGYrzr38NMLdPgs5iBSb531rqViNRkbPhzW7rWaUtW3PeVSbR4n8JYIgHEnnvi
hMaIXAeA/dB5HRlGNltHiUosuyLQ2ua1bkAGztzvDI003SChAyZckvvSuea9uiIEg135mDzJ2B2N
5trF4Ck1vwtYR+4+DY33TnN3IOTf98LgizKnNJ0K1Y93qW0KaWk5WeuZey1/sXKQEuE1GZz0W30H
Lm08lz9xamnjUdRoGxC074yDKHWFd0Z62R07fO53bONfb0ERZyeHq8usKhGpBO8ZdgUgnvyAOjsH
j7xxtKPWl9stYwueRDvp3CEb2ju0LagiWuNWU1WNXBte658gqVyax8ChGn3dSfOkFT6lTiFfufq0
ZFSngR6omULYTPNCYCqoLSUMvcZwIlmOH0hO9sh0QfAYQy9lq1U1wp9/xIG9cDLYQqudTveSv8u5
TZr2UUqiBTc3DAM0O1W1yp1JNLSYpEpqCwrE96a1KOVF0EFn1hkXijf1FY6jDzgKICP83K8af75r
en/FmFX969DIFADABClonl+AbaT/EQLCh+RLdaU84j1MekZxsCsdOQ2nTQkgQnNhbEg3B7K252T1
P02mCe9CICBsjlbmrSbYV+iPuOG83uA6QCEfICOiLLEeMtaYSe/TmXdiYXYkEjVd3Sd5+OT7mNmx
sDDeuG9DEm9mMXHRYEfXM1UBq2R/F52czsmPq5UHJ/TY8gVC40J0D9b2kqWXDWyBFmNNeqbkpJJJ
Nxys0V943t/xok6vK5Iq4xJZ26wcq++5jmzIQFDNiVwdmlyuYUbNEc9AHrgS88AzXCbnA5TlYnip
GokhW5pvXQ4fu4H4FX9bk9s9emEWJ1Z3FFF805/K+dSLJyBlLCfJxOy2Nj3daMpaPSe98iRnz3FR
mDwxKEhDeE+N+dIpdCsLWtKY8RM7Ra0LvZKwc7OpZUjxYvKC1FbhFrruH2r/AbKE602qT7CMC/P9
w1aeVGR5v/dm2PzC72t3ZjcwXvJVEAu+70UEEuD/CLOoYIyx3xMfSb9+yTS8trz24vv2PLReUbhW
ZHdEYubyD0+JQ56QW+6wxqk9EsyEVhkSRgitiqQ9z4RiUXXvXdbiXrpE0fxw6L6D6XjqtANZAhaH
jIEz3+tCrUoTTmK2GOaxu/qEB+DJfjqePnAgW3/XgaW2OqG8oERSXAcn8qC79ZDLL0MTfI0koEK5
kz9dedyJ+aE6xQx3uR55AgD+P2CZ6AuYL39uRVdFxZKjaJcrIPHgkBEKZUCePFhkwGBo7vDFe+Ln
8tugfI+JwtEnzZ9T9RHr9lQ2PFFT/lEftUfXPfUEObM8mf6/q+ZvEohAkUlQ909J9vZWFyfpymwG
48H30xu/ljP0q8LaohhCjQ/Guq5p2IFYjr7ndXxN9sWTKeJWDUJfs7Xri1Zzd7kFxYwphD0UY1Xf
sOcIWnhNs/R1+h7ST5c0+xj6eN/+KPKB3Ed+4IECZ5pRC3lPsvtpjNxI2i55Bk5k6wybpzFPeSMd
K9t3jmfNIYgkTuGAWy9lLP8vbrhv3XEIweBnmNsLdSYFSK34aVcfPGKs0mY4azKxA7BWfmlczYgy
6wqdcsg1G9ZhDmbe/HzqA1Qbz3Xi97s7gSdcaxwnowGnF1/fWcAY38ZKe34J1udIOMHth3rx0+Qv
S4SHi6a3CXE96M05nok603Y014F2cU2EwSRaaQoMf7dAghX3/RhRTHNxQPaujLuy2VRLp8TZ4JpQ
KUeVMukrSGQqxRqiTb28zeAnCrSy8EhEAw1Cfqkdnz8lmz4S372XwpfKbKYPDQ7DMVrQlxGmkc8A
oyxe1aET7bNV49EfM4+Hcfwvg10qwbfgfK7bepUb+lS36jNL6Wv/Y4F0EtvxeQKtuAzhluxZmrEP
jc3ddgPtahXM0s0y+Q+LjqUPP1dIImQKDRv3ZOkCJNrSwKtrlDtG6v4hlXnDaQRQUfVWRHHlHfAI
s206YNYD5Zbren44EOIcKlsiFfHiff9for6BuBFXvOkBPeNBgOqcCYHwWNxVNXw6/VXv/nU2+YsF
3WGlKCdFF3c5LhZZ4+CapuCdlFeK0tGtSCIyegmY41OnOC0Rytp9PbJweZAhJnVXOGnND8wadMoP
KPDtqUklF5Ki7tyA9jyDyNji8N+qDjlaH/LZC+3Ee1p3DF1NVQ7x3uHky02K2oC9vQUZpfTPeP3M
WQT3zH5B5o/cUd5iRrRiHtaNnR89t1IaHl+yFdHjOkdeDWfTySPpNoOYneT0h1iO9c2oa5iGJGOT
c5IiIKxaPRSS/ZmplQJHjtMVPl1oNjwMYD3tGFrSSlMbMHjKDdcx6lFn0A2Mb/VjQHK4fLJMz479
Q/pVAxoEz3nuCl8UT0i3CcxUyHYdYo5gTAIIjrKDGaCy2U5uBrxi2AghuZnN96OvioGpPN246p48
aN3I8Z5Em5cxvHZk+USRCiMdD9ocu/dkOmeSwoSDpc5JydpQy6rOKEttvaoxbM6sM+msO0mPa8sf
nvlipIPH7aB4IZ3+jbh3F2R0JE7zEPBGL/vHmtwC1o5kAJHoYhXWptN8RtPuInUCK1Vc6eQxzuTI
mSgkTZRdPdSZNOs8SmVcV1iHnQ3Pcf/PUBWSuaWyzLov9+60WlnyJcz/dpFLbvkY0cAOTB24A2/7
+xWnNo5NFxU/q0/KZPDyJ/9uwqC+/i8zimzjVNTXB82VJffoXBrgF0sujRF7eA0X3wD2Ile5/1+o
vgx9+YSS3nOiM+9XZbvX1NQcKhBtUfDCKGiz0vvtyQPCC/cNH+nQjrVlfClGIi+94SLWGYZdWSDJ
VkSc5HD70JI+cw0wJoM97z4w3DoujPoB8ii0LzHfXGbestGH5dkd1G6pvlFJ9IcGXfpazjMnUIbf
yIRdFa982DU7ONy/AfrHExvdWRUSX21HfFkKbm1oz4UGvPmg0UtYL90tsx4eVdXblthXq2bU4LsT
4ntm8VpbDEC7hf400tfnHFTTdPGJpceUdpLPcIla1oBSn7CYJCvIb8LC1v/vziLEzOPZWRxAGT6y
BPBAjvGw18/qIGbmd6PSy14/7F0Zr3ItpSrFZgFyYPi4qykOqA1NdCJR2VgIqsH5nF7UpgGMJX3T
DzOX/XrQMkPdaJo3oSxrtNCNlAkR2sxV6PZAidk7P3ouDRsMp7AtIAvPbVMXqiqpjX9tUrUpOy5/
WhJgWPt3FqUvDVWWPlaS/l/khqU5icnOiCw8+xxZge/PBEFIUIQFD7UVElXVXOKl+J2Cf/eyrXWW
ZNIubS3OiTWr/l7GAazcgUbRVzumvWbFKiQu+Y6JtjNsAdLqGZO5mXQVRfJaKJoTsRPrHlPjeItK
fOMMsGQRV8XCs1Vf9TjUlTRmWrFMgq1JYWSZJa4M3muooxgKzzVKXa78LNWA6fzbAoDYZRU8aoyM
jZ+P+kGNRWLej2bu6cNvgZkoxsCJnW+sGsyvJePFU5+d1YRtpUe8nowlu4p84gj1xdc7EYPhM3Yx
ropqtfn7t0xv4zOwMaWXnjSzC8dhJUZb41x+WRhbu0hGEubUeAblxZjPJAAPoL6YRHFAmZY9J2fB
4cEbhRDm+7PGLyzH8hwffPyCg0uMJyGdUYBwHn53ssv4ET1R53WxvgouZjYW0zFAoEEC5SU3c7hs
OBXWW+H/2wy799AAGe7wkzbQBrfm2qQX08ORc8XAsR6iX2VE/i+907e6RHdMehxPaoQW3OsTxAP6
O1tdzbOdqpBoASjWT1JtPmJSvM4Q1MLQtn7VZrDQbUhMP01VAEuY9dfwz3ln3A4FlUekvfnO+u3Q
b21soWdMjzrmcDgDufF6ke9SWHT/slosvLbxeOwwL+y+L9Ys5ArmY0KiPAaQxn1MKoogt7IQwlHy
beiXZtcUMImQLss1IFsAf+PzI0f5p04ycPYm2lQj0cpjGnHURiJcgXUEgqu29Qc3lBT/LJ8696nr
dHmvaxoP6+Q1owjf0WRH9suuyH/Hlhx7deDbNk9Nkzpa++TwtUhwIqVdbSTT9jk0wCZAUEPDubpN
b3F0ZY1AhQRSLsTHIms2Bq9XhemT+KMgk4rwgaRBwYne1GM86pvfy6ZTStvxL6D0xVEUSuanaqYE
wqEczs4CYLSO+a0f9xfgfC9CgqGu5pchk16so9jKzkx736anfgjvZupnA4RQLnX5H87pvdfzLOos
IpqagShbIAMJb8xm9D8sT0ycZ7tNCvFT/dLc2v6EfXGlj1dVP9hhAfEGGR47j0+W/iLzb6+62qVa
nUxCkZblKxfL4ukAkQdJRppvowHhJp9ddugL88QMqcIfjxZAxYkrU5g+17mSRDlRgp4sOaiK26cO
aIPCdSQ0Vnpy25ZkXAuIAxhJDYLJ86WdOqOWR5dVgfCRaXpkW/LZ5RCl95aEj3mGZNYUPdaoLV7g
thSRexIJLflcDYUuZBir6bVc8ej68TXlOnzziKExKVZZN546yNsbAgab93j+1Vb2zCu39O4LdK5F
Gp6sjkbVBBBB3NMJYbZNRku+mbAEBEW5GotGHCapjhI+Lr6vcnZm/IpkO5YX+8fV4dmOT+ajLNks
V+O1JU8k2sgagu1k+qLvruMN1KawOaZQcY+Yz3v/ur9Rj5INU2LpOE3vZOxjdBhFJZV1HvcbYbe9
qcx+/KtBGPysg/BKky6OtGrJudAuQ659802mxeWjiuqzYlHVgMYS5gB3GBHT17w2o3hEU3khPcJX
LON8If6YgUGpWsbdAbQkcmgJhrudmWNvKLazG6PnMz6cgShZxIU77R170WWilMgMk8KlIWSdsK3P
x/xzInEfI0uLAzWWiM3NkQmG+iU5N0hvUn9toUZ0p63vOaMAGW5r9iIe1ZIkqxA4xrfxdRZ32q9v
AGv66B63/gvaoaywxG66PFO1Ds929nHLuUsHLm6pPPQKmkalrIPlP1WGfFhBDJNSAbvNXHFQi+OH
r1Vbat4DCgZxNey+KhkzQ2Wa+4iUNYlNatXxssCmxrlnFQDC0x8zXzXSiaFtiGQWFZF63j5+/YWv
is8FdhRgjA+zweZhct5G/1corIbnYiv252dhACmn76G/TPc3KcKa2/+5mbutU0L9W1srfwn4DeB6
Zrh1cZC+4E8+m6A3hkYoTLBe2P7ui5HQEhf/4oar78GiDSvD/xjRvR8ctbCCcTSlbPuwrv21xYWv
xiWD+ZxBVHgwW8Wma0cip0AU7rSNmwTqgVQmfJmN956ymoRJ492VCPAPxHqAXAoY4JI12FUN4BAt
nvuOiVr2nTsramkyeJsnbNBvl8QeK3AcpheLubw1+4CEYKTO6og2DpH7l58I3Ljrc8Q0LaOLlJys
wRX+2pZ1hqpByGYd7Qq4kSipEO0kvwtS9V1WghTvfkQ7M2dRpDA05CesEidXSMYUdgKklP//K6F+
weqBbP2WHeHzBnBg+KRDT9fw3WB2hJ5hjOBCJtksSqvCJeDBMw0Podf8bb+A3H4/jfDhK/x+oz7Z
g8q256KWLfmGgo7Knlbp5bcVYBL6Kx+8+gyCaueV7tMb0QQi2j+zshS6OvD8lkvq/9vITC48zrl2
zr/rqfTu9xNvl4c/WSTFa7cTBkF3Q4tITcSClWQlCtFC6NphqenC30NWR1y/Qzy9y7peTowy3j3m
SszZCtQNFgdafMPre07v5cExn9BX361QDUnbLf6en8Rt4yCNgzrzdVGm4t7axW1BFGLdSE/JoURY
ARLOcIHYw7PE+HL9W2xW//0F/p0+YjH7H35KmQ7uKcJcy2itRRZYQihEFxly4b7GFpZ0Fguyw4AC
yquQDAEcngmUL4v99oW2U8xU8zN8AMfGN3Jf26//3woWmN/U1LEfBRbLxnq5tjeehMyeOFxz2lb2
UOsyeI1+tYQfpoQcb0J7ppKYnAdz1crBpAGoOKvGdzeaq0GVLci88NXuhlEoxPci1jxJILR36MPo
IeG2ELZXB4KHK8VfrH89zEfOzvUxLnCnFyTIs034ESVj/EhADrihpsbs5DA3p92gIkeIXiNPRYvW
25sxUtz4IL4UqqUIzAa3BLvfiuKEm+DAq8pzdt9+Qap1w05oZhgX3tfdTWlOGTfRvwoeez0kOhtk
alQPDNDLlmX7vGOG9MokxKKeEnT8ffybeOpca2ft9/g2RHIFz+7iE0A7/Pvu35azKxHXYhuyq3bI
w/JsHGNmBO4zlHHR1I2eQiwjJD0CANYJbh/fDiIf7ecaQeVaEkhmt4clTCykO7jh2O/HNrTt3sle
zbRhaWhmFaZcSJYS5n49KfL6pp5y4tlm8Fr2G8VlHd85IFfGdX/RvEeR4aeivbU89Uk5RvySK10j
o8xNTx6DZn88nsZ3Mtroa4lIwXYmG7Gac6pK2ScxztFRCOIRX5AR7pex2YXVSWqkMsl85ZN1dW1K
lgpO+2YR47FCq60Z+R9aHYTc+1j6hkDGwX5iixf74lLVEms9nyNLSgvkkZqRbBI4O1uAS77Hkt89
QRQLr4OaZ1vP6C4BtiorZd0Le6yGnLUiFRlJTAP89y4fn1mW7EqKV2gzKaTxJ4NJs9QGwsJ+SIT5
mjGZ5e1jeSJkaKJBCOQRGIqge6IbPoN8e1JO4/G9dNqWrcnPgspC3Yx4oIAWRHlZkKVIbaO8GB6L
xiMr9gKESt7jngieRw8vfoQx0ExKgyoPF2JNi6zIU3GIiIKiwIbpGngSTMv0CSArqrMw0Xzz6kB/
ZGF+S3IRUVXm6CZtXX8/IiQ8RO6jz1nVPH9cO/tjX9lOp/6d2taOihifDyDXhLU0v7ax3y8srIMG
qPQ27+x6S4o9ppQ0Ago68BFtps30O++nnDkwabqNXX0va1dT9KBa8IhAR/TxOng18F2DtSlkJZdM
wjqhta2t8ur8yMiPTPwDJWpD+ndR9tUPPhG5qVDtABoCqhKOeSWwAvrisPQmrJ0seEga0Lm3K80w
vGrvPnAP7SHYCosKr84vmxi447IGGJaeXjWUGagbKnf+4sShfy2HT2dwp88UYeqxE7riYobsjJGC
T+HSGeAYYoUSte67CISmXZDx8ivAR9xa0l0n4I47qRuzwDTVQqU4o0cqZ6ltfT+TruTfCeWsfJoD
9jGEJ/0//PlaQe+KbaYvdsLiB449+Fz2qgQ6jXZVlrlg1IasKMyvU8T4A2fa0I1I9eylqHW2+g0U
6CEXmlMNvE0FVYs5tlvfLW4qgcYbGH416bQwfFVDnySFn6ihlE0HwcfHqdIgSU2FoCpRHMmkaNSh
NtH/kBEQjrWOU/riIGvXfMjov5uMy+Mu5DcwAQf7u+03lBZAmBTjKYL3qnLeQFHrm6NP9WmMHaxK
s+TUYwDeouJAVgDlum9yVGM6gJJ+Dyolum2+obsZQVutQz1wn1zmXfrt90Fc414taDGm71AAsaw6
A9LBvVtoplVHR94YC97M/TejIcgWfTD8jlPceMBhbmpqc9jZfxKmHAElo20Q1yOAEMTvHx7D2SxI
glt3hEYOkQ1hhMApRWLrXxAOUmExJMbQXUtng55xFonuJdwwfA+oFzD+RxSWZArKWd0Y0H99e185
uTc7w0Yqhvc90nje3BnO8c2OybY71zRgmUpU1+FDs/adJXZjx33h60NyOe8rjJljkDYUFRawCRPY
AJG+GbUX++54mK25Zsc2aHo8z6CpsYrHUeTeG69f19QPTeq5a6RCYVQUhvqphiAM2Shx2MYm+vle
FMzHLmH4rTUPMrqP09DeDEs7r7GzsqrbVz7oTAmyYHQVCpVcrRmqe+KPx4Y+UvZqkd89o1xDvfnc
JCVl4DsxxAzMI/iOTxGSMq0nzBdt2qjERCEvx85y1SIJxREyvRyabRu+TyD60d9ckZs2KpMycsmN
opJLr2jlNO0yboXa8X78e+7Aoz8a5kejK7WNJyDuJtKxXWVU0yKS8NunhsAv51eGZ7fGj6Q1kedM
mjLbiKYWMaethYj7huzlwxsK/12kgquxhFw33mvdc1O56DDcffkpxW8ztsMHcdpYeqzQ5tyNZSRi
BAI3eTSkcNSVAXCGOM3m86EjBwNyiWLz/MriBiPeJDZZozkv0eq5L/TFyK48n5ukkD3t2/gjkpoN
VOz9y9hK+dj5A/2fHXb10DDe1eO2J65kQP+98OO21Rn/7T+RPelN9eHjtjlIYaozvFuL/hUZDVA6
8AjoGR0+ITnoirFKydCFY7c893NVX++g04d2PR+Z55Mx6jnufn3JzXxXMaQNqeN9VGCYFyXtnnRt
1Da9arLQb0bZtx1rPy5+YIj8BrtO1c/cvZefv6IPIp1O5czjYqfxCqujNWMDuRtzjHoQQ6UDHXcI
a8iGyJZOf4SOxUpmChgbwajczpx6FvOS2sDMPHIiFboV2LKiGKLgZqcVFYCBcPmEnMXyAkCH7GCK
x/hV6g8LkAvldLsOS0xQIcvAbuDEnbViyp78G0GXFm6GBf5PU13UDk2JcOg0u5qN3g6j7V2UXwgj
ImkVIAUdbJSHr9t+8mKnZpcmBpaOg75iGCQ3QgePRgWLp+9U5AUSUYyiZ4lIljXS02HTWxyvB/7I
2vDbTMvxrLGWh104txTrUwKk+0b5P/EeNsEMvEtBoKkfLX/TGxubyfrtw5Y01BJbPUVWFXL4pCsl
04EOUH8OwMER+xcbwqDyIwHIZk7LU6lgPy5O1s0B+1Oyo/RIGwo5PtkFiKZ8EsBE/XbGJGkL34gA
kg9JylsO27clTArfi9kJFMlY8uwhmbQrv1j/fAm4DS8I0a7Bkw/vGepLAmAkrtnVPuGszf7Gta+q
OJKZJ5vVur7WaZ08u3UwfLw+RMgYwClz/BFa7qNRh5LvqyaSGL65R/InvlvnDNgPdQ4YR0CPBoty
+mDmQMtnTvNPofowAoiUtTtzqt71Bp/Z66LDZ+Cxf1q3m1IDyES1x7KwZmtZSQaI6ynkE1E4bdsq
/bMO0CekoxtqxO8oPMi4R+FJk3Heq/Dnb+SwmO7l3gYrxKs0YxNeNQq3Nxfe1LuRMPHc7XU9XumG
4sCT0kFO0VF8byc9cPrSv5P4h5AMjVolC2flZxn3sVuPgSwixS9unH7V4r4isytA8z9qdhMQoLbq
a+awCqCBYMaTufKLXXnVlTcARl+el//jqSipqKXGu0Se+zIxwOoH7Y/WiFQgHRc8XXUCqIkFswhW
GUbUEaLOwEE8CDdZRX/YWC2dTVXth+YO98xeYz7L/fnCyY5U/QvgmLDGw5JsH7QiUmpXOgMRCBlW
0wOdjZKOcDpoXNlp9K6XuDNvNTWopz0DwnrZuWQqpW0pqY999p0p9RF7kpe/lUJXjR8wp2Hz4oA+
XsJeRS4A9YGZr834As/aZtGElGn0znMaYusk+z6ujV/jw2RNb/5NVvDU7gM4//d+lhS5diG+QK4K
Oi9Qt0hxVMe7VSUEUGDQ8esJZ46e27u26letdQDIo4Fy+t/mpJKCEFS2psbqcbMBA2kFsk4E+Hb7
8GczaY0aVwZdDKOd0+OUADpspmZbnSwIf4bTnpO2w/nsBKrqY0zp8x9ImTTGKKLNsgGCezJHiW3A
2JpdKHqAfYmzaadfic86Lq8htIFjY71vG0L+glOw85nyMOnIh4oMtz9wQCpDoDV5jRSqwDhEDWe6
o5lfv+l/5NxxnIQvUykswQOoQ3i8EsScAEL+ILNKvW/yhhaHth3LkjV4Yc5v/NE9ieEynRFI3r0v
NDafoDwqcZQad5N2IPLYTQ6rpG85ms67zYi+LO4h+LntfancuD+czo3rz2Rysn7S0Bx/dIkhd4uT
fpU5agpxpuKRqXV4/g6nUH7dbXvKCPrapG7G6Jsp0zW48ZpiLLVYGt4PBQ5GGlbZdAYLD0U/9OdW
bvM7BX/QDr6WCxbDzVtM97wDgU4ANZaQbb+jWlXQCGf4rmNzO96P2dSrVaeSAlguQI5zShIdwrYm
VNJs5xcNfE4BfjOWznkBIbZrNguQyP+CfjBwgExAjIco63Ib0D88Bp9aUL+hgEBfLdF4BP6k+wQv
LiI9Jb/iO4RP7YZ8kjQRPpmaQoB45dsqq850K77heT0YmIeMIq8J3mL7ernQ6mUz8o2uRjqcQVF7
KGYkVTaX0HnWzjWll1FAe9Oj6dt5kQL+j8iAAq7ffqX+UDWTzlpRTlHgyteSsNf/xTAzi7WiIdDJ
LCD1VHRkWkARfZK2r/6C7ejer9HPJNND4FjoL0B3KcYhhVCd3K8ci8Wozmu0GDYFQUZezuzvv7sH
oF8InXCkBuAP0RqlrPDBdEJWczkGWGovufLYRv1dHwePboA+U9FjnSmwoIyxjwUzkhMG82XmJT+3
Rwrwq4tRYA+fQe5nUqQkOD5XnU2OCBkfdzShiGhYwVRi75eXiMDkONTQrCitRRtMyGoWwkNwIAeb
FbxIeUqQp3yv4neHV/1GVOrY1B34fBNjEh1LubdZ7IuZuIufQqB8Tj5L23P0IcmSGXjtZzbW9XAv
CaIZ0PrfEAdjeaxIDXVADg80JAbngFfaQWIxrJwdWb9WkGiO3ZtpXSch2ov2T3j+9oMKTWbIqoJp
dd3MXAChRZsJfbXPYaeo7MxQp4NB4fOxv/j55kXCN4DwjeYT+ez2OswKOHQpxQSqLty8bmeRTF8f
TvbbLcHExBdS+LYJsPy4R7WSry5HJNtjNTAgdICQUfnFhJ0zE0hsGnwdzl9gCq9Y8W8jSpomW5fl
lLxCb429T9iCwcY9INpAGZJhr7sWL16W2IdMzRLDXamDgDuHAbAEoSVs8Cu2EXiDbul/NxJd110v
zf/87gCmivAgbOVI/rprogftge0ls3JHn6IYzoMeJYZbP4feimiRuNWFz46pemsDF+Dszba1C6Xs
muv1QKWcivkvOSlVsKmss6naUcsrgruhz69heyKp+DuEZw1CEWVCtCpebIi86GQ2w6PuEUNyKfGs
t7gc++MDqEJv1Pydq/JDhlhzY6Nv3wFgDiLSTDl7om6vCZJbqYF1idy0Rr8TmIZTxuedjWQyGjpH
R38gmC6TMTReE/lUePucvRWqrSR9CZrHpTFPKJXFgVdJUsYbyfPDuKzV9syDQXJ4k5f7lZ9OZust
ru2nPuNmF1DRt6k97KARCYeZiKwzn4xthUP1FcCIYqqccIS73HHLYRPnZu2Kl9QXRXsMxmyTK0V3
5pz0G95hKRDSgHv+iloR1p75kp+i04mE38F/PZ3rTHzl/B0pc0lcNCoAYt1WwNbxPapJ3PJTaNcx
pIm3QRKESa/ZDDtB/92Nk0DRxHyHF5VQFo5MVGO2kb2BYrFIqgj76stlZYMxuF3TwM7+mNqRE5LT
Y8RQzgYDVXwrS2ShCCDjWqJdR76wbQkhYdfNtnQNy+5mHn8TW5QB6RCxdVSNaCbdi/RtyQMViw0O
SuvakHm4LbZhCghs0yTJUVZuQH9VaMAZ7RP1YcaBIY5fcV+SHd9aWIv87xPWhwVsu5GKnbxpUtLi
RjdLJpIb3WkL4hBp7jxqdaxVhWsUYjgCK7MJd8nTok+I4mJLIA9z95yonhD9GpJJOBU3ZEzuVqr9
9VFy/c9sgpxTxeqUIkRdXcKkuor69VikMU/VLJbe1jIriZYpq0YF9gB9yod//EcY+G8RTcqGk93l
WrMZi+4Qfr2KCBv3gkuy5XdUmP17W6jO0ldVvLyBUzog6yJB2aA6mvxK9w8ExquFTT4/F4IGMRj1
LLUZwrskfRD4NZeg0yAYUyP1r54jUboIPNQAlykrURz0AAwJ4+/TJyyRLlUZsuTpfSW6lnwccvOV
/UUrM2Cks6UUg540Rve1dB+Qc0xKQuCTeEBINjug56BEQK5bidfDQp9RLrNujMVN0fCVZHR16K5z
P6VLCxzutjj41x5APzWqGCL3m/hOOyyIQGVMdC8DO69oE1NjYg7DCTw0XA/IoexafR1ax2gjHjNA
BXIVjmZVsI8tYJgpC4K/hEVRs9BaeCPfScCfmA5WBr7Dra8rJMwaVDL6OYxpUtFspvE3+7yrlNy3
ZNnISqkSvvnEqWlV3bcHvgsxdi11ILCrlKT4R3b0FInT7ylFT0r86QfPaVKajsmt86sWP+Q/Na2l
JwIYXjDSelOqoFzy5mMqnPYbvPjuVGMGMD+4pXm+fsyofg4rrs21zZWCQw1JTW0mjkW4FMJj+F2m
r+lI7Eu40oz8wSnzBYV+DtLfYFXhZ7xVZmXXMkrpXqgiFCSNLvlJ/Xl0Y7KyzFzcqd6dpv5x3naP
axVJgYceICZtS1J2QkK+MZstjHSfnJKio1pTEYDd9t+dwYIYzEvQTYf/gShO7vpReCk2FyHkmWE8
XBeQ0qxEZ/evmX6tEd/Daliqtu8nDtBYgM0DqBs4JYTKadZxrutSBbWthvAg1gPIlERqeMOTuNSb
mMNdKfHSkZxni8aGLYurcVEWvvvw3PvYkxW5zIh2rSCix6l2PcUHpFLzgP6Ie5KWj7VOD3/AZarN
x35j4sY9OBzkWDm2p4k7aOB99tp/T/Tih2bcqMt5Kw46BnID/jUDBjNJzB+db0SLvFW/Fh0HPi+H
HjE6r1TTyQ4NMIS//hyOYzCaQAAa5cmrZO7ejhWUKiG+qHiSchASVMDp/TI20dyb7YfKtUQGENN4
NxGWWD53B7xFhhZlhirH/exjokH/jhtG/KkZmyCOp7k3R4An3o4FJKdJSFF7q5OB1ZBm9hJGSaSN
IMDXVqtC4lRUHhJ3nUvQSrEDxVUjvmiXvs243I3R3hpkVtMDJQ7mvQ81aUVj3LTxGF1l4C3yBZDr
dr3+sIEEe+vg/JIfmaxVrX0ayhJ05uoHUESoRjMDK5jCUJjXjzPEvR+DdOKln2+Jh3wUj9sBq4s1
FFKLykuvLOUSdGzoVcyzECu3HLmW7YnMQ0lATN7xFkEknuoKmjak59KIj4ETcUhJXjm8UDN3eIR1
QHsCVmRHLXchuqSqXKkaNtkq/I0CSuHe1qTZwje3wB5jjXJ4x72o/kyf6YUATAh5zkkXdpphG2Az
e24JCcWBMw9/bKiLAOer1SSCWZAkD65AwGEOK24hHK1zXdJU/8UUYTQceF1ufOUVlWgQbgciPuvX
Xtsx2XPRlJkNkzEb/40XHOR4o6iN6H30OeYXgn198q/CuDxL7YWQC8lumGwQGRGghGVZ9oM6iq3K
B0XL5I3kRnf79ijzqxRyiaTMJogNFxntd8dXUOBbUkFPCnrdoc4Dt6Tu17CwJdZczv1QV4UOP/KN
zUy7Zurj4IT//wmxmfGZJosiVfmGbpiOzM4/oY9m09tPwKvmS462vBIjYdyo9seN7+sA0EH5P+PH
hiQBLRXBQmhXMW3pIJCoFdtzESnm8/CDeT+gSY5xDr1qO8eS4dbdsYe/LxmFslbWdQqEeVXnEpYv
02SpNQF5hPcM3IUy/8T7Y5aID9eLG7k3vhaPINyAE7vjqpYby4PSgmmEsDyEXT4ABEZr6ahQAD5h
U6NQDRO6qXGHC2cu/AIb4/EosgEYD1unzW0dK16gCBTOvnrOvUQf8tn7S1yizZLkUnTLGLF/c0Rb
Mm5PEEUquJ/Tep9+vaE3DI8LmaMeTnoaUG3NwviKb+Gj7Xt9cNrg810ym7nQtWf+oo6VRGhkoX/m
QcCqLW/Cd336qApp5YzwDBHwLEY5MMO8ks3z6zP65BSDAE/0b/lcu+0/MBYd5weGs0dJBXpzI/Jd
+7fW1UuW8Zh2XbOFRV0Won3rqRJZQEyJOfuQ54BZZa+TjnGkZT4DQ0oTqLsP+ToZSQGW2M/FKOXG
zOtTBu3NTJibx9ofgItwjLtfQQLMyihwA9a9VVKRIugNEgoaMR9GRiHFDSbqX3jtEiLGke/kVh3h
D3sRV7g75V8qAWyCg7Ow9B5KPTP9nIyanXge7b+YRfEPyfrXB2sN3Q6dQd54T2JXYNvTsX0sCbHO
c7hUwOtsiDhXc+Z6Wos6kVlnEgTu1Lh3vGGL9YfeR+2yKTtexwaYn7yYcyGo3huwhQKgNEiEWmsl
/yCic38/1XZTO0HlFbPQq8qioVVFn2ub4spOz2sUvXl/SZY8G7Uh0dXimSKKlbEiG/ivvF0FLB+F
ngo+PBR3H9nAmnwiIH10YAAErDGlHujUG+QcIAy5YP+E2lHX7MwuxO3f/LiAK64KHJy0i/AZF5Tc
xBSYFU8+y3kNwQQ8oJpfckOdy7YVoi2RXSehVf5N2RFrAOuuD1YhC3+tz9fOUx3WhTNrd2llBtFj
LAl5tkyx7WgkNwlUdFXX0+20yKZxduQSR9zO1bb09U7oWnLuvYXM8t11kqmX4bk4OoO8MyEJkewa
GTwozsOSOtRRJ92ILfpCgIOmuaKdK+2dkkBIzL8L+pX1oWf6rCQIfgRn7vFmphKPxq+L5I5lWttO
sV8rNMUhEhxSt3xC8qCXXOz5D2muQlRoo3e9MC4lMRJFxIs/0VC/gm786TiXyPnOkgmHnHcVlXI1
YQIUahJvppiG69R8TxNacjJsMluZgQ34BduR1589NuSo3ycCe2RWhCTJ9Jvib93Lon2igzApiTEw
LzOQ7XyBj8DuTuoStfIqUZ0whM07fA/+ZESYlQXZFgZYW5qdoQTyBuqzUI6vhHP1soYwKrNQq8O9
F1nhxz0CUw9CdOUqDhoh/kJoCpTmOUCE2y5bOvnMJtGFHIFhiNIE4r58wYdHSMrqVu8ZZMhYm6ZR
YAhBKiFCfedJDkbjOowKDhwfHi+9v2gR5Pc7PAUIcd5/pSqizHeeHT2RD/pEB6epHfJhgjb4s3B9
EavDf8v+nSK1uKTm4POC5BmcO6tyPOuREuYs0yRXnJ/isZJqyUBYGI7nqAqdiEiJaRU82pW+UtKm
RT+vop7hMpH47izU5DXMUNI/Dvddr2H/LHAhQCUR/G7wCpT3dynssZdQYw06WP9cyNDcVn0liwjb
/W/EIOX5rSIQuyc0kwfTFT0rtH6ML9IRyPP49nh9BZ7t/E12rYHnxn297/CIPbqRvz8Knmk5EDNS
pQ+bOKkfY3+lmd44Cs56LH5zd+pAHuJcsqO0rQ3Kx3YDLzDlg4kaAdj0NJ0pLk9Vik+gb/wXnleK
JqCZNrc+s0AvjHTGoqPoHon8auZtAnifFAwCn9pa4Tt1kmwKltC1AJvtW535RB7o87N/71DN9ej+
jeq5TOUcigxf+zEEuZHusvfoa4dD+5SPgMruzExlAr/Q2anA9keko8KkkpQ0F9H7FBxohadGXppQ
wuiqj6b+OVRP0pSN/fi/iMY487/CxoA819iFb7O4IQNY+9el593FgO4Dxftf+mekYnMdBGQXiEax
GUfSLxwRYGzzmT2XqnJdLmCwnYxyKHT6cd3aeinYEBEk17cciwuK4crcUqTVysT93YdPU5n9Pgjk
r4ZD8pX9dI9elBfhp7k4z41O534iFnQM7dLKh6MZkfBGzDGVM9G2NNbyouHLM0TjO3/Zg+Jbb1R4
QoSGP3vcZ9pmfxthB587NIUrkit48FTeOE+OEVYnesXa+CKZvfKRTNvcp3tCbadd6uXivRmIE/rp
hXn5Ir6o/EshGKVsniGH04i8FNgE75uu7iYMtdHJpxcjs+/Lm5UBzReaX8j856QM9bHYCzlZddvy
8u7BlhruBPVFPRhYTs6mjThrgeyznSNRCUyC1azkV9+Hl1Vpwgl9wVNXG74ZrD2xk6yk2HkEWG1f
os56++rRFk3+H4Qj0QOsMu8eEkUgrsxm2cQaQ7TkVmMa7TAjbGMoUZx9/oYI6qRnUyHEaQLRzFut
v9vHTq4BXFLtUIdoAR/QQ/EwtxUnM0vuSeSa+RMkpz94R17WBeJkwNaUPdt56EyKk6Z1ZF3B6Pz2
ivVs/P7KHe5aAlNfY8apzIXeLSwMlHTXhOlQuOr7A23z9YVvVGNLkggdES262R6gIwOG9ZEGtLvS
/wgz8RkcG7PjQSkfw8dc3eLE1sBy/Bs/8Jw4W7GnJ+oXCATfu/AFO5aZzkMme7PC+yJVQmBT3rH9
hnfImA1I8NfcOHcMeVowqeziv369X09QRgUwu4iTQUMUrQU2Tx04ZO9JfzOa8l+UHJrBP00ddxqk
PGTQskGb1uU2wywy3DPRNQrIGIaNsFJBETs8w/p5afTMevt0XsFOCWB3IZtgRB7ZoYHMsZpi0v+I
Tz8kpAMD6ZC0O0RIlupL+OMYPILa2R9UciOd7dMTmPYRS+pVDu34a7tYWfmR6nPyFMeq5YrcPuAr
bOPOEx+7GaCDhmfvgbr4h7WSpoT6xEI69719xVR/qget73m1StNJV5JRes0fTvFFUT31Aj0xZGEx
v1MUsY8V6BJaUmtBWwK9K1IsF9JEbRlXVZyH+zQIU+Ay1zolP2GRgM+AYThXu9ABZ206+XSPLuW/
MGOELpNQOyvEqmkaSMBIdwMJMMpJFnZf8FX/j8MmiRKVpGfFzcWJ97vcgdPgFDTa7igIk+dF008Z
lYYgSGFwBIqEDZSWkzK7BxYYIAE/4oDU6iR+31JYUPiyMTcWQlGjfmaI7BRjURWPi8/vq6GhSXjZ
lOjS6Zwu5g8lYbkN4s8rYW2MkTfVN3L5NBdzQtSU3cVSwoR1lLN6ZlzfhkmE9++6Cd9B2PVAQyue
HCOSkHXxPDq9LtF0grxR66DPcqEcUgN/l/bxeyy9cWiPm9wKqLS11TesfgzN2ALk8+xhTeTFSNYR
IJp6WnEg+C6oIvvdI3iV2HNtQQXfDJuijw+gjgZK0abCZzOiwuuaPC56sI0pPj7LaFE9nZJ2ccS9
QWn2AgMfH/PBEFCfJoCMN3suL9mjD+u/938ruwp9X3BFKrKjoCQP9BsYHcGmBtV+A+phMJ1Udu8w
RaL3YzBbbAPVHrxTa8qvTBfwY/MvUCR6XHr1jtE/jMRaqngVOHkQ9NwXt9T4cziKTNXcgA7zekx2
qsvSiaLbi36/e/I3o0dq9wBfqtvpGekSIyV4lrjSBo+tfkYZwVs+VU6lPcEzPt/ZSoFtXJZEelJj
i68+xdlgZ/McpiKI8g3k8+AjlrRTAP1kOW6KmnTpv9VzMacLayWngJJ1WNAVHwRGgvu7NxPTVSLL
Fi8JR30+RKCpKQoNseGsMirym70qzOmxQPumsDOIx/wWXsyQHx+bgnTODUCzsV/FYSY2Gj8Ako33
+WPOdcHoqtdq6n4XHu5uPrRQs60cIcuGL1rRA2g0Ya4QNqZswTQduNTKvQJQXCvxxBwyVK7liVW0
vAXfNKrRRymZqYqZEttfqfCpnUzPGxnxlFZ0VbTZoYIIn7v4rtMf0WTUTQAiIxHy56dH491IbSxY
a0hmasU0gmMH4UizLVP9SmWBhKtvShfxCl/hYz5+n0lw8l1BhV3CmXZBlUhFPtECpzfnEk4RWFVN
nCKGZNp66EbPl1s+9oVl4rama2PnWWpElX84eqUAEWbHFBG34SXpAZyRmOIFHHFYWf05GWsx5v7n
gN/+pzEINuyyAiForciOEMKno5r+vIx/LJopo5zXVAfwWOREYNCcjhAMDqX3u6nKdXvYBQSp+9gA
a3torE0j4XCD+BJn2Fk34U4pWlSvOE+zdEdukU44+vtJMR1ByEgphoO+S02M/yyLM/DkxzJkVOLj
gzmEFO2qplf1heWNvj8hu1ub7R6vZM/cnCd61TLO8g7SzakoWWi2gbr5nNIwPsne/GQQE4M1HfGB
OLYWrgfMq+U2aQL2cDonH3gQltLka2yIe+Nho3tiEBLDoxFhKGYVeJMQNDw/V3duWGW1LM6yvJeT
BmoDFlv71i9UyGC03CiRq3PXqJ78JPU70ob1F3TKAMEeB0/I4UgoGRrPrwF3XM7ae6E7KUGwTZOO
nTLtpodo8sa8z1I3JK6a6L3X4zXoM8vpLlSAdKxzn+E+ABcppJWysvPL8jTJtd79QFC784aC/1Vl
BKZoGVY35eNbpIq+3pta7tPsSCUDwlFGSOkoXdh5Q5DLJpFuGwwNXBrakH8+NYRdfTRYoZ08Po4J
BuKIBwrqx3rCi+a8QEZZ94GZXc5eWWKPOsId1eAJ7fegq94itfsV6Fet3ewtUMNxuiWNRCfe/zt3
2V80+YRSsKuVdzMg7Va8hBeFjHYWKdnjtIR7PV5b2/efhaj8HqIIB+AaTN1wqar+uRZxofUbnqPa
YyJgoAftyp2gtGXQz7UBg8UeuCfqs/3W11JMQEk0J+eYAJ3N/6dwHyXUsZcOHHkBUu9vXptBgxqj
TSbqN2mkZOUSF2dBPXBe7aaDe3+rnFKE+wp4ZKBFXTXhopvGXLnK7ezZO3+VshrCKQ+6M591j5Nt
5fx/k2m5hthnbuIMSaT8yXhSpD6FobYbHkagqKqKGUDpqCcksK+XkJx53k6aLDnDuNq33dz4Cbhe
yD1+KGCnO9dmSZi3Naareks6HORYHNE87Se/JV5edox5ULWEoecRWX4HmSEDgY8JxXfj1e4myDl4
7Kr+fyd3L2EvciaOBWrkV+RZlec3aN0If0ZKZeXaCV6uXyUi8xGgmlJi6cjfxud9/6rkVVIpLOn5
atxTxmzf7wHTwMzovQGPmGz0OoMia9586j+Q/qLFnTzyl4I9mWb759sOD+AbHOLd6P2kpF20E/Np
IM/ppLkq9zNLbuSe8mcPWBd48YkGuA5l5j0Jq5CyRYZ2QB+MFEDBfbN/NuPi6hW/dTJMJhNLHef6
jW4RzANf45p+3pvoc1Zy+d3nWmu0BR9r4S33jY3fIMzhILVxc45YawRVrWhCQGPoy029XUCCecYn
6uIUFkgkifxwA5FqsiOyricjzKd30NfQe9cpz3y1Tza+38rDtHoMZbog5Fr8ryFOxL67FKfXxRoh
8FVUE5mXu/ukoOdxAFD8d4LXjbCtcFO5keEGxyiIBc9SFyRAlDzSPbQeY1dU/zPQMhOVB3SteSAp
zXnONpLMxhd9rsPxO1NcGOM3SsKRAQNEJNoveyZkrE8+ZiktEoHJYIS9D93mtaVs9uxIANfdAexu
naXI6proXoecZZGJKplNJ824uevkN4Y6CFm9ACIM3UHAGQ9+8DDD4aNudeC7z14dvudxGxrAetfu
pUdeZBbn21gq7PeZC/XEAwSbVg5/FtUkqE1pSp0VAVnFlfW9jrts6K71jJodlri64Yihj5A2m3JA
1I2HDgYGmnE4DapzhC4CSFIGBgD+N1Wshk0Iz3apxtZ/reErUm+ugxbMDYTihytXKVCZWwkl3Fae
y5XmkDym0az77MFvTVRTgI1frP+TMi0qCGfvY/9qxMdzjXo0BY5hpw+qwlabKmU+Glbk++YHu4oq
eYy8RtgKJLqXn9beEisxOwE/JuQ7axl1QQFOWaJSTnYJjyLxGYHl5jtXe6BglONcci8kaHhrRHi0
Cu1D59Jr3nO2FdglgqICN3+inYmt6Wghe4ObuYqASvhnoVNI/pad8FAAl7kBs405Ks57b91lo+0h
qc8MolZ4apU/9ixkbNaI7vFMQCzPj1yliUlFYv5TUhZZ4zceIsvxFNnZkPWbMQWSdyz7iQFkxDN8
m/yKAZ/EtIygZZkgaoi7Uiky01ned/lVLHMi+QU4vo6lnvDTqh7ZHIRjrdr9k8Bxnl0lFbFiW5wG
HP+mvjr0jMghUth+uOisflemkpfgNqoUQReFfmZTD/NLYUzkiCOas+LhZVuY2utsVX/NMo7+Pxji
PLMPLd6QK1dzh5gaACTQ9zMgEU2f0+ArnTen2JBdCHuN8DkAUyOafDxw1cDhLDw2KYeyV6OdsDUv
p3dRZVrIUqWSLS4bSLe19bLFRKoZqnpHfAYOYlRJQhSokSFEAhmRr0R4hMidUvzNdoPJLp/f/y3I
xB7w+mg9wg71BtADECkwP44M4nk//X478k9mc1gRdbju4G8S6i50EZ9jTbh5JIvjF1G8Rtj3Nw5R
uMLr2cqK5k5woIXcaHCauFrGQ5q+xNNvBm2Lb/luehTchubdtaIJzdIqJq2Dhsb5UsRtpihAUmpE
BsfZx7G5Ija2IjPqDz31M3ekDc17x2Ii8bPXAQxvTXp6LF2yIRc9kH7Q5z3nH6gjIDdeuaHvhs4e
GBvAz4NaMkKQIS/cAyTmT2sKl58bZBOEW2PvQbnoOhAdWvCj5PUybgyF7+T5YrWoFwhZMfaJYoYR
geDb5v7Tu64u+CCw92AKP0Ik2cpGrvqCYLoRsJAifB75xCJKWOoVWlzXgcSc44sl93TRFXOUQpUi
LJkXqKviXzYrIn2nEGsIu7dF7FFHVBWeCOCXXszO+x+kLRy4x99kKJBVhqI/YRZnxIBvEtW38/Bd
JL5NeYoI36pHYp8GSuh1Yomgc8Ywd46FOa+2XvgwgrlpTogOsTS/IfCPyU3h8huQniFH6WICLC4y
Xk1BKZ1ny962NnehZ0g7qNXHZPWLo+/dJn1Pr/1f5mBOs/4yOP/W3tB7tEfYY0GvJILFK4PBM2Eq
m1HJEUPPuplkM3xM3ptxwdtHGf59q+NYTTehaQ5uucYNsgKb2LX/UFN2DX+Pe0A4H4vRqoXK8keQ
dsuOJYxWoFgMKzAh+6PguBLgeXJmVt7Ooq3zoz00L5jda+K95NBXRls+zJSiziUX4unrePjU5aKP
ee5CAWp3ItCAnPWrzq90ND2Of/C6IEU8Q6ACT+AoqCUyAbqunRIhPmFZI470MMI5pBVNENBf4gvt
bnwziFhO3s1CU1rsJj5L6/Dp3svWu9IoSGeP/TpY4AUeqwFaGTWLCk4j9DEAGxAQuOEebV/UV24E
lSJ8QS1EJsuuDOMHUg5Ty5LyH0l2uEXN8c4AAbQacnz9Xrp4R5hsUTgUwspIlpjOkg8uWl4rOiot
phuFUbbDndNU8R4ub1BTWlirM9rh1ffzo5N8O+ZYicuaYwz0TWOkq2PU7rNcVmPdObSjrYvpXKwA
CctffIyfAy/K3cjaQDaH/LtGHqdaBqFEod/HYo64po2mW78NCfni1YicnISbVy2d8BLG99QI342I
PKtv4VIIt/w2ZVJ1Nv43V1onXvlln5F1eANHqQo9FB3+QGXkEWPKqucTCtdcT2bw/TKboYj4Npvt
7emjybZB+iA64rDUNJbFTbZrEFgRPpmKJBaeQgHh7/Gzpe0awup7LThmGvb9VEND9uHtStOSZ5T1
nfPDQPslLuvoKlyV6aQeH93t+5D0Ysz+GsLH09iN2wcLfQf2/TzpcLIHWRw2TopMkBr891sc2dtP
q2sNADTNftNfpl/xc5BqrA4VUvlq122gtyZVjCIpys4z1XQ4IlHddTnaGn3djClZ5WmQ3Dtz+0MR
Pxw+1//M/Tt3JHYcmpd81DjJUckuOj4n//GP4ijJMS/Uj+C9jlMmOzEWU68ItBsktYUqlk4ec9P6
cUhroETGgh4kgiy5kgDz5NXhETVX9PZyJUoRzR8vK77WW6Igk7IlNj9y6zxYwkXtmcFAHfll5aaL
ze6BsnVBfYKpjHHT1TpczSH9fclIhcbfe5u2YKJlQSlA8NjHKAMcq435W0B4Od1WKGOH76+J0qZk
nYaHZ7dwFKjuoFNv2WJWhJfS+hWMgmWrnjf5kv65OYGYpotv8WOHHLN9bCN/nQcnOD5b0AIRhUsV
A6uLQfCzCIBgwlkZ6dcPkVpNFEJBAiGw8u8DELinZArNkSIpdh7Ls8U0RJ6yrOjBj2MVNg4F4Gms
O5n2CQIF5dCikLnlzyxgAE/fC4rqovLZrRZzxf+hGZHWHQCalEux0WVL6kGU7nyOwDBhhmu6iNmY
ZU7dJThBFWAXdgZ4BYeIbSeCowmn+R5Ic3DG+P+LgF65P4uDRN3TA8DgKO5tCLhif/mEjVu/sUMJ
FaC05qVFd5Xb52HdWP0TOQlH0JGDBD48stZ8guyEvYLWN1ay9o38NnzU1471nY3suGJwFB6cRsWG
Z3fGrTXJiOzF9F+TSzMmfnnK2LjuoEx9tb+6OkADB+eM3W435wRuaNndMgEr0n/Xu36i9zbfYVFs
f0GqfvZ0XLaxmaHlBmIO3pekXi/ANI5aFWx5+tH87/5c1LAzxaT895AKDJeSPaAIp2Ofj87Jr59a
18ENgW0lQNboA9yrAcjWxuANCSO36rm8NOYccLIDFa0+3xg9syw8JGMByDSNT5AcRLyIDKKkMn33
TNkj7mnntlrpk1qlM6gjivMpaPSvH2wy103U/sgNZsSHvL0RvCseH6t8R7kHTk7aBLyjk0GsrPnF
+RjFmemTcDdAZb3XLRN4EPWfrjwjVCOb2RAkmC/7Xm0OqzC12wlhot/PDRV8rofSs7pFgLE77nOS
hljG3JH8XzhemiWvN9gMAWJfp6OOtf26Bh5NCzNB9kPHfRUApeZn10buZpEgciC21hdmM0b/eXj4
ExiFND0qfhaHUZHI0JWuoS+k5AXvFcYaPwpm8LAWyiC8xDQTM1yJ74hqHQU9RM02HdZZgnhXYCCH
2cSxYOT1DprmEMnzmcKCATAvx4GliCtJ5k/wKCmw0Df5cveB4naiomYdiAWE2bHzqd8c7g1WCzB6
R51QNz2qzix+tXAuWkKbg5ovUldDeO8CHY1zEM7wifLOqUrm1d9ibDbA6DCUFi7ESpW7W5Ik1h5v
rsUT3lZx3qYnyCQ2HL6hIMNAqEnkXp4W/1SDTC/NahOFzkOyu5nYEnmntPCFJCsWvFJ4i/h0HWDR
x9xZvstFTPaloWoAzNYdM4Y/dc8MlokxC8yLnyBcl1dmxL507eHuzAKL46k4xtqeDBoVvfM3ZjLT
R9fJXxT6kSZHgDTa17c9oOXaAVy+TF2xkGmUloYHfgG2OP0l+e4+Cy1OBD9BWIe94HLfobQ4xeMW
uSOWxAdWaJ8pEjUy78tDQJjqF0gMVR/dY6/IlmB+mPFEu0B1slDkU9gLGFDRWEd2tnjfUXW5tWQE
/k8dbUcDnpHtzxVAo3BiViKSoMQm1ePBfN5jQlM4g6eCh2yXk6NgLYrh6WVwJ4WFS8HO17b8D/TA
ExAU5G/nqdu3qWcGWEfy1SBt7zBsqFR8VI+w3WfB5zCnYlTPQXMLsBVXin5eKbQ24kDqZvEOQGzC
djErc0znTYhpNNuq5Ny1wRdJ8/eLmHhIJeQaGfAoiGfaXsBBEw43XO37l9RxtvhpaNM6sArLzR64
mbxqkqOjr8rUvuLpSxtT3EvPyJtuYmDVUtcrKjdhpKxTVVUug4xJJMr7u9gG9Rt6O6PGNP7m9e0h
VRP4CsrvQTmIboabuPegtfQwLhWq08Ie6DPNc3qGxV4NmpOg92YGO5bhAvM5XjFV35PPAL8yKWz2
u1PTDmjj4tWjiHnPrM/sQqZ5M9f/OLFO3ilaH1fwnFc72dzGOIYELfFB+PHzGpDPfhb2SOgWxuup
gm9FWWxOHjfFMEpF8euKATczT54bLJmUXYIFt21Fzy//ct6+Cfo5jYGX3zJRbIiF0xIZGP1odSus
BkopHtTJtWFsPUNmPZjsv9mGjetDQRvGha0MRqyY1fq5BU6cdPIDzix2zPfRarcrLrtmGsddZf+P
zhzZXeHgpwSI5h5ADshwUYUjEGJoGZJwvI5ejcB5JshxW7vvLd7jc9mtJr7PsxXdqcIjnEHd2I1k
Aau7PrSkYP8pOlVHJLfdP06NgeAdu6xMM9nD04ASXW8JopV07COZm3V5VrRZWwI3V0wXARzsIvCT
m/UhPrwOzKu/4X0WvtOY821se4/rYHwsSFl4nphHPgsTT+7qylJHn+m2HPcKGITPSviJczdxe0J7
rlaq/jwo7SqVwu/5mYxcuPqO9lQ5DbEsCwjewAAHnjWDCE1Zx80c30Lbe7xWIXjs7QDRV21eXOQI
vhldjr7SiLfz8i8JfqIn2KYnrQrVdQvL3eV3hTj5Ll+djQOy1g+v5c1umA1Zq/jWivEbjqg/hZ2s
Uk5+Wx8TSP/zBwxc/RlG9qFgVJsXnhCIEJpE+PD33YhdWh4MMznsxGAnKaXoJUmgdMKMcbrT1vkU
V92gZXMR0lscz2cOP+95TqsOUoKFLbl5MFXVOLeXkqTcwkvuSZZoWKDqOZY2qvMk3e+34YY8r+oa
ifjt2Fcg8VpiwrbxOi64Oma68HXvfFxU/oN9xtiI6mQcTjpEfhcqJeMMPEHlcUWSuzMSsss3I39s
9wpj1ckzc6rllf6bkZXLDPK4xEc1+B1S6VPJLm+xwe5tpS07vr4Ao5UuzZiwxsrWpawfCWXM0Oej
rruBl0WwGgnJvNP9zZctGl5EuufbfwJWF7xMxaqciewu9N+ENQbqwglzuqByyGtdkwA0VhSWnBUS
5DFbTrR4iZj1X3Vri79D4aihjzDFkzlBr8q9yG8UuejZm+bISfdysKy8W+E+1gT/61ApLVfR/mWQ
K5HeLlMXPXKLCsLv+HAJ+qSH5vQwgdHYIV2wqtGmnxAITbLVDrLCdj7jdbygjSlVNHVVUTTIs4V1
g6Wg3uAQ3I0QxgFUewaN3zAPGRAnZFZTXA7L0+YLnHfsxLJU0a5XxjNe83gL2kKmJ4o8u9HfL+EK
hAoTYSsWbOdKZKb/cXxlgSoBQFV2Dfa+tzZn5wzDoimKdkYrawrXou6gvMqqd/5zPn9eFCdJKYPv
5ETb8ckCxX2dZu2q+jSIVcXE2GSG9vhAGmeUdn1gkWmEmWP3nha2aoXQttYy8BsPkhbBWrMDJ3lr
Gi1fKKD/q+M2XNuPseq1jDt5zK20pi+tLlt2+3v8u6EZGpbN/cH5FBYHR49PdpkalqlmHVWkaFlp
Wb2DeMILROrcXGwEHYtopQZtnCiJBR4UMbRA/xbaTNDAPXDMgy+oDVwocWoBXe1l1usfrdbBTElr
JxMpRTaUKXa7dFccWIIsfS0aorPuLFGdS60I1u7t5o/RCuhvORlr7EZITKLPTnr/0s7hGe+rTFme
NjSCPxAWHXopMaJn8sFU/OqldwKZtov4nQm6RdEuJvtF6O/L6gW4k8scylGCYih5jFv6SW1ab+8R
W2NdG3VDtLYPZxvOvZaZBUCWWb7Kz4soSfA5x0VACVyCrtpc7IFLyX2ncWqoTVv15TXYjIfpir3m
Muoeh38/4oxfvk/z2KYj0fJ1oumCnDhdFZl8/ribHIaTTWwEJ3ELnqmInCKKhiYRjFK/uEOlZw2B
ymHO5pq7DsngI1QWN+3zoEzBdjLEQ7kDqVpNXREZzkD7irTfWesDrcTto65revaK4w4SQdnffGpK
D/VAzwvJzUqodYVmDeWsTN66KoSiQ9tZ1ZH72nx1VTBnkxBn9tN2fNtCwy+FVPo5ascvx2QylnnD
Ynoc3dLJ5aW/rmYCWe4ou7uF1Eh3VauyfO5GoRtIoR2ZMxNLuX0d90JaRPu53dW2sGQFBth5LIgE
zlwG95SXXi/hw7DbxyJi0W426n/NuPtJWFVvXuY/v3yfJv55uWFCkvLP+ks2eoLnFg7VyCGoHwGA
qgZ+ZNuS0Wj2w16pKYFx53fTcBChVoG+DHavkfsdYm6vbTtVcKS5CAZXJovR2HQdysGzA7mJ/StE
QDze4EtW3YNBNT0mgm3XcabNh32UODA1l3HCqUYwlxiAsxEvAtgPPjmE2zc9KKWuVd3Eua9bzQ16
Gk5ovaeatwYUz5Gwbke5Q52ZWf4D6b6MhMvTer1+YdEY+4W1MGi5PxfQkxuQlhX+nOB6lk7wWpIc
cCg0zrUwCPJMBK58GHFK/sEThy9nXPsTxtEo7DG8O6cgU1bF9hNAUpecurCBFdAxkbheUnmOXURz
3DNYjonsyDefsYmqiUWKU/rrxUllTuApP8YbTxWmn0jGxVR1tGpGuwFwphIcFjcW9Tei+anfZrmz
xZTwF+tRsygXNq/aPLilrqWxnyLcHKohPsk9GI6DTtnEW4EddOeXcto4qc30JCZE0NIpdF8vqJry
pdTK/tC7JAgk08UftI7xWtBdLxKwgu2pPSs7/NeAgINjH2O0Wxy2iV/RCtcwTDTbg72u6omCYQFQ
m2vYTORTYM5iIctLs9XVTb3G+XngOFEIVO0GjdAhGRs5kn/BRh7Tbdx6nfWbqcnmZbjW7K4pn/pQ
8gPjJOUFuKQQfG7KokT3IckKU1sAOueVM/46My2qX2f3441Ko50aa44MU8oqCvRxQVJVbiyet++e
3Ey4nQ+5MnOuGgoyJ4qwB2QQVQBXbiinTl8K4iK/YsB/2hgXGjclb0ecvDXyLcBHcsPNSMgcxFpR
ckDqvtfzqk5AkLjfmP9kpEmLdZMPKIE86w4GCHlTTxu8g/FpBqC06IbaBzzbcdCwy1yUtwUxQhRb
eMURS4dHXNmHwyponRHaipkQ7pWvg17b+iTWwCqIYrcEexHGELwQfL2th2JTa9Ec2fd1/M+9cNId
LsWE5HkG+eC4TCI5V57E+QTO1Je2Musg8KuEhbSYLg/BmGk8x86ow5gbg2CdDgs2X70/oCv3JnHC
ba8/XUZCQlD71ZAG6PU0TG51YgNWo3UldepadUnMWlL0QbryIX0pFVEpLltYS4NfGwusXohTxMkd
aApQA8rBmt8mnLsI+qnU6UU3b/T0aswa+qQKiS0mqZZhG+lFdSD8NWqeKX74DIE2c1ManVn2CXpj
JXuc03L61Ke+YtUAmO/76RpM+vIJBxqImJYjgLFq2uAxgxLlPD+jbzK4o2OVCTiWkg6yeTOjmzyC
cD3ZD4L4FQTQfsW19jxNxqrtHddky5eg6kAvhrGymnS77CyPLKHW0ckN9b1n3JttV/0mbjENeeS8
8WYshkABD1inRy++etPsWjGa9hQ2ucdGvoe6oNf28caW1dskZwZX1oQIvKfNyTs38CekMklP4h63
oS+nCiBGQgXBMQ+c0OpveB6I/cHzIhEBndi5hQd1QLDqIctf8eF9XJJdK5GyaNkGVTZPj6irf2UR
wE4W5I+l8UtjKzw2wrOb1utB0r1RdwImDOynqp1efJCl3fQFk/gFt7NcLZqeDtgvK30ghVnIFUw0
08JGITchB+BUlyCcgqNB3amhon5nLJH8337MN4n06Ma6yBrJmDFHA14szyayP/fLHNUNnjelVJSW
NHJ6BUc5bHq8TJupSiyC9e2G5bwV8Dfwuey7nFVyTQQyuqRP4zsnV1o8q0UpIJqPVnCd7m+7MmM2
sJtf7PJSKn+UD4zQsg2V2qusQqpEd0ADFKeJCXgvy7XhH0lIh/9eBB1XCJXQSqP4G49K9OToeuzZ
HNTxyuvujXV/6ZfkpvR8CRqYhkYWAQQAC8sxn3Ik+qlAQyQ8FG435FbYcP4ihKAWGSIwQbcc9u4g
kAAjerseO3zN6u9Ia/IPnvLbxt7ni9UMBsgnDMOGRzu+EisfIogZoC5uyCHTAbDTxX0GnXj2vzCx
/O7Y5q6qYkQI1wfO0gJu0MAwdNmmOJ50bGYuUSe5gwuX9xocWEM+NsdfaPPHzlEbFr2ZfV3+2LoV
tx8hNsPLCb5zFp2dAGBDUARhidGhiIsfRcNqQjGJLXwaCQbWbaXlkzqnW9C+v7ZdwIhhFq24ieTS
P+KuUuwNa5xIpKqpf1lzYdQXuIA3+nrW6s36rEz0epvHTExbrt+S90hmX83C4yLNz24aA1iqipJh
Z5azk3+HWs789B6neuceFABdU2UDUXQt9s9r+xqrfTkjboQVkcdfS5hUrgXjF6M6ePchjTWAvUuP
GoSh0CRGfx7AXFto/jWb+8rv4+Th5bEopy6vfzXm8i3xDAPhM9DG9LX9FWXp/AwDQbLdFh5vnMUT
kAPMNjUyGYgl4nFaVDM4GzVSqA2ALNw9GcD4qYymNK19nQVvLPROaSwPfcaFK+hINj9Riqse4ful
JBJ8FPnhEz+8yFrCiC8qibXcLnDUPbDVquS9VLlHv7nH9nL0Cb1dsJ9/LXAw4y+rp/RZnBoUFZdQ
kWOyOkak8We+kc2+BzdkeFwgynlhW08Ygvd1tdN6kJFjuQfeqqx053l8sb3YPTQa77bN7lhuBbi7
FKcEPFZaadnpKOz6xIHeVgTwB3Stlo0AekzHqds6PphcLw9KwItN02Ly/2bV9S472BEFSre/e5i1
4UpyY//5OmNhBr8DfzJVq35sa4xdYR9G/qimwp/dRjAwGOQlzNeegSRhuYu6uEeWnB//IAk1YTJE
IE4hvfksYtOhL0xPrNkKWUrK5N9h814MS1OzymCP8TfMmf9lVkUiWv9Af7oWs7U3ehdhtAOJMXHT
wcpwkXCY7785lDNuQmSu67STgCZJM+au5Y1rgTkDaR1rNNFv01MHv8p79TIPmor7R1iOgvoyv9ej
P/k/RcYozIt29jdb2y1HsI4pT0h1ZyUJnJHl/OZeFwCSTwGFSwzXuyr2lZOUZLQdaepNnOs0kaFL
A+rSQkgarbWzfYIUZSabR3cXgEhiu9k0SGJOmLqISb8mqs+rloXpjTq8k22gXA7XuXXIa0i/Na3e
t9yjFYhYroomerdg3Lsb1uKf70xLvtGD7XslMueTNqUhOlP+H6grDRXZDUwz0mnE8Eo7SEdAQHVb
A8KdpdINSAIWxGnUomjGibv2PMLbq5niR6iOF9+tdMatZfdZJ4WiRTSJpRPfdc6RKLrdmYuClp4T
5ACTQWiv73140tmI5GNIjYejwHRDl2Oo6L+oaV6iod6wjFVQ+7e84sBk4245Wf/k/kVsDLXmzCNI
gl93xZZi55dqG31T/XXf7yxQeGsRNaDcP915Hc75C6iN9kzwh7PX7FwChXD4uBzH/l5VMCZkCIlU
RenWYrmtjByAbOLL6wU7GOo+t/jYsUlbPNUPV10XeVWf4urT3tGdN6q4Zq7LinuEmVFiK0ojgZzA
/+fELOdrTB+occzGKGLXfOvUlMePW8krYF9FveErnFG4y+HspYdZugICz7gimfQsaq/3LP006PIa
5dsOqwZ3kNExNTf4zy6uJMXB8G3GKBndQ+qkkdZpV5DNA+TPY+PTxAX9JA8v1sbmYjEwIlgBzfPF
DpvNWarQvqZuyc5QYItnUM1wc2ugmFa78kLWlm/yFm0b2wHq5+xyX1lzGQukM5+rkyxGVqtTkUif
IVP22g+aEZue2zWilqd8BHxT6MJbb9kChAVfaFPBal42jq1isnGOnwqScEnJctQQ8tTZXv1kmOK9
QSZNMlUnxGJ9TZUxPyhDIhht/y9uP7JqltiGbxvLRsnow4LgcwhxyE0yv4tUZYKueVPODTUL5Sm/
y7a0Q2WiruQxoFo+F2wn8Uk97UbTR5yDWIInM0IkUNJ1Nbt0UpmIQbCpOYFzKQmp8snDwA8gqMij
UFmI67u6hrU44Igm5y0WF8pIWP+uAdptvPCdlaYo+SAlTU+4Rrue+rNQPCSnHpWR0Js2Q5xlc7p9
SogjGtuL/XlyuMVSuaV3PUPrA8waIVaC1T3VI82MRIWfy0t9UDhhPijZ8PSK4kI+YByUxpaoBG8c
IBLzYhOHe7rwW/QRE2FOOHI1kiks47ykNYFHh45M+CYd6NqE721SWD3Zx+v+lk8Dijms5ncpdH+d
kPhRR+QVARlQG54RzKCV21dxSH8KkWYoEcsn1Urga+9NrIzIxQki+IbyIkp5eF3bZP73Bb/lmk4K
wOurQc1MT2KNxeRYHM1X5S3NAWDmISGU3BMCLIJNbBMG3TUs6n385i97quYajZ7m3Q/pKE7Fm7dX
Y15CRcddkIR+B6LPTp/A6H3DbwwPjxctApfXaGAw59aL3MIZVs/UIh0eso7q1NBa5D8WOOBukqG6
mBfL9CWSmKp9QWXs9BFkaJHTFZKbiZxZNISYa18ccX1M4tUPgYot+9VXpaZ8042TJ4UsWwmR5GSR
Rpx8cbAgfUagVBXOq+gA0tiMUBAr4WmU0nm4Rvlikcqa1EYZxz+BoWBKWs6u5ESeXhIwP9/Ws0rY
VEO2bwiCEMSnqRdxp+g98fZZ/DchkTIDaS+vXTwR+9Rii19rX+JuS/l8ZGbh3dGw8/CnFivISAy+
XbO1uibeHkyS34MBRILZL/RAjzvYIAFxFZ1dWQ9eRu7m8w8JQypSc/MD6Squ/C613ZHS+F9R3atJ
8IAIUF7d1gwcwo60P1GlMAB885X46uwp9OXzYPBS7GCUiE3cSYWblhZ4ojYjRVYrmSR0i3pZuAnh
6MYAoNnczv4VciMsHjLK7m4cjeP7pxyP4PJlfQjNBIrxZf141OxoIyIE4ze5Vh0vhKUiDazGAFe/
lE9MDOoAPBWphutZqppTGjDdvWfVgBdwMOi4BGqplggxCp3/SkKmmdidJpO0fpVuI8MEmaenefCo
Lsbz1rCmA66ZwVAJYyhFum0hOT/qwrSRP7dDqz76zAoDGjVTHmVxw/85CjCOkU5zD6iWJeFG+09z
Ubxfy0S4RWOW3GK4tWRF+4InjeCEfrFWiZ7mPqXYGMZH0rnkxVD6SgD/IjJqNaKSyS5sPvP5kvy0
JR4VKLdMcpgqOmr6ah9tmKSD5Z8+pO43GAXOlOa/VJpKvThwzbfCEikM7JtvuWXggxrhXhnCMY+l
nB3eTWIi0tjf5nhcfyigh+1h4R2m9ZY0fb3I33U5MKP86kvw6kgQANXMUqFGhyNG8E6Vjkh/egtR
NhkHi2H/UY5nqZT/2/NAFaAGBdEneKVEVY+mjUL2q2+7oaOIhO07B95hAOHPhGfCn5a0F1vKE+dI
fgM+xAOdicKColKcd1kBw0K+Lon3BAfHjGm8rUGv51d+zvCvrb+HbjyNzfSQktDqKKbkcV7d4sr9
XSa+6guGhQa5WddUrZCHTLIRfhNY4POMzyPqOpLRCKenRk4jPxGCgtyDef5gSUe7keHaV7Vb0jhB
JGXkW/OSnyvPcXx+7bdP28zOYOwBQ67QF9kdJzz4S8c+a3WaRjgI0V5UVMbeW16OFrf1kIVSuO7n
tRuumoiV7m2gxio7KAA3xtNjDThGgiKyQQdbbvqoJsuHIVM2RK3Oae3UUP68NNjo4Wqryt/lVhgE
wkw8RqA6+uTTP6luiFVQe2nCZ7pnGcXijJbCcfoxMNsx1/QLzmqJQsdCKlYAlTQeR2kmpRMHthLg
J38LAIVkBrZhtiipMFdZS2jl7X8mrliQNdOhG1akQV7RpPvdiRe4jQoovywoc1Z3OM9ecPgS1+ID
daUnUf9S+MZQ56SefC5hzGZdBX0FWqp5Hw+7Nu3O5mEHcSX01JWfbO89hTa7o/0CmEZAnzsR42WY
ub6t3Ysh2N6UzWHT4tujlDUwIfiLHRZKsW8WGKB4EXI424R7Na70TWJlEKG/KhhWWtB3vo4ZQm4d
7f3OwhUhvGOMwvA6CKZIB85X6YdQhzLQmoRZWXOz0AUUi/3Ece0PN1zgeqjgWoTGoNUmrlvXeKUq
M0wla76bIiMjC2SwDU/MVu9yupcMYBPq8nzscm0SbFHPihZ7pl3xUjoHUvC9KZH7u09qQNi+JujS
MfBJ8x5TZqLJSIBi1bD3e5AC6XwXqMfM9b0CBqDpnhaFN+1chZYnbBmahlW/MNAqGd7CapjSqvB3
MYWn8uRrs4TAfigtvJWZ8o6HONGtI99/B89BbAFhuFTqpG8btkY0dBMM9A06mM7JzArJYcYLMIuO
VJkdD5taTmdCDykW2EePzDZZ5ACXrC3tgw2jtIl6+yTEfOHgBD61geGn6XGSq8aE/eSpSa6usGfV
XWcgTuw7BzGb7gLZlgAUMxI62y/meOuH8+43LsIdxQLdjKNqEfZQpZzMNBNWgUt1X2LpSObE17Z9
YFBVJavA+LTT2NFPOhA2IOPaYoweB/vHip+2RMlGAFZY8HwNWCPPu6PdT1ezg5AlFFQ3YZQ8Voc3
u2qZPk23aIhbo9MAteWbAAcx46+IIp5FNdTzlmGernk9w3Tz/uzKifSLVCXVKs9l1VTUNLjSflY7
HeoYos8DNb1zmfSyew+ItHZkSfSZdDCZY0J3bLoMpvHfW0NJ65foFvAsgVyWNBap+R/FuZcj4dPy
eaYN8+1wkTuupqn7gCyIMNzdmVxQcwtiF4rmMEvtbtw7757daXEIO+Zu9MnsIH3YI33gUvNRcMbc
D6rp3ln30Z+N+6onRNqj2726RxR/Tf3SY6ABJHeh5A4JDgS7Y58MxXnnpWXpcLoh6l4wR4UL3bnV
n1usZM56x3QdfK+5wdK+7PzXrsD1MOiBolBn6JZsWF6Mi3OSbTWKJM9UOSJNYnrYJ41at/Jjre3x
wVqexi4bnnJqwSq2HSwGpykIyTXu+vwVSJWLRr/O1IX3/vIz6qkoVAe6g9/Zg9P4mbUsnBTWQCCt
i8ta9Vn5EAGyzIcVzjebH/c86HCUraK5tn7/590MLRNYUgt91RDZ+UJK/B5gCIsuiRV7hXKxzfmd
XULbPGXLGGGsLA/WmI5fnmrCwl7Ia62MO9KKSALaFW3MfRflMkIZRCvTCZFSREeS+dmIcZXCqzYg
fsuTW44P9rhka6ErjMMAH1zWDyo+Sj+bKcwHgI8ouaewmk7DshkgPcKCwGnm4zly2bJ8eMny9yaY
X+L32JEjXm/7gXjDGCpua4OXJn0Yha+xOhWRRoQ+LdRcRy8/8jEGiXSsG5cG361h2jkgNOhM0BMU
jNWeArv0FN4+2ELFcIx5mL00DQbiWVYuLtosFu69C2KDbarNd1GDWGrYTxxZMpMHbY7LOLihJx9W
5rBEUo4gJtMk8Blig17Ay+ipClrKRT0c85CgO6OoT4I+fnilSNYyuGuZxWURiiEwGDIwZLWDVCP+
kSHuplw6jm475VP2xr5Eh79givCjuyfG39opKDa2095rCtuluSBvP8mdl5SfGmfHi2dboX7XIjft
R3PDTwliIXaLZGIcp/fG1mmL/ZQ86/NTMLLUqKqh3ljN9OcPHJwWlJrmn5w9PsRqHwE+S/GRXnYG
vK5p8iwk1gKmUqEcOTTj4Vwl8ckIh/u5BBgTCxRl/M1M7SgSSBpTsp+JRAb7U+gKu+6dt5Js1vYA
pN4qRSxeRSx41gO24SjFnx20P5Gvvz2RwFNgS6QFJPEJzzpdnf6M6rhC13cl5YbcNGsdJvVwgg/L
q2xiPDW+w0d3euhih6/LjxS5Ckg0LoJemzVKCX8kZ9CghjwSgbGdX5VosdiTzVTEDQfNGbzlRJtm
0K+8zV0FDAdNAxR1WdrkLBe+f8PNk2PfmRggC32M2dddLG9hxkhg22B0zBm7G6q9H60ZlLeXSfIb
booh+SQpHywOyQ6ZVEEKUdm3oTLzJ7F6GbI7UrvZ+JjmLAAndq+fn3DG2oblHDj5exVngSsHKreJ
HPFHDIw4QF3qnH1vereaYqa4d2HLINHW/Wa/6U4CgRczoCG0JIgCTomFmW8VuMftUB4arsTveCjy
dUXIRyM+bK6UKFW0wlkln63I6rBaUORq/lh+rtfudiv4K8GZmZ3mRQ0moxHJ6/j5Xa81uql1APpj
zbGPApxu2Ucw2Zcd9/YmorOdeAp4bobQ6l/HC5lvj/eW28TzRucgiHd4IK2x2NTEXuKvf+PdOO9y
RTGq89toAoxy1Fm/EwHBOzw+Vl0iTuGOLca7kf32RRHJIMWOGBq3h3c7dS0CAHdV+KbUAWh5LAtq
xbmCHw7MTT9VeLM1ps6MK1Cz2qr5Nez6VUATlPALQ0+8uhWdE0EciEcfCi6kjo6dC6ZclKsoHruz
p8Fbtyu7/SN7h5stcJnTPUkOVOQ7ojwfgQuN6sQ1q3oaFqokhFEA61ZSeY85FAwbdGEWNA7g81uU
MC7JvZdAl0ToA5sEBgPV42vCWwNFTt5ZowCOIvgYGEMeSWTeoIwjwmmCFkKuUVwz/pnQLhK1pPZX
vYfRkM5+SO2/5nJbFEk4yhOnoajZNsDp7m+IpgFm24H1uZT1s0d4/UXK023P8IYt/xizsE6MHnzU
RBB+qOfm9esAhNycTeMQmv/HBmqSLoECsivB2IvTTG5W+0DRZOrw7K/MYQgMd10MmFfdJhTlC3/c
IwuIy1HNIY8OhANZ16ZZOA7jwCW+1kK21TORMq7f93JdzKCf65aQoCWC88GSIfN4i8wCeaF9J3oz
KyMbTucoKbJ4V52Qs6X35jddQzRp1UjNVX4xnXkb0/0meKjCq9/M0SGUktV6SkubkJkeraJoESay
+7yJkNhVqYV7EzJ2d3GyrnvpGhjIvABO4zdBtfRh0vc+OrxzltLWMhQSdXqrGVp9/pk2afPX+Cba
ePYPD0Olq33zeyhe5P6fzrMbsxVKvMsSi0+YqF+7YF8xT/E0TAteChTHnRkg4UR7Oi8Hc0mKGdZS
wxr70Mjzvfqv45p9+KJQQCzhrVsr9C3ocp37Uje4fZucxr6xunFQa9sl4SV+Vu46puFgYvcEoORz
96nX04IzZGlVUmlNOG2gPQj9L3Eosc7NllTRD+i4KOymoWR2afKVZJCgN4tupsbvL8Ea8kLAwF4h
nA3zmPXZiSnQL8Z7izbYpUPBXG5NxTihdaDAFL2SsCNVtrd4hyhLsCNRKXhMMG+S9xZXVoDKGFVV
fwISLgIxs/ZvDxh5GLqS80sATXGOn1BwEkxecVn3gu3s3pcEur5oG1ZYhp2hLRF5QjGPx6nt6akG
FrnFOxnA4WaA/8GmOV/EOuDOskQimBER7i4C8kRfvWqVTrzo336n7nfd11uOLyUPsFaLRLY25het
8jlOGnlBXwb7Ne+Sq88i41Dul1PmivsKl6O52R8X3wa/oxDrFL5mO6ed/CB1knEywXsJi1lyyH+9
L/+PY2FxCpIiOLTK3hXYu7AY8+dKkRItsTkETlvcpt+UvnVzJ9lOB72l78nVASgNzpEVSPKJAsdU
6tujWYlcchPPOPquCgMKwhvq19/gSF5oXSp/7JPttDYAmVZyFifKCBMLC30cgy2T5uSzBJN+HSxs
YTw6Ax8lL3F3I/Zx95obOCXKReOCY1bxg5PskW0RubuZWx7Fw2RrenBBzxpF231JjNZrAObEK63Y
EPBUaObcqAhdRki/NWaIoUKeqxl2XpNywONp5uXYA4r65mbsLMSO5bWSmkAPnFlkW9UCkhX+9Hqg
lPPAVD73cWmPwhmwKg5FHyYgIt49HPtrcoiicIHDHpSzLph+WMzvCUeKAICvkhuxKo6sKrqXyArk
MUcvcTucGOD6PUdtnAQheHl8ud8sTGtifFUWBKZnRXuDdxCvi57BsPgyqb4kU52nPwfBOa10AEXV
5YIuDda0DL8E+hKZ6wPnymwbfEgMsVlUXajpjCgdXcAKKlr3aO+6dj1F3VR+hAQwZQDYl9hZc2No
+OFU9XUKZAbMwyGl4rRl8dq6C0v6YesuC+5xvk8BuK6MHUtPcp+Divbfcz3J0eVHSYZA4AkD8JvK
qDx8jSxzStw66Wzo2Dj8C+HSQFiXL0VMd2mEv4qwGzlYCyHIdzsIWYv7sQWjcXUi1aya4KLX3+Cq
9a98WFGvZS/UMT8on0lsk2xjX+THBWo35L0TzhsDZXQv19ZpkztyEOEgYQj4EmwlxjJS7akQkFFk
WvDQJw5NRM9fuZoNm6WV4zZHxVAj86CAqBn4EEU3aDCZY+n2ETKL08xQRuEK2hKWe6ZDutktV4p1
CF2CL8lWf6vjC5YybagZX4JeF833K3+7aK1hRPD35YzCLr/CHQGtJ+Q7UdYEdU3vB9rPM5aPYQyf
Gt0rrWiXuZiklkl/D0eCWmXqvF7c1jAI/61W7a+CvJjEL0mrb4dPRlRnjSY6crva4oKNlTcHRq7V
fgTzsVvUGgycIgW0x3kyjNMb9P0En9Bd20zxOBKB/39mjYhCqklDqaJ0hxTt8x+iZkoTAMIlbqoP
LUonbYBXI3GsU/kSJCWY12FHFoMdRWnesv32IlIKSBEuwQyEQcgrEuFYXVIyvwN6AjgkqIUEUmRh
T7WZzIlW30Yd/iVnToTbj3ZAq8iI7zzQjsDu71rmKcPu2Y5Vxzzg1vDtZP2FC/7mY9Ne7sTSGTtQ
RYJevWbiOm6d7X3sKk/CxfAZCMWPwZF4O2Uvu+6gioFKrPV2jWGG4Ct/nV31cq2dr397ME5xrFOB
NyfKzE8VPqRGrQfbeDIMCwQKjxtAOvcZgGYwxOaYogy9Tyqvfie4colmCLjn/eldWSX2FABtZnmN
Bh2ewLLnKCjw8ubaEjCEKhbfo75DaXDcIup4gTj/HUzMBtW1iNpgnTGeXFzkjfA9VoIUSTx1ETkA
AjhZAn9E8N3witlaJmyd00cji7RJz80c60N3OwUZff3o856ktVx1fjs9Ktfcr6RxMq1EeCR+Q+BZ
ypQFIbf3bnz23JLtsOWLoFKPVqSpvZf5g5v9vTD0yH8u0/gr33N98wgh2i/2gS5HmM488f4/yz4Y
1mQKpeQToZpRSjrHLqDxpop0+yK7FDKNlcQPjXeMkfus2nmH1j19al85DFeOb2XNGJe4LFZxgVGQ
d3128/Ow0XkQnLkHCfHXnGOcphRe2R+/cQnEx2QEqdYhCHbBsswtwAwj8freH6Y7w5yWjrR8TdNA
oYcjcJErm4GrFBPZTOI8Rl2/MJHstkktv9JUXM/Wvo/j+kd9Mn1QM9Z5Im/SIC8MoZS9J/7JqWij
InxyB6r7LLGCrRUVbtGTEoA5xi1DMlY/om3GVjg++jS+0QFvt5c78AyTRXBPvGo4Z+6rkQhWrndT
0UopqcYO3dpWliuXWV0GJzCv7L1j2abWiKZy81yV/D9e6lOShk1JYMnvHA2YJnRmJiSCm/Uro9W2
aSE2qz1IUumikN/RjhYFtEMIMq2stUj/0y2640S+/WdqRn8sP814Zfd9GYVh6GB15RBhUoAWADi/
sqiipCMBi18Y8Y+0nrb2DvqMWvrReAlNdazHC2kN+Z32tV6LQ3K/KR0d+kzjnwGQu9gdYMmCezQs
zZsL8oA9WvxqY65wpfYrugLqQ79Ed9xrroZyS3iTMwA3tIeEkP3dcCj/9JGfRKfpdQUOsMVHUZ1y
/l+a7J+IX0zkMAzbPYm2RyEzDJEGeVAUxpst+TmxwC1bLPDUOFGwa7u2c1Qs3yZxfMI4A1VDNRtx
I2UsVK3oSIMkp/j7sP82+8Fblmn9TENlh3IPNcngsrjwXp3lpjh7wckybBBNwDGpvB7axvxhP5iI
/YXcB5JkdjsdwCdYzDxRpGjU8IZl133DK3Q4eTql5m/YDfLhTTFpdil4xwldebAwumoG1z0wlJ30
vC3b/l2X2kd3GjSB3MiQOvrXmW+11U9Y0ermrUyn6X4kcv4f3nFjie4Cjt9OnD8xtJJGN6pxllMC
MZZP1NXP02WvA3fapR67zC6CkK70Xj+l2Fbg4VSngilWrj1RZ+9j6LqIyosmGsGCr+QVjcumjCfy
TyiVjxpA6nFvTZxfjbSYBzr253qZNn+NyHHpiOHPQxQprT8lvwRJc53LSn99J28Uu7a5ZYZTti7A
FlwMNdZgQAqOQlih8in2kitG4uaW7riz0yozDTj3D5ipI5zRpsniKyp2Te58YWjfVfSBwonu2ZNy
VxiW6lQEVLbjGXQPx5qYMH00fJH5xaAfiToDkFh2RRv2PpV1xUt2rpKRaNp9z81IAdMPWgiB/Vjm
Ror+AWT7ciIvdW1Xz1MP8wAO72NA2A2SeuMl2wZo08jiHYxL9pfJHcE3S+91yHp96330AdGe2xK7
+8f49of0BQj2gqBiZj+MDYcQI93qKcCc6+o4UUy2JxhBi61jEzY7Ytw0smTJ9yqkvgCSHyl5QuGX
oZ8lkR4C2uBKAusZUlSAmvtKck8kXlfZ/2ejaOUo/DG0jngABy4yl7Po0javQZDubFFF2vioYjRW
VsbPItiNDthvgDc3LBvS+gjQgM0fXqETKbeJtUAx3lM9UHaTDlKGRUfaxNAjx+E2lDV5ShlhRrzI
C1kRu7x93Jn1QgvNy+iNlXi+4OMaba+3K1RgNRflaRvuVWaxbkQ4zh8TMS11LyIS5OT6UXDa5xJp
/cdLOHPb8dECIvserUjdbsk5hY5hbREC+PFIMJpPRj82+KgDHilmpdMKpQkJESByyPN7G386Fe6e
1O7u2aO21JF2qT5TOx0j8DbbQWmBPBb6dqkalVT4Yei+KcJ24wYQNk9v2rw2RBLa9zJH0UOObqIU
gNVA6mToXucSj/MscEyIpOCrF3m13QYwwUIZWKaqhfeYO56zvayYCjSMTAdyuIKdWZF+qJYBF0gM
NeYWVL6wtiUcjF9J96FvMc30bQ3UuMAMUvv25wTE7nQCHEwj9knVFG9GBepLr4uTbPeJcEA9xQH3
lEo+FO51aKN2pBjiat1YmRtFzNm2tj5kSd95vRRc6coyw++/4ydacObmhMj3sPfv091ggtZYzPMu
aUaHKpetxWlEVOYVaSDtKnuyCIlR1Aycw6qZpm9XcSDUe9I3y0eLbmtqMS0DAlgb0fdhAJHm16o9
j3Mcn0A2dwEc/QwwGdE9oyzMkcMYPCKjL1TXo07mTLe5ZPY63JaVz6IdUfrPOwFR9hRYl/6uCnAB
2WXXpEMToE2xCbLGOSNSQT8eW2xLmENORxHtZXYESO+7DRJq/hO7KegtJrbzatjL0StAD9V4++Vo
3W0hvtXEYHvnG9/z2LLEFFZ+VMQ/V8NDCmri68kNoHvGSVwVVHJxIk3jrULBuzr0hrmM4q57KJz/
FcY8u4+yz+AkTFAqivnKg65qaLWtMSZfl9w80zSIlSZlJHVDB5dBHxIm51ef8vTUK92n0N5jrpNS
kImHCv5RXexplxDMM0SpRT6rIahTi4CBnQaY5NbHz6MEAex3JZr1qiBJXPfZCiwP0lkn8pMxO6pN
/o1Xysmm+qr+duV47S/DiG9Yg+MQWvJQhTeydGGsQPRWYSBvfrkhdHNbZsuTtX/HBuiD96skiCt1
jLsKo7H7ARqTCTTqmLs5Aeelnw8YSFFmzk/HCzHD2Iqq3/FCnfnPNmf6euRPB/fGxx6GXS2XGuxJ
0bBTPQ0LxVEPEz8DynhphQ1zSiejlPCIDnxqf/Qmsq5tq8TmgC42wqL1fOSizhLcoyrPXZPPkQ6M
FakaJ9Sa3ERwY9YqGZ7lRxcV8rNZfEuRt8vUaiS7QMEV4hjckAI750C+gUuNJZSaVXHHUfaq2Gh1
sAki/E50GVPlcPL2UA+T//uouZR9GKXvvlY1Zgf/6gPZeX5yfuyoFiD1QhI61UE4m7Uzx2p9We4d
5MFCpp2h+1dN8CDwgVO73vDYuWNlsJoiwLamnBJBvpNn9yyHBpCkklMMfYDEgJmpzUJXG8U3MyZ2
57IVKdP8UhJe+RQuzV5MlXWAxxbHomQ1cja9uTysib6mx6KU+4ILYJe/a4aQFGn1sPntbuMorN5j
q7yF6JRw9mvYgmOIIoOiP9THARSPPhZUi0dTK7bqff3ILhc3rUcq+fMM15Q6n+uRvHPhpzqcCKsV
026UXAe1z97FZBuTVjDr/7fa/9L3seZXuUz85DDj54N8zJt5IOKkkoDoc9wCpUTHEJu0b+D8kPbb
1RkVzephrNoKnm90gHcQR+ZVD6Tjms2BSwb0Eb6bnsOIqusdYJQzlTq9HG9P5Jl8p9r9IUyZgvC9
2NimXa+LFrLYAGObuh3R32KlK+RPI3i+7VN+Gf4IVcMcCE6jvgduaB7XqCpjqnKAFpdrKz80/QYR
SE3xXwCAIgakBjnluasVA4q64lEeY4Jixwt9O8cCveczvgPcL6cvSDy8RYFz0yjQz1FkqYiCae1S
YE16jmYa828FzVYk+H9iKq+yWulZCHZgmjX0D09cLbcTsVZ4dU6DxpHmqnZKVVGtIX+Mwpw67MR8
StYz13cIG1aD9Q2g8T8J0bv0NEHDB3IfhbLp2gHAag6u4k5Vf5Hec+6ElHON2k3oJE/jr2VaTByI
GrBh6IQGFwpvV2q07IXJpLoQcQNaAaK0Ux3Qon/j9FtjbnwS8KGYWQJ71jD7it+vl+Z9tqfDlGQU
LrTcTYoZ2VYkzav/x5l+BzbMzpcDRFlEt9h5Ed9GakbUxLoiHVHDgkt8dHgjQX/T5DMVntZBCDJZ
JZvQdLUnNdzvl6utKXlg8TTf6wzPWCkuJieXruG9j3jCJlwyuDgMYZT6zReoZ+TA6fyTGywdnBpM
YLYBZaGkY+/vd2opsjq9sw7rywXjTR2/qr2AkohQDDc8y1i0LirID0BXeqXRKd+NMOltNCBYQ24r
fu1ER9kXcTOU7F7KQuNthvQtYAmqyaxmfXUwMQTECy6WEMk1kVHeA3RcKCRghx7EdMgrRuZQk0lR
H+D9Zam7QDT66aLt8lwXrVbKSVubQK8Zpu1GAJimSsST0FoY9buxIhVKqaHt6gbyu2P4/33M/QI0
MuRnWM5plkVni1r5+zP9i53UlYbqdmdRPQKsbzDSvx6UhttZ0lA+Vj2FUDmd+7M+m5jExKn0RAap
z0fvLbgDwya328aHBs+bmM5vP/j466Bs5Q2jvCun4gaIxip5WNMvfw+edAuh+rKE7JKvjILHj2bC
0XOUCDQSp79hfUwnDZxAcetsmqeCLgdz2pc8TqXN0TM9MhpYrXd2jcQG1C4tZUx13Uvsc3LHwta5
3ulsqV3SAPYhJ38Y7NuWz9iZlII53vocGUABR3yJrcXLURi7k22R6wp8n9Ya/QKalQA3l1h2X11h
WvnvLzFejmNjwbGUrz3ILjmIFHOP3UFDC5YojTXqD7NMBMvvokvFsFdipEUchC8nErlpi5mLMDfL
W6FwdVv8mQf9md1kjErFXAPaKoENBTUb7KFq4KSOMCxz4R1lWACyX4p2B8XxL94QQuB78eiY8hgf
//hORrrSGeIByKEojfYmfU14cOoMx/AAPY57NviP+uPhNauXhnphK98dXnSqWfHFP1lEEFVQq9AK
dFZB6NLowA9kvCNVUYir3ABpJe1fWCO9YVudKRj1PJmmoNF2iczCjWfLGCXSpsz6Z4Q2QaDuzFa5
HffaIUs96xIvaHTo51nuK8qGziCLSKCcakdbBA3e4ZbMM3NiN0hMuDh2xuXrxRr6irHjDproOefT
DR/7hO9XaaN1nVz7zlJiY5XLxVMFnNffziK1Ng2cJ0RF1n8X5QE8/d9yBecD4+s5X9+8i3ouDwHE
JL4lh3wW2xxbr9cZcwNxkA7n73H7OfY6/4R+5AVCYWc2ZoRm+09iHIXpo+NKmIjjpVEjMX2yyJR+
fzSVdektym0Nx26Id5Xs0FvxRIjaNSj53WybnPA7uLOrcShizsftpDlMbgKXPoiFS5wWIrfEL3rX
vIBezMHhvIBbT/UUWEB0ws53Df2a++XiKA+lMr2ocMz0lD7Gl2BKYUfdPzTrgNUC7Z6YnQscWrEn
KSvOQI3Y4PxJXFlxYAd4h4j6z/6Pzmgb8pt3OffUNAEC/eOx6GXjyTZQ70c3S3bdXXBmS/FaT8x6
ujKl69sQlvN3ZStFrSIrfp5kWrOMou2j4hd/NnWPGqX66EDCARVobRfYwmXdDbQ+DrHHQSfGKAhv
9NOYQEnOiNB9uPoTaSnhXSGiOHAbMN9BRq+OIl1LrvJZhaJRv7zEqlr7PPXMAlVknPnLTpreB2hv
UL9+4ig0dFC0HP/M63dk0zQD/G0L1jIDuDmIyXUiIJmZUAK1q/TUHzp2XGn23uKx7jN8TiHV9xbW
abxCz4FcIEN0vm1CUWQH2HnVOT9n0c2/KbaC1Zb04JYG0NcreJzDhO8Ha8MYBRQ9UM7IP2bpge/E
OAQZhel5phIjaDcus7yQNWgxBTdWjkCqHLBqRIuifzxFi1hXSN4UtoJ+evDoeNogwjrBZDrkfqXw
TW12yA1XXC1UJ6KcqVGiIfb150YMuZTYmc2fpTdqerac5aaBeDLURByz533S+r7JLJzCr+seNzje
5AXzpznX6S55gJpF/pYr0qG5eteI4U5XQYaFCcov1O6NnOF8uUIleqso3dPoauj+PfHlOxj7KA8Z
Ymv91YOxS3wK7DEmVYK2lxSmxuqoHv9bAt/J3/FSRwBOw4/xZT348zfvTBEgzfoJF2l/fTTaLb0D
A88Le5kNDqzR3unRV4gKtwbTqw/aZilalC0TDDIzIXJAdaVtTnfvTx62E5/E5b5HTH/zKXQ7lSvI
SK44rKgXe1hAE7sqajM9UB/pCTdAzvn2Qu2lCTLz3sTlIFAvLOu7N7Bk4Zb3QbqNBpjUY+Y6EBjI
COOfKsaNrZWup/vBRS0xx/SGBfgxcxbGExyhs1vWcRCLvK4hVUvEIr7Ja01V8qtw/0pvbuBi+CwM
2cHrXTPLPJquqqA9KkRn0jON9c+FtPKsxanV+IrpQWtRYZrFvGrOo6dvatKGO0xFjctVBW7vBeum
B+Zt1b8+uMQ8NYJvc914q6xM96W9pYoxGMD2TYD511V0Us8f9yRbekAYTPeo/QAwhHN7/pONCWCf
Qel4mWkDSvZYHnHKk0JTIpBE1FU9uAIRvuDJY3fyW6QRcjMCXuHUjUbhSRgMAUw1lvChalVl+YSG
9V4nHN0KRNrEgkoR6dN9wkjQOwJVricz1wJ+KCR+8o71DP313WwWx/ORwn6YFdYMqtuJKjmHDlFd
p9Wkm8AOdfoUAZ1lxxOnPPE+8QDCgmQp7KdYFxLCmLi5JSVqd0+2S/0MRTflO8z3fhkEP/Thy78P
bXzNkCKcgbVTE0643ywaw81xQ6Ap68FvGSym2Lmb6lARErTc2WunXfTYyGG8j6n0P1ZqiaLdoCR3
eCQ+gqSqw5XVq/t+trAQZTR2asrj8rwJ53vqbiq3juZS5cW9Z6pEZoU4tISirqTF9rTh1zmIwSCS
txtr0SLr8Tc+v3aBexCgRY1SQfW+SkZuLd5ZzvRFwky40C1pWwwQ7xEo3ukAxZH0YbzPEvgpREEJ
rULEBgnlYSMq6aWY+fwj6tRmpMj7W1wAyXKvURZOtHLHgG3dV3GiqinHYZfXH/Xvm4FJKxPyKpzH
q6PLvX+1BGgFWq6IU83GC/QGa2xRhgYs/XDKpTnfpQQv7sNinvO0XeabvFD+d5MTyUY4/A63qavx
V80jqvpNaHB3+AZpfNMnpVWhAtqmXp6w4QK2l1WuKC0kRMLOvTbcIy5wbQjEreWwOLMXXMqspuz1
9CLhp3U9krp14X9NbPwuZ231t6w23uGsUEEjLON/PxJSCsWDc6eqCWL+p1Q8sNrG2Z2azSFSMPjD
e5E66b2m8J9UiMRU0XLbbj7cch6Gtcz2KDB71cAK9u1QXlM7no5SNIsL9HY8FEDsKKC7K5WoKdqy
RrQ1adh3CWLgHVtsT71PsbJIoHSjHFD/4/IsA3YIJo3uReOHt/E3EgOSTq+nqlxvokMElfG98QIq
AhOjQwDvFURUIsa+Skgp3EdGzpiUGsXSI+vYcMTjK3NnnfIfHhj99AlyCJT1nh4wj91fZXP/BbwY
P/OLf6Cz1g3cXEu1gDA/DDHNRWUABdQXgMe2rJi+CUAgC63g3D04kW6rEBlrzpXl4ILKF8eWmOCf
2PxdDVtMGcjiOkhkMaaWGDDfkfFMNEP3Dsl9iaLZqu81VuCRl32VzEyT09BB+6VAAXbzycWe8tI3
2E+Mc+tCItc0nhdlz4RATvoeAe6bT+dsxR4L/FRpdor/y8o+92Gciols/tZZhDIXakVvxBYtUT44
YnUgySkGerxhph+JbbcPqz/j/6pN1ACSRZJUpaQj6GKMs+1SOWhHXPyv+AaBrXbPpFceeqqUDn1Z
ZGEHXjasSUBEsugg3VRMqsPxjMq3F9D7kukPcowO2FUVWErCuOmkh/F4BQwHUNEsbmChW4VjH0OM
+SGy4H6fUuHI/Xb2374Iaha9l6FUWxQFnZUP88v8S8pAQVjT5ZgBEIqkYTq/q4wXn4ZF2UxsPgxe
kYaL3jP3eKwWTkz6OpILS/Qnu2fea4hHc0lYIjeFaDQojwzmLSo0za53Qq57sG8zCByMnjNi2GtD
glXsexo+aLR+56wF6VrwNnkZ3Qtayv2zbDPZ6c7huCQuLJLr2JNdeuyJYizgU/632AEB9h/X43RP
bbCJH9AbeL7rcC62et/N2gxKeDcZhpnPLytLXPfLMCTneR1/ZNZ6TnbOhD9aYBEkUf+uBpO4VomO
JAkzeCe1cI0cMobfOr02PY2at1titBynwCQvFhfk7TZIgI8Qr0yw3t7L7QDhYp2zNP6NTfYc1epW
JexsjcV10zZIzKUqKjS2G+w03sC70vg6ErdZAd10jg/i01TTxRWsYTFz3pqsFfdCTsvkHO09+HiV
aqUGOIRsAYcVSo+Pf1tShWnsnnngditmLVreMdcxdGtLQetAQeZk+1v1vU9Ai4aYxU16AywFUmGH
/mUVMzZknOXMeZFaG6N9Y03W1/rWOGl/QbqaQMMNEdf7naEyuHj8cDW5OSJt7ArL2SE+her6yu/W
WT8xr6orH5HA2/+DJ8GqsLuHS7UZq7thzJkf/GNNI6Zjzkj7MJyPUyc50t9qYrCDfmZ10b5KZgdc
DE7tZ/iMXBEf+1Ri19R0MN0x+eFjE7Fp9cEyUha7KviU/D5XUa5qd9nS0/3wX/3Yi0T9ABWa0kDv
/LORzsvIYMssH4qyt+bLcYVyhyWYFIN45wLap8uFlc+smL/o/7fXhrmEL7irwdNEPpD+OwWxJtGl
WaTW4C8DeUiraEllrbqqeVbEanUtxIhPNG7gIuCqVNfY5mUTfFPImwiadax4gZZyiKwFcUs7feuB
XrdQhoahNPUsLSlB4fOCuV/31FkX2uWlQ0CNiT59WA3NbsJY35rWeFoCldwwtV3m2HLvD6+UMADK
6FQ/sRfoQQc1PHOAYcnkZwG9msNSx51Un8RdtlVk8k9WesqeXmP4VJz50kMLx/6/1Eu9O2cY4AXX
oPXsvkp9QCDsbmuFZXW3ye4DkUBoZpKhoEPDZjtooluSMQmH/EkzgfT0WccM0LsCBOrbso8OUuSj
dVEdA1j6pd4gJ6UPpBbxzbUF1mqaxa7/Si9K5hy8t6wno2FXOJuybHvXjIeyZsURgOCTIZZqQzkE
NvUJimlx8tcx8h4zCyzt7JGMBImI8vWkcClmrZ7ZUwiUdEs8mmLPyEaUn8YwuWHkmA2omkjb/7f5
q+2UBtLklbmsWSSSC/WpWQ+VasSF6mNOKkCKhaaHg65kb90IH9lFREhRkGU4V43ANcLgp3W1kpqm
JBNVHQlO6miLi/vm8BNtzeSLHiEQ4dYFGG16WWiaEyCfTYWbgTsxC/uyJD3BhiziYWSrvxLpG0/g
Lyo5mgCLZah2w0xXxzns1YhyadP6/cJTi/aVJo7WFGwchhdlnLZq63KRnFH5FXOqxeR/l37z3+9d
xo4svSL6MiFZmT0lDIfnfItWBpTcLExeIefxDb7zTnYUoTbemfmxv8/+acKS1neKJy4stXXytAim
RORFYEvgXYlB74aTu4Pm0FaCwcvFY1zw9ZI0Go8fLM+o4OWGq1M0piMILU+sZZ97BznOloViX6pi
QRBesD2Dg8HonSYtrQ1v79j+13TncbD5eefC6I4PvjmhQUXein5GfcMh16/+y1Sm9MEjJ9gN7qaA
/5WH/6mDlVgudOJqeCrWXglaLYPD4Uh+hF0M0PKWGdPzIid2Eh9ssu8sD69juvZlg8hZKmNyng1m
bWvT8IRw+KztqVk01MdOBOEGCRg6sBtuzLpt80qMNk0sI1bNHrwivsVODxXCXipGyGhwzauTl4eO
1hK2kYikM92Ah2rSBDF428lqvkBCvSNV1E9TS55aB6AytM1Bvk6in9rZPpmDU70RjqRbidXoQjr+
I15QkJtD/mug7z++Ee/g3b3v2QI0dchL9K2c5wtSp5pT8gth8TE7N1XJPfQYrIFyKHMQo4m7DJih
A2st4v/XTWcfHuIjKEBEMhZ5uf/BJlVvyr+bN9OHsMp+ZI05jVi0ObbFtzFngf3T3qy0y/CCzJzA
MGv7NhRyiEMbG2KksUTLE9ZJzm2FiqSjnPa3FkBXsT43nVw71uO1uwhzo0KnwAcmsSbYFw4W3b3l
32ZI7nnmUcjLCJEn87u2auajKQARiv+9h/RE+d8W5uKjyAtIzs3mICChOHd882fIX+HeqNe15U9s
vFMdQAjp97DLaFJeogJFQS//H+9str4NxrehDDvXnRxGgJubzHzEdB4ANlAG19o08KIfwXZoxsgQ
v0gFIHleh3mcrCBlTIIXhQ0eE8H399JIxY+QfBKy4cetcSHqDC3lTVTFd7DftKrn1CusQWrnR4md
cmyqZ8SozJ3rbXU8AXrqPwGMSZIzcMQa5++aL64gT1cWu92RwV4iG1MHQ/sGtH9Jg6sPf5/qohMr
2X3TAGISOKaOrYiWxaTd9+L8Ews7BBuA0GZvfJl1sdr3KXGpSwmu350wxCtxsv/nUvmDDoxkxk3h
YMyLPcwHyYXGt/PZ/StPkxUqZ7nCuqUJx/YCHNzUhmxngDEBMzW1wSICDL6+jDFDMnzFRhzXQXsA
tVr9Z2AD/Uv5kZLX+APLvJZP6tFQ7UNcxbwtozFMfBImCwqT6kp2ZEztCJhYuIxQPNEc4k3pjWdx
YZXDDVT/l7MfMu9HAw79mNWb+wsvzznXBeUm0uRGFCchp9yi4krPmgh2faIzntZwEoykRgBrWuFJ
1ZLtyyehVH7iFNF85p3PoGQlmuADCpcwCX9aAaJlqufmuk6C2u/K9d9Rsx6JYgVFmryGyxH+POJN
cKpRbwCNwCib/8FHNZSVPEI+LruUtRgk3Q3aJVPI/sb6R2XNaItU6d4o7ykQOZjQzuPBQfVDROKB
09jpwitQ1i7TPPzKb1GhVk0j2ZEMZBf/0dd65P0mi8ALBcwguKVcLc44RiEaOO6vf4rJfcwnwopB
OrzkvSRgCEjQQdMH0dRA2mhTHV8NxNM5fyA4+mRj79Uh9TilbbnBgJrTcRwF0juzwzg0gwVedlj5
JSKqrt5+2LGHO/yEqK6ft9B0AkI3zv5872Tj1roGYaBQQ6ZPHwj9IK6L+xJtJT2+J/bQt4eVooSC
Fc3BROKijmlfu1XoO5Kp1p0wKObCKEObyJFC+yaMYIcZXbS+kUsmeYyc4gz3pna6FmMcYjdyC5xf
pl3Ib1FgzMNhje1tBWbZ0kTA/xkyKFaqnlYiBzlm3fETKXSuYfJdX9/ZYPAxSslTe5EJc1QmTJsS
cYozH4yy49XPHbuBuxiW8g6EOCEgtOendceh7j41FsZdHnAVVTjaLlLHxTcgUW/w6/qcxUefxrcB
gp0nUudm5OOaK7DuVRH+D5cN8ZYWqdkM4kdhdKyAbha1dSTH/Kdlrnpdy+IukJm1oBe/FfI/SJd/
JuZ4EOOxU6UX2X56S9rC7sk6NdXXG0l4Cwspa3LYHTuDu+SV+rEjV5P52RS+KM11sFznCgsk6me1
BZZ0tHB8PnuaJ3MCA7c0ybCQLjwT8j/Oo8qiARmTmYSEhGxYTENC0pkqrZq0oO1rVPAU5wtOWNJs
rPwGu44jsX854q+JFdoe8k9pW1v3R3rtNXisp3R2QFWh2e0GgSDs5tnS02jLKuqLNhn0RjLpNedM
ppR5b/2NYUct+PPZBX4qUu42XgprnmRieVZeTQ6o0WeHoB8RnmvJWplnsU6TBoZ1szdcjKtoncXP
Ivuj+NyJzf872BRhSi1fIhX0PWd/KtXLLfihtGWocQ8QRpGhTe3akwT+gZbLJzLgc9bO9B0djx7/
0nhBdnv4oRgz02h0EcjjgRaeu4CJP4zdUNQCqID6YCNKRVEaF0T8wwnYPH8zEH44+N9vnPpQy1K5
XJVq6gKnAjf4KxNVbc7xLefEw2RJCPPQp9+AsMDS5FTTeYXMVmZQbENXHjJ/kfksDET7fA9Ear36
wL+vCNOISuMXDIBcGPU8U0CWcYVMZl/GKeT1J7dYGHBCH4bRKC1GNFPvJhnvF4gDKPdtkR5QfbkT
nLZccJnfSF7hJoY+toKm+DP1bwxtPa7VrDZjJ4myCK6PiH090bI3A/ggdqSnlFKmK6emHXVJJoT+
Xk5AM14b/Qi13+/5hh8gduz+FecG2lvLNntouDA90+KYLwIzNTGzc3bBcPRvqicKS1byQYonqp3s
kIzqoloYd3/cBcogcqZdgg4ahxvT7MODblBQ5pyjQvp+yTfCSKJiI3jIqjaQ5v85aFn8DGQbpv6m
2xL10OwAMtyCExjj5jOreK0WZeEyVHiZ4SYYeEcP3EIA7G35agdpVzx6jAugYJQ/gRKyR0BmjQ2c
+2H9OAJUpfNlr/+PQJv2cLbcWqOZMYmpgzCGleR4jBT1XsOtfjxyIjtPBAElcqMeoZbUNoc+Pv4j
b+AaJiKv2TQ2C0Krd6AVPQ6y6Qh2ieGX3DkTFntMjPW9h4OOdMcgHh9Ev7cSU8t2WQvLILrWGJ2G
sFM9mOgF6F+LwWArIm9PHFFsXrmtewnp2bO/ncNjgnoyVBK5Obh+e79v3Urm2F0PZ0FYDt2ExYqO
WeHsXSRGd4C1x74e/cUD7eo0Sp+6pGfDofCzDcK1z8G0+7x8lz5Fb7zGvD8XbYilVDksaSTyeyzT
C2KdvSBnSqISB7ENQZeIN9+bjYNEyvzsqI7vA4UPNF1FQy845jOt4BfojWB35SbDKrTWdIQ4njDY
fWUTVx4h2NfR9h2A88XVuDA1jrnfJyEo/ecmOBGoYVsBJONj85cevRhKhPdBO5sSj9O/zDGCExAD
egxYvrztHaFicoJQV8kBcNQPS8z6fQGbRa/rSKWo35ZKrJdrFcaAP7zptTxOByz8JgY/LYAFd2Qs
mVFfzVX/FhUGG70fmzkKwtNUSQq7S78LsxtNZoeZiazeK+0z0tFMhBG9QnJcuwYepGfunOhZaW/Y
ek3/3iRFcVLQm5+6agKCa3i/GAqPihDxFGvHH+b/rEr8vEV+Ht6frFu8kPXg//n7G5REzgD5ckNj
3d6VDvYPMbqzubT0qu1czja27W1fPtd6TclX2bj1YhaM5OaccxyLQ182Kb+QDxpHVC5OEbnU5qBS
Zk40Hka3iWDLzbYce3ZW+l44fvQvDbSawfbYWzoWMdXD8mYJd3Om8GLjTTUYebKA3SEul7Ha9u43
Dn7fMiyvG2uDGf894B3A+GxBuE6oeRAwkW2pYe9/5s6DlmjWzNMh8+izQ9Tu4xdE83+ZpZAQtfVw
DYuWCCcxBzDjIYiqiGgMbA3DGPZOiLXtF+oaiv5yX/zzxw8cIHo+PPu9oAclT1kSWC3CNjE6v4ov
fMYxQ8J5ASFul5MLe11PVOIlnLgTFIxtBbRCpXSmZ98PtCHsNFrDQoOqWJkDz7So1UsFhT/z/2oc
KmrjLp9BHx0fe3fTjY/Afv+ARIsuVWmj8mI0qNR8aEv1pgTyUmH+TS+gOi/CIviWdtuLmFDlGX8/
N2WiTERuwuvz2Ib/G+KPi4FBJ8PXJ0cVBQpj5fPrx76JKkhlnoUuZKK4EOUd8AcBbHSD5Xxw8zwE
N8JboMg4AYxge5HTPaCnv1ZmTx/SDwUiDOrsYwrdDyXk75fg7CrETWtyS9kLTldKhIbRSUCkDZjB
bYL/PbPgZWjCcHHs788v6RNpopzZouz+FdF5Qo0tSY5IPRkC4itC0vXY1FqFR8hI2SnGHWqpstS/
OkZ0xFyS66pX/zUFbTDUIilDnF0IY/xNqyKCpsjzbQ8HMM8PjDuC/CvSI6a4xyeHSSzg80jLqFO1
31trf3U5nSSYjwPf+Hq3wp0dANzqc1AUtAq5oiGC/GE5bXvEXCbhj2AvRVZ7xaptUir2OoZXExxo
wqDZzIiEee8E1otg3iDWGXh5Rn49hWG84eQxe04vSAM40dPI3LhhHxkRgJ4ynUQWCBtYKd2HeA5T
jRJbL4VS2cwCg+LO5+pNxvbBl81CWEJiRsaGpauq9pe8euy10q7TR7ddkRHBwWncgQ0IVN8NLhS8
QJgiaab+b34DTByLGuWWpg73hzgsnOtTScmD04/Mv1hFQkqM5tG9lCpjcowG4aQsNy9S/rYqOmJP
dyqtRuoXCGwb7o8P3WVOzDHZLf/R81ZSyT6l+hq0mnyJew+zHz+rI6ioFb9kxg8S60L0V/b8l14k
9o53dV8uSyleN/1iuO+P9OVKE1ZtnsbbDTe2y4zDjTWw/664p9gLUWPw9RnkRtG4O9QgKstBrb6K
7H8O93Ml2i5Jpv4LwB3BptDIhWdwHQU1JZz2jaDBEYIxkDHM4RBxRLREXqbOc5rP+6mylmeFiBuW
3MhAAmRY7ana2r/exQSoIB30h+L8QrabRqbwePZDYYWMcDD7MdnTtZw2osY1trohcyWmU4/EUCBK
WJjN1jeu6ivbGl7/mMD20wKutEWGmt4yqLgOo4G3vbuWu3O6JUeSzQGlraBqqvR8VPe7KLfjv9eJ
Lmi9hu6UGbTM4izJQeCA+Fpk372dCYQRBqwImFRnrdUE6JAtYY0f7CPqVP73i+NkhJKnFGY/hSkF
oqr14sTcvsISn/WVwjKkPiLM44odUQIAs0s4TY0N0WAtdn/3esbUbPGqM9FEwC61GTaaGy/B80i7
V3vs0j9agzKs465yw0mwRZeQsgsulB0/mN6jJY9p3VbDQJhRNt0vIMVA8sdFrWpj6pdY9KaUZSqy
OoyYXy1C+NcyW5BbTh/IncZYe8pXlSq+x61VBMWESQbYSd3/4U5oLQ1/d+ABnaExj/1aPoF8TsS3
TTDOzs2VJC6zu7OEhuCVuHTIsC4KTwN0fyDJ+jfet8D86nA+egh2caEgN/l8Gr+9p8k7LE5GB7tl
BzOIRusJjPpHtmBJ8/bp5y220KCcynWA4mRZk4ZEQfXUtOUD0qdWMnMmQa0jhbQw0RXJW6Ixt1vr
BLDKxsEgrDRl3MRfKC+nmJW7cUV4634YFQjzZf/cyEmHS2MtWIwbZqrToJim94/Cq7dRl1gEKpZT
0teggWsEx2wvLwmzbTB7gq2XnVVBtEgtRta4W5w9hjt24Nya26mPS5qaxlf32ZJtkxEh1+iO4HAG
jA4AWSC6aQsVFW+ErFURkEgJtEeAoCDYGENtK6/g6n/VGhLnS2ZUvEKHZsicxiUSe+2r8F8+grzL
4Cq5dIhZjl4pYm4fiNtmCHJ+uFJOlFdyLBu3eJCn38f+ZmrdhTAR1neSCUxzWKTbDYKRWXO/hN5Y
gWNGJf28wqmM9PSiF/rg0oA/U4BNP4TNitUDimzNMq/7kLG8oso1kR1LryT65wXqNSblwDyj0kA8
Q/djn81MMsf4L82JbnpL3IWvODHc6lT5UpgdSzd1zqxCjuHNv2Iy9Ci7h/1flJJ+2m73WN5WCoqV
LMPnFAuNslkKnZBKfR2OcLZK/juBAazAOHpZwajUvdbnNflu3OVsND5snx7e6dECZ8xHkn7nwShZ
CNwY/3EewiUuRcU81zU+IdDSaBjGGXx1XDRiZPtrKlKxJ7oSE8+wBcDM+/aKWJm+p3j/v66/xnf+
KA5nEXIWcODnmThUyfdURgrEXeGGOqf22NDEdX1h0A6ziot8c1EDE62O98m2cd9LhlKq8t7JXOxh
UJtsYuQhuWgfiYDY4/0wqt6h6iE/5p3tx/01a9s+7tyU4IH5F4huJ13ZIWxLFnhXmL3HAXPrahZX
Q1MKjY14+YHadjQ9wp5hBbYNVovgZ+6QlpkoYeX0ZFxkRhLbl8JI1tsEpJVytZgp3+zHgJXE/sMd
Wipn2e5MMMSxpFGttkx4iaXed4rQYh2HTZu5HVxYc/ktiD4VgPkFYUI27/Os4De4B5hpFEOQuyF0
WTxows+DyB6gj7UMrdZqbQ4rvGpLFP5/lZ4YAsX9jPyJcFNf30Ica5cIISXx6KDy2iwfHApE2VX7
cGb5tMY0I1jcWdy8DFvG2k39NBEBooCmFFNf8ghbiODKkyColRN33l72wy/xRzvXv/HU/1FTNCQ5
C2v81NVBrruLnIB+PKW8KhYZXgXQllXJzRHYPMz+scsojUL5IpEDNbkyOSjFJ66o/p7kpXdUPLa+
fvEOnY31LBQLs871oNi9xydmygFdZleZqRkv8BpWNJxQMgIb6jnRAAEdnCJ1DdOL38uoZiuNxUpH
OFEcScadu99BR6hA/4RCQtK7DWIeM6NSFtWkIxW0XSec/85IOYv+Dcfeh8RIzOv/xAfP5JQWHSPa
MEzvbMSmetI8rAuPoSpuAHcuDhfim8GbwYXBFTIHvWbGm2ipRprwZ/N05VFYUuTOlAvM1DO/s9vb
my4B+3CtjGHBL+r2uZu5Xsk9edTb5eP9UmbBJe+mWWS0uaC1zIYMhjzgIFKSx+McpWTOp3NvLyrp
qwFzStJCwguT3ArCB9h55hP85xBsRsUdc2oyInChVI8wdYPnOT8RAjNtmThoEdPHf1oE90mdiWI6
Yr27mn8Z2SzMIenxAmNUtXzATrHt+ozokro/ZxtBpXZL/hc3Q0YrP3XIWQk0eH+twd1xFfdUg+Ec
cinT6NrDvhDVPrQFG0yEDkKR/9rwdUyggWUksdT5mJxMo3sywOfcq3OAsMnh/k8EBC68hDwzyhnE
2wWH/6TyXzLU1a0duS2mF1GTfb89Fxe21BPb0+aRFiF+ugXyj+vpQd4E8I51AievF4sWD15jJwbz
z/jK+fP89eex0nsled+WbxM3wNNWM1+z/8FHoaQSy3JweuN1qMwntb5msUgkSN3qtl7blC7QN1EF
0Up0oKVdH7PT3rfgY16RB5mzOdRPxazPzfgngO/hw1sHLVsPUacaQk8TF34n6k++oVykT/o5OITj
4L3EYu5vR2eOKVPnnhkpeEXmWMEs8q2UsobJEKVclV6x7CK2bH20V2W1Z8NYT70s4UerCM50ZNVv
xxvvwhXieUUfVg3zzxxaLHD2Py6CIyjmTXNfpImfP0doUFpZMikNyQ0f9XdEGGXg5l0fC7UktNIU
f/6ArVdoEAa9nK+y/CR7scHi98Yq6B7dUDFYs278Icl3n9tYYfQ7QSMANrnv0FruGwWL+f3B5hPQ
sPhY/yHy+JkQbdJ1W6If35iySMgZCi4zFBlG09yQw4hn6dK4Zg0YuXzZCO6ZUshWKlFrYQMH1+KN
+3NVPBfVm0Z+5EeDvF6RJvcMwN02+/b8LAcTmNDbyPDaVaOTBOOQ10yQ6Bl9stKvnykPiFmr28Ej
sjxE2S9f4WHOmRiUcKRbu/bpUGucNrci1EYVQw4zZ7ka0ers36w3zYbiNnvYPeNETgluodJRxkzL
FjABoI8XkD68pNwTz2T38KR3LwwrukRyqJADZUW9N2U/5djFo+Br+B2nfmlvl8wm+5PxA5wXi8GN
4fmL548tvbLQ7IPIfT6Uz2xdqdhRVY5wced9i/qjwN+D5hX4fP8j3Hvsi9x0/4L0tblklj9+LV8V
yKH+Tqip66RFTqLaejZ7wbCrpZnT2ojbS05VQPWzDs3dFPDBJHp6kFI4cni0thsPeOSZeLcaoXUC
ncMnvOWP02lR8GXSDKot70+4onHvuI2uYV0dJUl48SYQTn0C4NMFlWA4nD0TPmUaw2be5zJ81dW9
w8dvKz+SVu8gYxcgd6RAAzwlTtYd81rgFgpJwNTj5GrtA8uWKh/iJIpkpVqiamywoY/ahoNPXk6U
yptNjHM1YwH3PeGq7nUDcSyB1ls0gqpaTuMKaWGQTxmPXAPy+Oq9YZs3D01gYI3Rk5NCssAmldS7
wbJwNNOdonKK0Cm0hvt9r6vANH52Xcc+ESRZUMrqCvBL+KhuNPy/pIKngKEs/TusqpEHPFZNmmBW
QvaKe1VuI0INyYgGx8x7XLt2X1XHmcBECDbEcp4JuUNSVTgNSE+c5uPXjByBDbkYsgCh0iZ6WJiV
FFygM3XP5klj4AdwWqcEqkzcPupdYbIPQ1Bg6gFjpE1znpHxoX1fcbp9oTiuhf0Yu24Yy6fDqPnO
5wyXcHXHGnY4jVJ6vW/9GMunfMjboVRENSV6jw3Vbaxsc+LbTpvgiBofq1Py5JhTHvLcNXMKL0aH
pQ10ZfDqPt2UtaNduaXSVtXJ9sd/H0D7er9OgiMm3twf/dqBrEhvSjuS5fqRHYMuM+uF3GOKWf/2
6IPMsYxX6xEGka8qkOAHuY+jkjRGbWt+Mu2sFED9VBeY8/p3+BY0WHlwDndjndb65YEIzbemHdSj
uL0/NQ3LAIvcE72z8y2s0unHmyGnRkUmWRbLByNXbnD80DNy3OtXpnRnQ1s8Jf5Mb2PQJ6FD5XCt
f8qhP92dy0LHurFxIQc3orxkWy2UZFTircppCdfp4KyfavAlQhGKc5Ii/gGR/LL986OSz8batuod
m8ijROwd4IDRyyFJZ8o8e4gwd5KLhm8EPzpvvTq1iWfWU9aE0hwTWG0emjiT1s0BqUbIee+Rrlqr
xgW/ynMNrF6xaWF9tubpwe6oHL7lW80brjQnP/lM+OBidBAa4R2F8h1/wXNdd511M9DyjlQCqdVM
83i+CA9xOl7ZWe9dX1H1cb+OtFfwIy47amZDXfSBVx41m3NiRPm8oZ2TISSLKcrgaUc06frRpOpK
PnEB5TBir8jTNpENCDWBMIieNY5bopA1Tg+OI/WCVRc6Tk4d+irWtTAL4DG4owm2pUR7CqKwafEy
nnEA4v9nV+hWEQdE0F1g5pup5XeJHiS7qT3SUUouvmErnM/1yGB8j6k2tXi0Zb9z6VCdDD+1W2Oj
AO3avDZ2TxccfNFfSCDqYw4JOGEfdo+FEe5ir4OiZlJJBPS3iD7pUFDcJthCFflvEj3zAdpVZ2gP
/G8z/I1omM0k+8SY4mJtPnSf6L2d/fUpwfPL5XfArTSETVAMjZsJm2A8Jpsa+KCyUBfJuBBLkJHg
qJ4rIUS3STIrjOkqJjxgDINZ87UswIFboxSKpLbe8rqpTE47mN6RbDvHX99/4HlNqehHqqn4nUhC
GQ10d6Zn5QTIo+ICigbop+sovK4yq2nh0yOg+lnvgXHwaLHyC5sWgAb+FVOpOW2ZmmEUK9FYzMlo
Gqn3VpzS0KbtSCj0qyopp6dIUQKufCybnw5wRBq6cPZzWYp+Kn/UHgqIcMSPl0YvOJyuyjQzwbrk
0GBp4jsXeYTQF2E2kFNPqOpLJIVq/2Z/XnMpmSm5awmu+vB08ksWhQ3TaZE84HyAyIdFKDIjPl70
I+4lvk9IGdf40Jy4hvqB1XJP6Jp+U1xhZUcTBk9HkI3mb25LgbFfsbMy6yAZS6gS2b6GNAfJErZB
Npz0wMkvo4HkzckGgj1IPM68+WAti6/uyehQ5VgA2kgn5vzHw1F03MOi+A/ehFaZspxsIpAQphHJ
Hj2bQhIX/7IHQKjtBOpuAFYl7UoUjzHeWFN6uB69xoIbl6RrAsy7OPXjEl4ActZQx+aJNbIqhIs3
/Xsb6IDoxTPC6NB/Hh1hPSxk8jhJU0+PtUI6wiMDfyqyNkxAbKKrVJSvwzjkfiWMTf0snCfoQkE+
NNl9rsxSXNE6NVHPvD3OU7rSOHxZmhINa50E0ILpgSHjNjyRaIcW7w4ErXP3s9cyM4CNn3pIXh3g
zoQthnFVqSMLFemRgs5Z3aXGBqiO53yK2MDbOiTl9kxd6neEHKuAiUt4BPdcvLIRf7pg803kQKmU
mTEJnZ5G9253Gk8g8rgi7DNQaf2hSE5Q5dg0ZSMKJ6WEFE4QKfONn6Qq1bkapLSh84jqF6XqJqwT
Dx2DjcJXNe0uu/vRSXDYGGkvxDPEQCwBQQlFVGg3cVOKwKisAxniE0KFAH2bjrqlC/0oLHOcOa/g
qZD/WHY2fs1dr90PJ36aiulXG4M277JUvz8uo7n5SHrB54m4l9e6XCMpSe+3Klu+xjoL+/r3htxx
kgOnqJXyUjFHvD6ZcjNAp/eizagMHM1l2LC/voNSD4ZWtRjQcfSx2En9a/6VIS9TUEGzoL69EjnA
KO6KX3wISsJ5oifGeWx2M5bD+dLoPAblnWhAAbIOauPCSU31LB1ThVnNU7/+3o+gO+BKVE1XIC1k
T93y1h8lIVxdMacapeg9KNbiEaM44UhRIIQBQkpZrcGB/Xs36H5HmkNaPHMQRA1x/yFZZLEQCVzy
cHSF2/ve36HJOw/6GfTTWB0ISq8iTx5NB05WHrgIwcuZlixqsrsGSP83Mb9U/32es+lSVTDwxPTF
uZ2ru0Uw538pJPPGzYd2U/6OIxlugq5SibkgAea1SkGnYEM0nBboC7HTH+YBqRWIgKeWqyoI3X35
K/nABdT4FL8Cfs9kP5Samj782vxYcu1koLGJfr9cIdvkOzLxnR6Z89cib7RT7lNHYLwWTa+aI80A
aFLdPdbXMm42gejaK3ZWDlf7haceLsX63UtRqj6gMcdKPGTC606SL0kmmojfNlDmn0QR0Gvzl07f
DI9gwfKwlXeF9QrUdkwpAHANe9vrpOddCabLJNe9yv1LY9Ol586RO9ww25Zsq3JT1evApQaBIixp
uafMRRAMB9542KyfHJaubMfzulKp+JpSQ+pSkjDg44RWJm6lokY/fcgdt6mtCIiWecKHsYIMpjQV
nQofJCAvCsmPtqwYVRbJC/2gNUYSqyavV6oMb6husgqn6H01Qr+WeiZQIjfn1mNMcb182jZi5eDT
ZwKfdCdoxp4Mb6pAP4SE6jY7y2lHZwO2ny9HEj+5hz4+HWRMrNzM63LIFU/ylM1G7VG7mDKEk4uy
U9Yvk8UZD/oWJYAlxNnwPpZEOiBrCBU1zseNsXyrh2TxRHGH+oZgUPXNQTk8PravOa9A2GBSqk8D
fBx1OX09Q95K32LJuc+AKtwrraCwrDEupJLYh+VYXc+3UpZ/6zfa3V2Jl2f6YgasgDFPVLs+MYJi
l5EZFTpstkMNhaEz82N34lEHPQfaHD7Sh+gsiSuYUSAAMU3W/pXq+XGQ9lvtd1hcnsgbAGiOR0xQ
ToSF2sxVTYwkQL6+09dsnMd8StqDWF3nIQ29nJ/RLbBOvfr84FCei/BHO8H6VwuKX7FfK1f+WA1c
vjcpc0mmx1ttZdUBNF46nBmrsxIxjOXGbR35Zge8qPcXaYlm6y37ep1QpOjeXVl0yp8xkxMyfbaB
tfJ0hpDmPFi5v9TX3hc+TCCeSkAk/Kequ8GdsyrsI5OuO7NlAXApY7CS2ZlpXR33US4V51xftgGk
DOnNY3K3Gfzhy2ze3Q1NKkRMG1SDuv9ho4DgHxUk+Gr8FzSVdrv4IIso0duX/kpDD+Ey5GCVNaWr
sL4OW7jpJbHfJUUvKiO1/SpWlkruQbMeeqqdwAcx8hWijFdUlEpJLOWdnCWvUVAESieQg7Re7rSP
IO9zcQFn9sLuk1yveBtHSPVbmde48JGIyUooib6bSTAP7H9onFhi1h81LcN3v9etVdVG3YRKvbxf
CDApQaiCnOHF52MN99pbtSit87nEAaLdGL/axKqGzZxyiTe/Ms3n1uELZL6R99EwalXgwlKp9nYf
Jn/dS8CuQj23dgYYSE2F84SMvH2grDsd5vSE3H2yvewMqcZBpAsjDM0HELX57tc9he0SA+sKiwXd
wS+D2AKp4O5MsYcxfa78wIymvZkTnlnuGUOn/tMj5QcJ/eekpK2z+yhTZuRf5WJLYwLWrwQFuZR3
zFy2sGreL/wd/3sNnwiR2cOpYiJDgdzMNK1QY0ATKftjd3v5m5fv+EPt1dD0WVzrbaujMOJPMsNM
GQHBiXwDex4IBeYh/NZDX8GQnZRjDlpwris5jrqvwJ7MVRaKn/wK5vRzBhznAm6ixO+pafodoRnD
QhLRQVJB9EZEN268ObZzoLKYJaGsENKXnZjMz2gJpo6faDDa3fyKFL3y94x5MMrdCQQV6RHKdeeg
80NELfOZHkcaFlPv/ZyJZE0nmdKsK1D/sS1bG+agF6J+FZM7q1h1SVFMu/u0Lgv0I8cVTfcQBbvM
l10+onBm2XnGaqvSDOXImBKrSWPbevKmmxrzf4M9l62PDo/OOa5sKgozLiCRzQ4tpocHV42UkGxC
bFCt7PP8Pvy6uvDigXrPnp5HtBVczu3Lg1RDLgbpYdSKH9gsciR9Ht1UgJg/gkaiNGVZil/vSRBB
QHybJvurz+OsjqgMwHswr+4/j0HM1bQQGyOph4pNJ/53r2xHH98QJkc5O3BJ0IYszztS1hU4Sl5s
iCLWZgi/J6kzzXMBdwHCibvA+i92DRkWDlMrmzEYafb5MHLD7WZgQ6lr5kYA12kp7Ihyn6GfIq6L
m3F3H2bc7exs1uSAX6SDiPHpKnjhYBX6lcJMPWAwIPxWZnHqImWHyVLOQBRJ7lv0WLw/5F359TH4
ZNJLMqmDCCdTAlep3Z+V351yPCaiwvnULtBwhKsbfwPB8iYTSXcyGooRmH0hkvRQHJbRbuUChgRY
cHJIOeOMprMpH2adIrIoAO/RJZh0VvxacqQaLGFKbpm5AGBTtUEPs2Gj1aHKtoibzddTJLFgSozP
CstzdP+cdrJKb0ayieisliBdVOICieZUVWbfs9wBgNYCM4hzFo6d+MDnaZ8aXHGpQOA34yywWC8o
IDb8W9LZPb7NDm1g4thFpA76NclHlOFp6rcb03PI3s7obXWQbGAdd9JBVkv3ZcCcNrGUPf3VjNRG
cZBc6WsCNJvzUDXGIiRynC5B6eadHbIvu5PLj2TBElEP+T2SZzNmJvDa0yPUy1mDCZ/CRnPbFEWD
v6jTTaSC/L57t4m/IW1eSEIh0/IQu+Mm+nAPsVdBK/Ic7nNKKHW+9xzCnx9fqD+WlFaoS5uYUmaB
bf+Wo6albBN0mln5p5hRZhT3lFhmGeI7FuQ61lZSHUnixW34i496eBnBse+sVRvis0Psn7X9kmHz
OwXoBWc1FQvpAq86MupuAGxRTnhKgL0A8bxD83Z+2lWFQLwRp3wqKpzqa8wt98rgTWlqT43mCtUG
SLFRJenWPJcJ7zG6jFIVbE9xShIhzYXL4NEZPXv9stcnjPKO5t+ebiX2F5lkjN0pZvxtnrztE394
hHQ4/B4bF6LgrfFNQTH04lq/IAxBtUpPYJsoX0ghgEpNhkegxMgx7MtTesZPUo6zPWqGhl/1gWFm
dJDewekNYK6OskbfH1SzCC9c0bCchR/mJIv+zcRQGZ8smHOennyph3D7dknugyga3qtMYiTsbGbe
TrMBixDxrIfX2UhhCN+7iSY+Qnn1s7Krmj14m71kU2IQdYcbyzjhvkErvkuu1ynsnXbmuZ2Tx43i
B3e4G01flu+efOEKStkMjIFCyuTn3S7VUgkmqLf38HADvnLrNiTFnH7ccQDkiq2KszrNwucocIuF
4QBL+aQIo/QeWMts82mzRR/9jvPTPh62GsKuLAHcvJNdh6B10JJQGi9D+u0LXADk66Pk+5tSE+mU
psywYV5og8uGmbGAp6a0hRgJNmS5q/8NHubmqivo2/H+bLWCd9CsJ40hU3iPxTLhcePYPA7sH2Yx
PZRGvdTJi+yB40ZuSCE1vaYIPJeo0JmPwE1ma1p6kp7O3A6djq8w2LpP9mtVzOKEGpoKPruJTJDU
+i32HlhZvkC9N29dBUUsO+kkI7ehaWlblUAjL4JSHElgL+BFTkJGY7GWnsFNd8rWXb1Y7v/LFAK2
tUtXiSAo2ZMFa18Ju2HSkckE83hhAChfEXvd2P6CmSgYD/01PqbLpI6vCaxEMbQDc/HQubWOdsrW
DSsZr3/lKrnG2dUwAdxSWdb4+MxbzoDS6RzabfuQ4/dG8pigXNYRGJv4CAsnaPhIaqCM5btAIJ8q
Gm53mjht7Bju2CtvQAAmTHhVFQavmYXQdwX7yL7oZUSswsSRY79LJLDFbjaAoJwrDb/Og41UseGd
jYuh1IuhkVL6DQjmJC4MTjZjG2dI71uUICCs2pBGOjgkn+0KcF0bW/7ONZQtngq2Rhs2VUAY4FCf
ubMCQ3qbGrNkPlkT9E36FMxtEWTSZwAg6jlvLestHXEfxcRro9vvik5LYoCWiJ1S/wy3hwz63LGr
YNiMCpnlJ+vOqFvVB2NRJby+3l2WsNHi/x8jp6z4eW/LHoEmKvgwm6L2utQDkIhByjbIs0YSJVMd
8M/GHm+UWwt8YeJqZw703uClBDGXvpMDYZhSN+F2xncp0zeLgTHyIlOQGFa0tGXudDsvpDPKToGF
x9PkkJnqsrkq68hqJsU0IXcsoF4TfqEByADIv7jtUztoyQqDkkjXnxsr6lWfkY8wICb0WXpv/Lki
YoxRjG5FqSpTJQqM6yppIkOd2frIMs7sZRCENK6EJpsg1qZn3yHSKgjzD8ZcYNtws2fFHE/5LtbT
CQYhy4jq/xy32eKyBfL23T+jhqCDgK4STF/xoFPrHhQjD647n6xqFc+HA6DK3x1HcOIZ9d4wfaGY
nM+lvvnmO0cFBLarGTtxRyZmHFq/OzYJvoLettX0OIFOUK1W42eOr5bNKOinlvX7aL8cZ1GssgnO
Gj/ElCHpu4aZFbvnONZ261CjPuWtIKroboRzbZK+BIeixkSQO3zwipZiHUx6CmQ+kYCn2i0OT1lR
PS0D/e7CZjaLHqXbeo2DXgR7/0ExXTle5ZNn/TktW3ploeAo0Ex+JuM2r9q6h7hNU8NfWKY1rN1r
qECGPjWUAffsT5NmAJ1FPLrouSXSP7+anOmzBxaIjtyZZlMMrq2RoZI5eOfuHdAbyEwxpQa5ASFS
o/43jmKCyFfFV8hljvRZjHTjT+/5LPNCRIUVn68spoisz0gbeqrx8BNlrRZjlWKyMGp5uHWolACj
13UfV2F4ZCOGusqh98bTCNn65STvmCqz2HZG+YPOkPi+c4LwOzXldkb5rTvJibOYsBhLBqWy96ke
Zph+1/NSBcoWd4Aip/bmpR3onqTHxBe4vk4WELUEPvaVMUNIoxzr/yjQJNHlVIzb52XKkcRSV7Cp
X8a+4cX+arI4b2EhkkC4qq/YNwqTdNeLZGBxkck2UeTnWvI1iyb8qGxEyZCVo0wukcH7FVCGYtFj
gw1Z6AxDi4MRt5KPsA65K41F2LV88ffUXcAb6pB+PR3kH6kCs/xWhHzsCKJegJqatBlSNstqB1xV
fOYfQY3S1A7Utkemn1V4iFTVjTYgyHz/+cLo8+yjbNY2GX+e0rPb/g9zngowarwnxQSEYVU1Fk3N
+2Wr5Dn/wndYswJU8Ih7UI/KRc6iiGxH3CMg+z77xpaMKFZ1fSTQ2RRb8dJ+Aso1dzVoIJZ5y/Ig
k1nKJwkPkTvm3bDsPdojxtkR3Zbp+kiUCzOWR9d+6BYWif9SNINitR+0y5CWUzEW4C2qW+3Gzwaw
5wyDOjb4lU5xvEembyre3SA/420lIKytJJkvLi3L2lPKLhXgP6/WcJRh0iLybzn9o9bpXjYrZXUV
y2DqrftyDBB5aZpIsgjT/pQUCPowyJmCAuuJftfBC10SpJy4mRALRNkugIE++fjdiwV9cvB0mYB+
uPoRxZDaS+wA7qm0oULGiDJxYgD6POG0PAaIte1cFpmK6hVU0TBL0/Vam2sEA+6bsDYZNqK1EgGY
n/IKqG36vTwqyfRjMmQ6k5psy/A4t1FgGJGxtkCcxVHYYftzoHjQ7xRDRLax80xUmpRercr2q9Jk
esVgNOeqz9+NRDyN06y5Zqru6oqDpNfLz1j1EyaHnA8kFaFyCYbyUX7e/DnHmh66ztkzrTKafBi6
Sn7OjLVvxNAH40P27GmnhWmI2zugzVUvIbWTfv3c9oc2RM9YshLdiQRZfWAnYiz2gDiq2uRPygsf
qsyLmVosF2eeymrWMhrGiJZTemuM63fJHqZDcUKCHpPjqfx/RVQ+rgarVVc72hpwla7118t55TAg
9QP73b9tZYf5FRxKnSu4rKIejNWFdT7RTDq1eS5lXw8Pyh64POin+msVjBg5gkRYnXlMdh2jmSKM
nQoZ3K996cMXt7PhKUDZnO8qtOUCbQquaGaQ+hZfxoOljua2rg4q2Epe14hQJF0O3zrxDFjqXD/e
TX9MTTwwrLD350yCI5SiC7oBlLhiv84KsYgzSzrnH34DmeWbmgb1+bQlTzvmDaN87iNM3E8OWYqT
gM4LDQ1w0OSEhurALA1Jpm+niA9s7Mi5iu8xV6XrXivHqTM5K8IOmMENgdufBRAtD7yAMZzqAChw
6q6IRmDNZSAlwDhazYZh6MatTolpMaW2x+S5Au0n9lFQKY8AwNgVhv80euysKg8w2vbU2EUgN+5S
KPfErLbOfcsGhE/4Tj7z/chW9kBgyc0hoHPWzuaW//0+hdpjDyDZ833zdYZPeDRIdkJ46cG9VUkY
hEp7stDVw/aIfQuo1EXFb5bnZ7PDBOgr0mJvVYRbs2f8x0S5CkPMoVTkT9p3rVDZTajMITFWD2Bx
UguguGv0E/E93DMKxADGkhTeDkKOG/0i/x8sxE3KXzPsO2uVi16xy4MwA//rG5CP8qE0+kvihvPa
QsKL5EmT5qDc7jXyDDdKJxIdQhejpW3e2shbD5WELFAoB9tkq4CvINTa6r5A1wGBmVmsNY1tKgu8
XC8uSCImNfaaPgmLnwyw7ofPg34yaItYeEBFLq+qJ/zbQy2lUHY0oMF3niRsOB9DYWh1mDKssmIq
FACaPUD+qpk+cceeNiMbT81jiX/wJJC/r+6k0Z9cWhyrNonK+c5UZdgVjX+7qYY0KPsbZP/+g2El
Pp2lfTw11ukepBG/uD7F/sep96yV8hnYy0gyuhC8eUm++qz/aczq8XXXSVeBjdhRxHzJJajoTVWa
Mll22nf/UrwaUk6PX1W3low6OxMhIZoyuR9di8y2tnbGDARIFCa8Yocw+TjV12Bz7sw9svb5H64I
UwemSqhAarz84IjkuOuk+mC30g/o4MLLZI1HZ5WQsd3rC3uesnh6QW+QCo3elhAorxcfqEayraOx
lm+1RX5eUvMGKiiq67eJdQZdg5lndFkIHepwU06z1ko9kOH0tDocGp5rfjGg1yGdBl6HhOtvml4M
gg+llYviQ17TDfBb5ub3+ZQ7Ww3dGiekuv8hg7snytjCDMJ+g9tgdhEP1W2xGv7E4WndrzD/exzd
4SUmPvj33fDOrXWzCuyMTGw5GTpWc5oRxeGmLn2RJnMvGiT+5p6v+t2M2W0+kYFP9fLtfp6QCSKY
csh2vRyePjqJko+jlSI7QH5K96xvjR1Vrn5ZB+NZA64iz9mgT0z94VBVHJCMN14/avOJZ5SYwdLK
rgQ2umYvaQEz6Zh4sHVCrqpGTsnQIfMvw1Nzjkulaso1S7ZrSRsLDwHhgC1DAfcE4aWoRsFDfnyx
IYWKLOPD3DHX6CWGXgur+7NLT+PAB7kPYzsP7mXFjBKJOlSrKKaaQIqLYnOfDyhbqf9dGrXgQDqi
bcyc6YwrOLaUk6cuGQQFJLPkPVqWKIJvVUjPEIf+jYunwnwGetQOIjiLtuws1PZmlMTmNtDb2N0k
wloFbBQZO3yaH/SNyjvgsXCu1nSHywdq9CopAQRPIT1yBijooOq+T6Uz1boXoVkIzS8DXY9FkwoX
2dEclfBTDsmx0AJh2knJwO6eJiJOoGAatej9Vl9JF8hoSAjMq4P1ZzawRrNjUijqOBBWrkkiGMi3
EpkgR9qQ9ic8+BbGU+G763PIACj9eFl6WGycO1Q8pQ//ecV3NvHA6hctq+VlKqorPAouP+qwY/xy
1et00SE++FWq+AHvp5edq6RtS9/UinfUcEaL5sgg90UNv10cgrloG6sN8VBNNf9gJdv9UizzkZ9M
koyf+DX3sS3qmIXyoYTCad+TBYKAc8W1+FSvavGsCfYW6Rz34qqbT6P6Cb50ekqv7iZ4VJrfN9e6
8oKdC3XvaA3ENvBIby4kiHiPzVX3lCjYkY9X8J2gC0BLhcNZwFokkMfQxh02O0yoK9jkJF3sq7pJ
JVSomiBKcXgSe0lHiNuMWT+qOKvozQBSpw8Mp0n6TQy0jx4zIVOUUp+XWwHfNMk1OP8lbqC6NKcz
JbFAxTviW1xLg+Sb4PURgUSWwZZnqUa4ipKAR1dgNt5V4AOygX5hapZVY+kL5cPa0M1z6JZs78cJ
fbZxVSuTL4xqg/x6ZbdTbquqe1S98iotFhJ68bHxNJeLPiLmFv3wguuez5l2yjMMG1DkJwW4JDz8
51Wj+WhJf5mYKFWmw9h68Um6oXtchPi2ph5rd+mZttEq3kCIM5VAz1i8KZMRPOkYmDawOtyT5NiM
1swepektckGi3+pZL+6lB4oJGkdgSg9/rdEQBI6s7Rc+sG/Te6XArAQdUFj5etBYohvQ5wO9qEYY
hBkJ8D5L2l3sveIabn7ZcP4Rle1B6RkivU5xB7PHmIqC7jnO3BG8KTESVt2f2MUL9j+6ftn1sEEy
QWX6uYFQmXZzOCo8AxMdOko65wd+bnHQcxOtHIkUYibcv/HZn3LWx23YI3zs+Jlqkt/octW2ArlH
oHCiCKvqncv0tic1Ylt0gnqR3Zu+qqgHtEIakqOmFCUDWoNoT3LLaEwMpd5qTmugfSG0iJbe0asC
AOrE6604MH0HrGk5BC3c5/e8W19clbSXQf24+gN/ogP6Shcnj+fFkbNO+GhsJKHvCydWKonrT8Zx
mldNtVTZy/vr2XqobiWGglxgjVA88JuEomk1HR1Z2D/BOQ8CDs4sb+znFfbtuJI8n0hS+/STOwre
2g6PR34IAHY8ttgCi0DXBx8LtoWfDlPkOw+a82tQvT1IvG36MOmKkPfN0+CBupJ1hwp1AjfVu93p
CWiWUx9DKcPPOU68yRTvSCMcihEoarKTwF85I7tc6OV3Ag1KuzUwdzJkECAY2e/9+B0USaH5OeAk
oxyUlNEJlp80BFnqQR5IqfCXOVaLz9chU5JmWVMSc4uXDFLrD+cvxTh3Pr7HtZXnR12CcOhl/yud
zmm/ulfBC0c++BXFG+uztZksda65vez3rwc+dm34eD++l1E49oMsMGdg7f6btBeUEj8e8pI6VVSG
4t2tvjQqbLvYAgA+JIUT8v95ljtcwQKObzvXX1VDlX8WkK7p3U1NUml4DDlEg2hWT/utuEBZlFbj
qVV8YPxDToHBV7pVKRZ5Gs/YsaeQmYOF7/OKlr6+dqq8PmrZbZqUj2nP/j6z5TBSCDRrqOTxIvji
wH2TD94FNbD08OmHjOOQ3LUYXV7j3WW1DUGa5HGRWUsRlvIHOT52b9we0EQ2HiCau9nZvJEjQgN8
uhRkHFIbMY+UbaebK7MM5SwEJS0B6gnbnPT+dTtHBeSsTKhk8qr16wWLW1EB2AMOBR9xtCJvMR9v
pRrKoM3IQa20iBML43o28IXjmAEdIz8Jp/uJoR/RgPMcrDHJsLjhFocRPqdzb2ZyJb+55VJVMtwa
1e+8CpJh+fr5jLpD5gx0OHfBkfTAsCkL/jySJB5ESqU6nTX0WSpUB9jhtj6HWoZPAOxxzEw6uTab
LyW59tpqHxqtVgGKMUKY2UK+qgG/OPF0LaTofQMF5GTjDbbwCfqfflbZp/VEopkbPOK1w/clAizR
mIG+UWTZ6sNsfMizQ7PANXL7PZ//Kd0Jacc/NpoXksRQ7jSKMSgIKuSrMKdfZlAo70qHKdcvrakE
LxKeif1FBADg5QdBAb6IWc/bqksz7avBCCouQe/21NXZxbtkAke32Aga8qquvk3rdsJvJt3zIaKg
Eu+lPCY4SonDXhxzk2xvoxclTQbQULox3BhANqVAl3DfwGVhtdkl6+7mlVfAFgtnOfe9rl+pUD0P
mLNedOSdE7BLFZa3XRzWX10SKWythniyI7zx/flOzm5UBYs4HBPDrMl5o5Rl97rzNuSg9reKO9El
dGx6rUnpm+WsLbla9WZjV+H1hIjVvN1ALKIQIpLNjTlDP5Kf4L6Wl1eTIWfYDyHSY1b1NW0D8fI5
NukGxAE002IIHMDqHIGu/bq/awjJjSsoeag2PZdsvY0RpMG/KKe8R2nxcC8ZehMgTw43FzOEoIuU
Y3cu9ErRzmUMwThm9VAaa3tLC59z/+SacPfY26Pb0xO+Cow0z4BudXgIJiLvZ+UbS3qLjA6CfP6y
JEKwl7dMW5EYoqlyQya8/4RGOTGjX7vWN8YNbCeB4aa1Woy8OazNWqk0EcnEFULPcfh5tWSQ4K0B
NPaP1uZouwGNvkNcYRyR8RfXX3ClVhwwnviHiT9eqPJLQPPnf1FLWg8WVB1+BHwuzaz4lqPfruiI
KEx1Emd6xFB6hNAgn3jC6/GbS+PlPH+Cr3FFj8LWkuc2dYAIbo1TdiRZZle+/avEIfJFJPN8Itd2
2k+PSMIYbk7M4+AFf9voFJ7voOERW4oTmWdpLDwZEO1dhkWgfecVnz5i1ZssYuhmtK1HUNbj1z9M
pvoWaK4sLlzKNft2vQYwwo4ViZNLljwm8yf13py5HwVlUboafEyz+e9c1L+/+5XB+/lUmX7Hbsse
nkl1HLr4sV0D57MfqGfvU4DpkJXHMOUvqgvMw2xkvkHnWaPNrqZ8/TPx5nZJ3gN/29rJOkkpsSF2
sQ51kprZK7TZr6JeaTfZMmhugwThv0ubsltkM+gAAljtALxMRwoGgzRGKyhIeP0vTMiF9UtOcMkI
SHb0MlXTQvJ6lSVtWw6hSmsQBo6yEGYBVnrvAPoEYJpqpZUgKAOzgdBc51X92lR/7U6229dPfH82
ot4t23UMUXj0RFLUpZwR7CUMgAY248/tLLnYli72CPjKYcDODb4eo9cEVLKju3b8yir3jLzdoBBR
A+bnYxNLB1QmciOu1bysTAABykXhRTK7dhlIhP/WBlVRZHwPH1VSr+LRQGFpoVTnIYiI70MmxCR3
JrhVasnq0LeRSwiZpMbrnopN98ghjuNsmeq9HtsrnzNXpDMJzs/P+Bnvv6dyglBMuApyBgJYZti/
dE++XYbNBX4jQ4NsQDHVz4tPQOVfnvn2OnHN5WdmLYXonxYWiQQ8Vm7aNmfQIdWMpCy36u5znRoQ
661iSchJz/hZN4B8ZigKgWEOdoXYl+9C6vcLGeiKEgY/vkuCzn1ijVnRgmUD6j1fiixK7qoM/sEQ
h+SMplpT7JErjtFpTH9w6JD7h1gLcyMEXjqDybch9rIA7vC0cfEyaaVYFmkP1R9fnItkSSvyb5Zp
OrOdZwLtH1OHMZd+zt3I3EpmN4AXFekvRJP+VGoXIKrnvAdizwosugDw3zRCcxana/05OXe2joFZ
gJPL6tDEXyWcsSnL753cefFwfoipXo9KvvT0hj8rkwzrFucgYY6Sr8OkIjaHq1bmrOBkoviWd1FQ
wMaDypxsToeTufbWgXtbxqopr4LkMmbBMNiEkUnD2Lmd5rKtHkgxrPcGNMgU/Pu8obRZsP6ZUnnV
tIT4XKFMutNq5OPDuEX0UMDfJyS80PrWjoigSrjSgtnWQ3/DcZCZ+Ol7dmP7kqZk07qZp0x6tksJ
ckj0G2sGf21N2M968aTwFdSNnCBeBPCeX5RndCwWNvY3AOXkVUIpuMLFm+lxLXoAqBJ/2TSSY+KZ
/efd50d1TTH33OpK9Z+YMcF12t6gi6fJPcZvOQmH6tM69KDJVgtlRR96x5SnazIW/MRfO4LkHaUJ
s150Sl3VzM/JCnxnnIV78x/Pae6cc+4LpoocD62CD0FJ3ZHVANJr7kGipQQphRWp3nS913w7d+Q9
BpWC6/tjAgmbSAEh9hMmyyP+GNHtoGXyTWI4h1fV76p8qvUn2E3J5Ku2lAGWVkoa/t22Dg//IxKi
IYOCJUWrgxrmLnvECbwlskNccI2doCv+e3OR/3cW1Y38NQ+X5gV7UIBB0twUXML3qFqybrcKnAze
MgtWwB6zP3ePpHX1pP1gf8EA4HBplr+9uOfj4QHMZXbWAZVRx497ixpr7r35Rvg6EVIRhNhwhtLV
GbyOL4PxcoSEDxuUmxPeyxqsuG8AVNe7I6x3ibX3bX/UobSie7YfUZzRPFh8MMz//AQ861QqHNkj
nwtLvsDdy3UfzCYV0IwkIYeedRzuK61swMW21EL6MmEIgvgszrcyznGd1fnDgFdQFThDvfTqS0z1
lb6ec9pdzngSeuEnK2D8j4Mk6icjGAudEJz4n0B4hA2USUbrGS2UsvpuC7Bep+UQYZFDE3QQb71y
9wPYDdpaA5owMLNmTe5RlYR2R876wu0ciubnznFLKYXC5a7Rsvp2J0rQIcHtvGdf/3zXsu/4LZQw
WdjqFE588ojCVPh+JLzqsLjfv6ywLvXZUGhFbgjDXQqsKM5/pRyylHqIoRfeQrwe4ohjR8BW6fXC
O0gLnRiHf8mUFUqqnzBcce/9HfZjfeAHKc+9yk1JFI49Frc+/tIk/dt7SX55SqDMyDynNJcP9b6w
xl2QKB2LeEZqoJ1X7//LjKmVgmFN8aHgwsFKbqrGgsbOVaVRp7fPvGQfS0aYbEtx70rweRSXvGsT
QwE7aoVwXneQLgjOjarDf6Rj6elmkYmVStXHpzJDseqUh6k28lWaQEiAlQRfUFPErH+5+DZPuAZc
YwuhQCb7aZMcsIuIO1WIsxLOO2VdRzSgI4QEwUddgIHjPMIw9C2J0aTy8gWCsZSitdqWU6O15sVg
T2xbAtn9DU7VMbfkLi57yNAIUi2HsbryLYqIFEipiFm6SoU+JINcYqYPC3+YFbm+pP8tNwSz00xd
WSbHBAu8jaJ9sB0qW5C89QoI4USsx47seRDbi7koELtQvK3Mh+jpmSdDSXeIrnibuwVslfj+ofR4
iKJJkrmS1+CJ+XOZt5sUlefFnGyR+vsQOz3p93mjNUhP0kL1I8oC2hEFN+4Fhw0m19OfwqkJjqpD
dO9QZWmJtHG+bjS1NcND9wTlhJy0nH/i0UP0gr0rQtQlGYYBKx5VOMhGJ7QBNTDoqYof4Xj5ji9l
t+mFwD/cT5Smwe6/G2HeJwKFE0Xp/5BuINZs4/7rBuR1XAxgM6CRVrjeqgWymLZoEIYyHTe8cRg4
83krSjEQEmX6WBHvKCMtREJUAt0Qt+Av8LqeqZUUJg6w/4akEeTCs6bZWFqKJTx0+J0JbecRIX+w
8rlPVs/j1ynxCUGTenU+Z5WTnCoP4/JXxj2t4imIctiU4e9C3qq0IneQj3ni66GnBGnrfcom2I2R
peJ05i+CKpNQG8A51BjjU6VROJX8rmefxUGihrIndn+mfuON+4ans6GVhEDyV8akPeSxPiOsj+8n
8VJT8j024myOpvGf80AKSu/jdM6FxambE7pYmEgTdXq4pbMpSg9xgC7Cn15AVBxrK3ttkAzZ4bRt
rAUZoWqqROJvF1itgRv+07OubPC6iIrYtvFYilG2Bn7qeThqR7CqwEqJ9sNvBPfSce8H4BQqKoL+
mYbB2R+wjk3JDnAPkNo5HFI+0Ft3yb3ch4X2/0o5X6kmt/2QH5XgsTSEwUPnUq3kR5BWtP9oC5nQ
cRINrcbSnCDp8xs+abfWoanb+Yiv4177kP8d/7JSgA0ZlGno8d9hAWmm16D1h/LMBWi+KWaYuzTp
4E2OIjsDiGOLXeRz9kBx8G6OE76O54nTwJUS98LaRUPMWnMNp5vC2Lnmx2wbRU0/2nuzlvvjuj/K
ueQH6GKj8jJkmJFj/DRd+6Rv1zFHsPvn4BNe6dWQq4gVM61tytmH0vWFL0kye7EXzae0Bx4iRiG8
Pbw5cQNj8/BwQULKT8fgfOMIvrh0gecfgTZOMdDSfQycM4fMUY1VgLNkCVtB5H1rtF45SrbbT1/J
9Htuf1/bYuq7V1SmIsc3dWIRRUIqdpgi6oxjwKTkIiDeUtn8T0ohADjagp54A2Z+BteZcaQjI3+i
9VaitZBfii6iSwJe9Shpawc4dWlbje6QFY2S41co3UQzu4wVt4mEYpkv/OJUv70CRR+nk3IwH8Ux
pMcblb9uyBWGlm0FgAj+2se4RzULW6YR6/qgFh5C10BoZDFAFxlgZhw0tHUYXjVBgXzgBam99Kwv
9KZkMvWdUnoxw6JYJKpW2dMVqDKldvri3/dddztlnOa8UPIpDS3uOECzMw4glkk38qjW3nCZjqDy
/m62jnQ1dWk2zAS0i/bVX9MbrOamK43e/yDepOtSGJ/+wPgDCV6CZwKhN175FLtLFA0KsC2sopyH
An4NqkKP3Pgw8hRGANv7QUzkkBHdSsFRZu/VMJeH+dowEqqXbTZi1KZC8sU/nLtZ+Mu9thR6vslK
CBU4u8qcTw6W7d8vHVgli2nunaDOiDLm89G1D0cFNWY+G26j0hSGhXZ9kSfOlGWIWR7/HsB7het/
j0UMkcHypz4JG6d3+UaAbF/aliXLUbkv/1O6MMCqaln005Mh7OksYwDLaDj9u3zYXH6w88KIT9Gr
szK98ENfSyQEwcVEbCKIARL143fMxOwbl6nfPD4/7tD3dEt/ng+t3lZR6UGnQblzJ9CTJocKxAhM
3YxzIWJL0qsIkqFAVA1qrQrfnu0uIG7q/+Uhn6HLK876Ash1rt6BEK8rWc93W4XedcoE/K7gJJIs
9HgmTJl5GXWk0IoK71lXzgIg/c4onYsmJdNdNHj2DIOtum3N0/GIgWIbKTJXJPuqMJBGA8GGIvtX
ffgpN9VaTznEOXNU5CwfjBUNXbhyBvuNjUq6+XBpi42JFJrIv/fASABOsq4FhdG1ninlIe1uIG9v
GRngET2gxBl0CRaNClVa0ncl/7muROozPmbqZaDjrdH185maBRyZLidAKliyBCLA4R5K/JfmwKI4
OtdoSqXe8Y16PnL1CCdxo3NEUnoLuT/ILlTDiUY1kT61LkZwfVgmcPVESn6kXYC5LJiL6pMzfp+A
dvm+tHCvF6CLP1NCOYRwlandTIuXZZjqc7a4+J7dXAogzD3M+y9+AJPd3QwHtHhYa/oAod8kEzCS
xW7ziHT8vXFAqqlUHUtQ3nAm6EwQk5c1+BMu3sRPGWC+o7bc0Iqjordlvx5P9gQHDT2/hy4u67j6
0V700t47iQeF1ajGjeQKdy9VeMwtxTyCSFSiFg058DbVLsgaINz1g6sFOjBf4RK9BVOY2voQ7a+1
cuqqTnkIw/tazGlpRJ7NDSMX9AWB/bUujCbLROIUBgSnBP2hQpA6MKhOOlcGc8WB6irbvJZVchlp
9ZIpJnh/6Ygq5mWm1NxIltCztYMbmIG7GyQbrndC4NmE8BoOEzEh0KFZE1Y56gXvHr7Pgi5YIw6U
2ezRvNivLPD8uZJJ40pmZSnrSqHoCG5nUpFJt4XUJ6Iz+EGvpotw8vOhUf3WyovCyXWbFpIV7Vi/
gGhit24S1Pq5wHoBe7X3acXe3ouj3fx6l3ceVCqrOUp39Xa4Sj6Xx3VYKkzbqoqFCEVptl0Zf/iw
2GwZ67/xHhMtZfXvi+WJHCpFXUH63dxM5FYbaHeTNlj0oAnl2rsmbKYgEvoCgWgjVzynTgw7iyKg
fCM2kCJ+a7ZUYIJptYs5dl6GcmTKd3XQ6s63glXkQTXUbZV60I5j052shZsMiLHAnV4oviVD9WQ6
oWJbCVXINL7ukunnoHp3koCbuTrD/hFuYTGVkkhFWUS9L7+SqgBu7QHiClH6sJFPgWGqpzttZCrc
dkXLH+3yyYQM+37uIxn36tbWkqOo3xRywHl/A9nODVBrR0gHmhI8FAIykA1eRuH3/+smvW9wKF5U
sRtsa5nkRUJQZ1ROUwBhtA7BYxfsB5pRqU38n72rCYsralIT1OMo5yogckHl5od+z/IUnmuUPxxm
NU+86wPXn/MlpgwQhqe/C6XqYS80/JoTgTmFkUYYKmklEynXlePiisBo/B+5YnmJxXd/ZbeOy6Vy
2oWc58f1MfVOTCTt4Inef+7xkWBZj5HV84u45NwRZdDHpwcPdQx2020MQoMDKqiId4ZiaOurD1I+
Tc2gLlJXEv/ayWEoTbXwqYYLEgVLiF5gRppnyEaiTm6OGgDTi/qSGNBbC0p99j/GcgRM2yzk2HrX
srEHXI67eNfu3ePyTNeyDYzkDlcAkWJM1v6e1XWCH9QbmXmlWafOfY0oKu+8xTMx8subFMHCwXRB
w3JMpDqEscQ2c/YdG2KptCEt9pKXli6tjS+hvXwFcvnwCMKTU8dkgCx22VOT1lvelHdys5YaCkJZ
EdZWhA2TyOMsbrEm59/p7fx67yeiu6aJecJuXEi/64mbD/q/PxYivXNSCESqKZwKojCahd/aVFiU
FG9g5ShTTevMFjpvFQ+OSUCOkaieBgwZXezDqMvr1E6poGL7cIzU14eGYOSBh4HSlP2qYLM8kjx+
AtUduB98ZeKD8cU/yJ9NHLY1jBekrSpO74yaT1IyRzoXZqStrT0vhY3mX25KC80XCMQojedyNLtl
3gYSYEgHuakYGLniRYoWDDgAlAb0h6Jxnm3WF4iog1Ishs1tEndzvXCRcaa3gRAfs8yJdACU6ps2
Dlrcd0cTJ5NBMtdLWPhfyeLlVmILIilpvA0pA77v+jKRempJ6bcjhSqhfsroty14CCUUOLwXUG6H
Fof+zWazhabcuC1VPyz14WgnaD+oek21ke66cusGncz/VCH+TS1DOxB5o1Pso7NVoG6Mhs4hGk7V
eV1WnzXiCgW9BuwDv3bwpxZTXYeDSv7mn0yNLtNc3nr274U7HK8dKx3iuJvXhhAWVnUwkFsDlYr6
5S0oJFvobA0zNyJpUFhvuQPdWyu9uBJgJNV/XCsrhTNTDCVLX92QzVkq8vTgjOI2yXowVUMbIb9+
k4o7qk1/+zw9IlJB1kUbFUOdUGgzkUPHdk18FvkNtxOL10ZtayzMqVNgjdRZcqvZsKLezN2i70qi
m/L7SCab7qV0Ij1efnmXgh9a/BoJavMTkWxKDAWiFiaFFzgMB/n+WfLE67lviMyfcIgQ9uIj8Ars
VtAmE0x4g+vdxPMhM+d2Q9oxrTTDvjz5SaUS6ELYmw6cO0M2F+aBBzsTWTdAn2tBrXYyGsdGaPN4
qb0wbykY8xeK+CXADHEPjobUp+A4RrSFn10WiAmVBUk/uZL09FKf2ksqADR8bAelcMpfBm1LZZW2
FsVzBMst85YUgUo5WY52Aywo8IjY5xxsUA3BDFh4kKuqObfwu9I+1vYRm8D9hS5Ob4XfmDjBn7Up
ue2mnKtyvErZUIkZpPC3ABPK0746gK85ie8t0kpLjcPu/HEOWO1+jNHfawjNJzFFhHcxUKf67cGT
ZzWykUHcXBMDvHcgor0a8Ipkf3foMOHUmSrZyTzBDMY1m5wtr9mNIJsD0J4nWWchsT66kz/L2RCs
HfGkT8GqXVRQ2et8jVvLs7DsPrXVt6fvaI9RpOGHejN+86T1G7PicTzXL7DbyZe0SKhHZ7UfF3GT
EXFCdFhjttm+/xcsJlnFMvFSPwEIuap7+nBuQQuFvuT6mFgEjG3FYIA9Oy52m+vzGm3YqHGffRbH
bkXI6dt+mrdwxiWzg6u+72e0V+sxws0fUSDXh8gu5OH4OEXliYfGgoMHmFrmHsgfUhzAr1BUtEVa
HuW0VlQkSUlLWFDOOBON/ZSjSKcvn4PUpNMLY6Jzh3VcOwNHOSyaAosrTpvTwFGDwSBXtpDsL06s
xDk2v3gvCY5dCw7BUIg2ahu7100TB27A1HXig0L6YFe3KKT0p+Er+0kcdhrLM372JFAqLPn6yhgX
oIncGhkuP+mO2+wOa2UQoy53jzhG1s2Z7ChxBqHVq+4fU4+cNs/WIdJXJGpZjFX3tfwerVM4URXN
gQlkijtS7QiL1/fPZu/ZBYl18FrsINgAt2gam7iZg6pIIhk7UPM66jZKPW0YaOo6luWw9uHA7R5u
iQj8tXfOjXA+shWZo+RIDaaRMWUd7q4UdzWNCtnHiukX6KGAnBHtPeY0m1vYseGa1N0yJdnqEeRO
CC8bbVaQIbHbiT1wQvbJATZLNIcxSX84ajSdDS9i7uHYucGe1oCnjSTais6wfKIKKVu5vRCOLHsg
gx3COcYg9CuRaM9zSVV3YTtSke98PBxljnIzLQW4ZKzX4jshISUKMeOCf5VS8XaFb6yWeFMUCtxl
PlemQxz64g23GfJ6BM6n0TkmOWp5heb6ljrBk8Yhkj2Ey/6x7HPmCIlJ6dWZG14UGScazd0bdOTv
opKo+tcEvqw9YnAxe1W8+KYS0gPRVcLWxrC+NzRaHT19p8d4MfFNmNjgKDtqOop1/dcbtLtvp2xo
4epthWmrPldu6fpwA+u2ez77rVF7omcMdhR48JeWe+NsaI6LFCXaytnQxyaw9VRCribdruSfqYIc
Z+bQNoC7xm+M9M04HZM9Fsv3UzHdtNgu/YqWX8vbkX26ZMFpg4MnOoMy4rptnBn42TkaGFcFW5KZ
R1+vlO9RF/p0jH3MwJ5x3tK251W2M8Vxjfl31owOc4KOb1nb7airfJL+Xz4O+6dmHVO7PPONLvvB
Il3Xpb1XdJCqQg1kQwqRnAqm6KSFVasu1+KCUAJArRIHdoJ1Ehc6VAOmfxlWhdQvFEsel9WUCGWB
svI7aVTNk38HP7kg3K3KaCiCB4j2apT6XVGicfH8P5z96YXMVLbZrxNrw1wUmTmnoL3Kl/8BYecQ
esUMEQfaC//sIAUGf+sieNkfCGxG+WN5pmmPSupJxpfe6Mq6x6M+zYTKL/29eGsP6b254se8/nwV
JrniCJL5aUZxAVim0fvfvmu0CCcDcFLEJn9Csuz5S9/VuJ4F+6wGnNGX4Jd4TKuF62B6w8rjHexr
S/TP3lex8Hzy6AF0Dnppg7LyI5eH2Fvc5x3pt3BcUySAOsE2riQecJ5LNjMitK0wbi4CQa2qfU7u
xSqJWzGkR8KIfzrVm/Es5BzpPUUL7HSdqwKUl6QqmE5OKa/Wjuois4RBvcInX5kCyqZeVfyIqU5d
ELok18ozgdOnkMDIKdMUBLpNHFNSm5gYRLmCnztjxoynIKQnLgZzp4AqIm2158LEl22IZFDVIBmx
8FJJDLjSN8/2kWPXBjdA88X0WCXgKHB7QCy9RFdnM/HWVHnqvE/8k1SUfU/DIj827yddgRC5qA/f
VZcYJtbs8yKOuXA0P+IeTVrqvYa2ed6Wm76bet2OrCerQdaoByS0MdU9GlyUBraQ72nth4g9vhz7
QtPK4wujdgiHFtgsX/Az5NuUMSvMRGT+I+y+PiuxDJ62MeLAYNswUxx3WEJKi7CE3W4+FTnNUwGw
k0l4mGwYpDbFV+ZjAoci4dON26gR7LHp5RYIxa+Oq8wtjyU0Az4J17lplN7MmPH37mUbRB9YAfKN
7lKtYvWC5syk5bjgIRYwKqtw0CibdanHk4v6jPNL7kdJCYfuw+NZa6VSawiZt2wZ71bgHrHPGGCL
QRUBrWgoso73lRMxGap2DF6aSJQkak/D/oKNqvZDz+JQIZbYTIC+DBOGEsi1KTWwzvLC22eg6wZC
9t9k18irOccmGNDlDfnNCoxKIWt2DJ8sRmVHCZnU6ftsobq6IzJOzeDZXXTsRm7kUYr7Bv/UuzMR
XaN7kjj2h6VAhJU1G+muo7v0/tBkkTzOfOkIq9k4p1qEkEPMQbjQ5D9yy5hXuAJGWQHwOPtBMChL
gSU7rrSA4YiHH0gY9ws/fltzQdvoWeqz94PGQ2jO97C3yPyIYU38rGAnU/SAwQlqz/8xf/7podt0
M+2Rkk01Mn/ulMaCDwXm6WXFiWaW2vHHH625U4lukAl3hAqq9M6EOyVPRY+gdhL83qltioXcy+S7
rpBVH4f+H2gACrT7CtwEq7EB/iENwUYYEXXWsb0CmZC2HSF5KG8USgIHBn/T24i+h5MhH7xA9qno
7rbU7CRjnYb950EGWnduef1jBurPp4WndPzh0tdKhSdxHtt9Q/votqkyST6cbJY4p4ep+nj2w2a5
X6iUetqSoawrnswn81eBGfSaNxWKQqD5gU3E3qkQiedPUrck/Qygpzq1jWYG+jLfvNckFp9pcDfD
j/QE3D3KkqZzasLNjYFLlD1D+mx1WLTSZXyanDS0NK4GntYf654ScIIRHKdBSA1RdNMoZpH50jho
2SmjAA40iJLLVTnTDm2ZuW0G7Z6h9qlUSinXZu/vXL36HKhkRApVPG/SDAuhyXfa/G+p4EmKISe8
NTeKDQrNxtXlxWJ2H5OtZFZVZx501Hfh2QTjcBl5JSf8nI0qHuHS4ABOjNkvKENwBaH2gvYyq6AJ
BGnmCpe5hWi1SdBK6Z94H2oyyngNoeMrcGPdmazIgIVLgE39a6CLMPc7dgaj58K23ZYz4n1XDOVc
5IMFC0/Ju7iOcGVMEB/itVOJ+hs+35rqCt1yJ8ecZJLO4CMiwgSCuQcDkkx1anVGrSnZi0e1GLNI
5kh8OGbIcLpdDNHCP19hcmkKlXE9sShGErkLllNyDgmQ1kh7k0wrN4m8r5dYKBQkSFPG8ui/NmWW
PtafbqQTxXGREnPv71d1cfuemGjzi5DRdRLCN4l3HIEPCUqNSTQOiwHdQhltOmbjE2SuaBhks/nE
AAqwWg/bYukHOSKPryMpnHSs9+r33bQO1y8y9NrYTl5PfkoBhY4YFFv/0u7sSl2UagV9fU86C8Ay
gGBu8d1AhO1gVAS51X4lHikbEAgFcb0BJGLj5L2h+ELfoBkLE157JctEI/tgvz2pGmEEhnp5z6Lo
XfxQQKlb5MgjSwr9dhxle5LSSTXMD5UFbZanzgGZRFZlw1rxaenWeUf9G2B2P14RTGSGcM8/C8ev
v/s2JHTlVJt3F1yqnljMOfQkwN4KbGWtGYeAjf9D+zohKN7bmSZLnWA2xZwCgEDeRgBIV9N3NzTI
qJHiUdxaXG0tN2XVa6J4gauWpCN+99XplQgRDvRdA5v+rk9FIPNTBORWo+4BX7HbU3SljyKYK/C+
qAklfxPuP5/o6BAmygHb1sQP9zOGtdwRad7fXmZ4Nz3nP2s+FbC+g7cPfv5JbH6HJBa+2OOtgkdj
BFsLOW+GFkGYyxy6nMyPtteXru+F+FiFeeBnjRgD0og7U4lzFpmae1CF3BDoRsFkzWw5UJs51cau
7T1aVFAGJXemd8KjIns+7cxthD61B1KW0Gub2yDLPs+FnsW36IBLNqH0URBNeEhRHXSWFJJyWpLF
MZXk0JMdNoaLhet3Vd08D5jmEman8REEBPGKCByqM7yAPI0wHs+TJqfQb0dd1cpLisLknriXXSgS
dUqJGQO+DzNtgDluB+QFF6QvnPTy5sSzxklng2YoUaGektFDXNfT5qirGKPoRsG9wLqKk7KvzGPz
EPWo4n4y1rtzOvb1ZxrgGEXB0CGdAUSCqxrUPpRmmavMN//qCfjmt7ahemUXZBzyqmzaW8O1+CjI
PrByFDJc8hWJWAvdTueoit2/6psHJKRtrluLbdeFH3nUgjdj6STldYMCO5KJNS4KDWJrDHZaEAhw
tegONIlTmT8ktwPli3vhe1TO5VljCcaGMgkGFiIEAezLb7Ko+GER4S1BUQAZ9hswgG7W5S+TuB5G
C9cyE5S2waX4DN5OgpgGypW0J3x07iBVnUoV9XCcxKIC1Ni1psDBFTwxpovxJlXWqQos3VF+9qlt
g1aLKh603ePyT1o3iEZ05Qv33hGecEdtta++XlESRVnc+XAJKhLkP+fRfUv2mlKzooQ7AW6MrV6M
IFgDInVNNu20nTspCbTE2FJv+Hn5mYWMKPpoj0SjtVYpdYsnmxVYWjQC4eBhInvCivGV9Ndvo0WO
s1FsL4Ef/VHxbgBK+CqtDHEl2DPBQWf71nrNNJ//ABpl6Nyj3mMJ/XWcYg7OHLKPjjiRIc6ZBChe
7HvZgcTihei/HzL828Yz6MaiMl2Ut/ubgHe5GsoI8hfTIvmbiEUlQOY/cP/dzswtCS1T+TxYlPND
aUabnKzuSyLosJFrpTWPBqbrgBrmDjka3L+cAyZujzAbOsh47bGVJiFVu1fXNmcD0KfHDiznmbOB
E+j8d5vlYgWrsxaoAFBQCQ9Lyy2Tfyw3V3/O6UoobF44NjhbYNdeBLQrPuV2sz1qCN82ktZAHyTb
8/ijX9Bji/DV7/htAO6kEZbUUprxq0MrL5+8gWOmAhQhVw0615tZ25ZWXYsDH4EKGRZX89AS7fFB
f9hAGgKeUuZ4nsEcc/jV146MQsC8KYrATswrpqOE8MYzbQlz1feazUeUTgZ8URlVG3L7PHCivOAu
0j63qnl7N8mZqdefWNs6NRODNOKGqkOBvrboNtBOvLWmMiRcq1JaY5uPQK59IGKWuOq463tqorEk
49QYn1P3QKkMSRC1xPzbUmBN+ij0bBg5nRE3R+NJ2Syl6X59ac+a1uaI69n6DhWJhd568ceUS6MZ
x67Rcci+z8IhUdP7tPg1MnaFrhnJGIyQbgGAmjfQbHdwvEKiThOW0abZfjLAl6VGaxnVJ/Z7+jS/
iH+NEvGZzWZP5fB8WGnGBooADUwNnj60tPQ1OX0S0D8+bUt16BuED4V1n+1GK926SXHAiIjYQ+CM
NDYiLUX1+EQqdMnr/WklN3fNdxo4BDFEIYwtytOahi7BXnySL4OYWJ803E1qCEC1L6EZDgZbOByL
MDnVt2V8D94m8lgTDNpN1c5FqG2MKlcLzyL1LP/WmQQyHLAq/EoaK/NhlnmUOEAxXmSWK7Ucn0MR
WaUAsqrb2zIx6rQ/Ks5NoRmQuv9OzS09Kd7osbE2BJa2bFw9praRALs6Ib7lPohG8AA3ePZ9Z13Z
+aqgifqhJmjqUtn4EdBUK+ayoYZLPELctux0mcFM3t3lKnoZlXf9EPTHE+PjjD2/MkiSbQ8SK/qL
KlGCXdqnbkoyKMbfEagwAFp6nswsHRGU9AFeDWBhmTpp7PIm937aUefhbXgVl9xuvV1RcpdiKP6Y
+NxFcq9QKxA9U3NDoobo6C/Y2IZ41bsiT+DeNpKwPQxiQS1h11K/ESithNcqiZf9MtAvetRrUyBF
x6XqAvNm+IIab3X7ng4OIzsdlURZZVK2SuABLICSMovIA0TTjG0mIpGHA9m4dvobviFJz4ebS6E7
kQpjzBzi88zBLlZW/cea+A6bKSWp/EJ6XRC3qnzyq9kBGWad4obP0e6KpplXGv2gvmT0iwt0yxc/
jx3cEnEibwqm4XdQhyOnp22o69YpaNAzXEo3eMdZMqWtHcZ2WJrteEqVZipAKO0a2bO4AhOLcJVm
O4dDxEthBf1gN1izo5yVeYnW2McockWP7g2heZA26MBcnwIay2M147mvDJ1Nq8V51mTHCJyaUq1t
cKm0Wl2xA2l+aOC6TPcs9rRsCQBXdxD6AeqKwfcHVGmL+D4Ng+dh+/kNAsWxPezInhO3t2R5/QHC
/W95wDLhcEF1UOn3RfKRT8QMzZtO429d2NUFEVRAjeTOMmSPyDnplLlhWucitwUkB2cZtmyzHMbx
GGQnnR9jkYbXqbNyLPWVnN+zX/BTJ8556b0WJdm6UmhM9yLcdPJsD+PBolKLHSUL0FHWTUp1YB91
HS6u3l20+0zmlvnNOyG9OinMxqRQgWtCEXxJ5TVL6yEOZ6pEG+C6+tBDqCpRGnDTSwZ+ii3U0gHe
N6yQxHWbsyMJfuCrlgfHaIZWaposhbsS9QAYq7NNAupf62fmOherHivO4OD0z7V0rUp+UaXFVu+2
0hP0v/OROAYNVdNRS8FlPmo7VkNV9vs/pD1Nt7614JKJ0agMyLfy1JF4HlQp02VCeIg8qHO/q3gX
YvSWEDQZSV11rF6qTJXPjGV/L/v7yeEGIlaIO51A39CWhuIG3dkLmtjeG6dhv1aqYrFdodMZG5ap
UZNBMSs5giIbqVsUiJ22b93ZHcmxkeJbFRJcMsYtXsqAeTqghm2Jd59RlTFRQTjaQsqum8CcdFHP
54bGDFoATxEtawiP+PBvio9RRZuYynUfugdTbslV5vGpByLVjqnOrCHebrtPZpb5nBD7rVx3X6o+
ZsFn85ViIqg3yxEU2kceZALg7XnOBKAelS+ivlI8Vkb1IR35Utc2wqDG13+iHfBSqCXV02e70/WA
inaanCnNibELwCqCrIBwOmmnrzLffDo4CTY2ftJXMdEno4FfQFHbyXxQX2zbN5ciIfUf+p9FFQsl
ubhXePi5TksxitDSE00BoGZJ3K5LJLDF8xOwU5Azu3R9vny6DXI5GPQM0Q5FTngOXSitYVDPJyWK
6wlQHh1JWQESBRXrVszSBWBsNyFT90oyufaGC1sd9Qz1ITGrvWFUpTfsFtA2Xic+sh9vb67sIJVH
qLkts3YaEKJU6vB769evW1do8c8Y5BdmU1z77k3+tieFWprdWZCRq2v3oSH4hqfw2mcFmlGd5DNg
K4zFk8Gfc1p7qyihBpVCRYOv4c9bNCBQvhFfJiYUz0Rs3fdMbU6yGa9HzEyOq8sHy/m2NXeAMbJL
OT9rWR234yxOVMaOmDDj474BxtEqDpyR34w8xNW+cxIDMJd6SZQgrGoutO8JMqXHBNQahNP50Hdd
N2F2/RiR4mUlxasTnsRYFehnBsLc5WAb++G1O0C7nCmwU0Ki0c3a/C+B/6xO+qCcHwa14ku9BMRw
DxqJXiE6JLnhMt2oF63c07fUUqTH/852c0AV4L+ImCy/7/SKJCsxe1xst3tNQ9GYlqm8R4LF4zQH
qRD5KWnVRfYwZyMJtSt3MinROXinKHK0vWcNYxCMo2HrHx+mpCbj5o/LQ/0KeGNN11YzuM0elD95
54KWsfKGfIOvRlJRPyepWe3+J2zGexW05vUIZQeWIIGYHc3Azpn5bRjgal/Jx7bg6zdXdss3Ujbm
fl4BzHZOhKYU3gTXRCJSGeECtleczTtE+hdzaElcGktKhEiwcjpwxbDLSGyjFEjd8IbfFidcPwU8
Y3M5RNjOE6k1fqkv5LAUWlVMG9NneBt5tBXKgN82R09ZJ8hPN48zpvRGRefZpcMmFjpFEVZImsMu
iK/Z6QHPTd9eHmU3tM0tQ9lWEHnyQg1WChrbxXojwMpm81M+wqM6R1jSAT3I5ezptWSy9QpnEDcn
w0zjgTCR+hOhipAeYL3P2ISL4bToQ0LiRP8817KlWifTBVVziFGS/MgB8c28zA3bwDIxEyuh/S6o
PEQMtXf104zwQojK9wlsGrIdl3BOm/5RMDKnrUxw9eragNX5xf+f/PIKNQh66aP6N2ljv1kLyf7R
oqikZAL3+UQKK+XIETKSbhCPfwZiM4nw/2nVubMtEqU3YPWZHMNaZrkVd/T6zPQY94UD9HuTBFxu
uk5BZtZMMXQsAd7HbyPugevkK7OlTGwIC8TDBtvHWurC6ZDiw4cOyiBmy2AVwoUUNm9ApImd3bXP
1wmzsO925ViMIqIt4ZzLG9/aJurg8ZSsJxk+rx/fnWy/YwS6gUKf2RpLlH4g1Ra6cLAU8/lxpWHQ
tb6ek1p4kjgy8jcf6YqyA7z5Zlu/YZF04GW7j8PkH9VhlkWeYhiEuSvEX/91SQMFrTYGFYQtnhyh
fkGG692nVk96vmM9Tu6SkiLAfy5BVg9eIYnyCJr3lvIEhgc/LMTjw7oT6ltE4mtcTJmYohNfal0H
2PCTKxkXfEoDSpewfxTvg2c/Op2FVJ/a96dzqRocIkwr30ABw4BrHf4D1NvG48M0WTaE/0BFy81f
uUivq70WesFeA+U6/Jx1GOfcuggsHVPYaeVv7D+LolLD75ucp8K09oIO7OjIacqR1/Id2J28wGNx
b2b/weUwlRgZkdHt2hQWREV7SiF0FkCjnaq/73gOGwVy03nmjuPYZ+yHCDXUQfKs3SrbFhntlOWh
Dtc3ILyDq6PY57fgWEDoppUA4VNhycKvxUTwJC8j1M/1rr1WSiE+hrZ6SD5dXGzZbS131TXgDgvJ
7+FWv4DluNI3PO2qpeClFxoPm+v+IO15BI6Mx511c6DlUziGgYNDqpREBuXb0hW18b9fJD6pmjaL
EbnRR+OXZbEgjv6nOs2s98xl9rhtlvP72wI1jaDC7SsvdVx4e80LQBWv05YcpvAaEQvnmJqzP+Hd
EoJjLtgyyyBfAXHD03nRihmPbtTGsjVYdJSrrtQN0bOyR8cKyGLAjlZXQIb0V/99HdpqtzsWVrIY
g2agUFkLbtK61uGa1hoXcMQcPXFWEzr6Z+hLpQTpZyCq+DDWPEt6gCmCPh3r3m8VgZP5RKqe9mFE
13CYG8PeduiCvI+fe70MTXAQKQ/2Hl0oC+bJ5brcFnUqFCcR28SAipMpiEIr/D1PXKdzHEUt66zt
QSBETj0TBhcUGJ38gox1pEnwJWzkXiNJRReKvm7CFJ9AAu40snov3y3o2vQJHTHPRmSuvcQ3Mto9
9DKVuQPHRAIrymmMygdqrp4szo5rYBBhAjhSubQ0Hodlf2Gtkxsw0bepLb+KUxepL2K2arxxBZnq
3zTGmpkjnAlhbZ8amBxy1gthHahUGSdeUo/tPBz+jSex1z5MUsAlpoAlntQCtujYEUTqTjdVZzs0
d66HDo733ksD2n/QosOMkBKpnBpYk9fAe2QPz9H6EOjXfi224RzbN1/inUWdVAX0M7SSza7ahepL
UT1/cOwmG0n942lMYDJk/hCVHYILgMZP85jPwOXUuHFhAv/AcC6uRC/FwPcPmuLkyGtmiqAY9kf3
BWwf+r5k6uEVeNmx8HZ2hZvhn97ehwhHgggSYaRKIcob8WEWnhw7V0TMYpYb24sCNdX396QpwXEr
ap5u5LWFE/0CaRA4X9AjwlwoG/dsxZC1NtAse8kZ120vE2sRFQJrTnwcW7hipnPGynyHpvE1OXRF
cr/pW50ONZdoHqk7CogBQ5ooVP4lvHQxAy4Ee/iSvpu++UCBCqGDQ9AOGicety9kAIkT3Ps8Dc8P
qjVHu5NH9WQYHV2uzSznoJu3G1Xpv1O76Y2wFbgSF7B0ZzDuqHceHbOxaEtRcqeAFCwfV3gdfyOy
VJqiycorOTfxWUvHbS1dD3woxn55k2H9Lrb/w8l+UJqUdm09zeQfZPxQEbkIAlI/P7j0e0NtOKxJ
FLlJKYkPt3EYg47nRvH58Y+3AB30o3kNXu0w4sbnDrjpsvGo8g/NogbQ5upaxQB0HuPsgMeJRcz1
ptZIs+GNbQhY0yhIpyq0qh4mzfthe7UwztxTcHNz6ooFlamWVEB1Zm9jhc/O8drQAbX+D6qzRo7a
8j2wZdklYuC4HSAcqRC3xPfDAQxEUAiMilkheFpeOEQdCE69rsxBCi1fPYBtS/2FKCZjkm24bdlr
nh8EjfwreHdHiuRy4IXA+bRA/zw4eF6RWBf3j3E+GYBBkPRN34FTQECVoSX+JBb9y4pRydkBXcSj
U80YESON5YAzXHzNZKbUKDNHIttEJACleAjDG1RA1gsOxthW2YIrRnK5vOOuSZk1eMFCMrOwmxRT
2bk3vkl7vW2P55GBChh5bE+6WFPPXLxMMH87IhEndS2EdozUQIdWGC1fsXHWH3XEANJ0TzHTYOm8
GbXmt9ckxSjug00kScnacK5f3phTt7G2E6yjngweW7NU5YLTX+h1ENI6akxzx3CJyBlPiUS+0lOG
0MrdpOBtcMXVE7XnK7ODAb9bdDG7schb+wSgHp+fA9YVvUHNTDhJijz5h/9VWpijl6golyXosGA/
dLhcAM/qHmzqwBJlwLZeV848yBX7fLyMrfgx/HIhY/vM4TOGUzxw3EGtFjMX5XGPNOSWsqAnWP4T
zlnppZqL+LGWDeoIDlf5hs5z/HWlpQawrw6X/mvGCM7gWPxjQ2osxsMzAZmaCaTI6wTbPxsQn9w4
oF7LC8FBoVX6yF27hpPJehw5vTHz9hsyS8zrwGW9mn83mxByPRXHvsgQZbwqVh4DrgpzTxO1GtiQ
Sg69y6aFzTeLxDisq1JiPbvYSAln/50p8yz8XC/AEUhAF4k9tu4G56XBBqsyeV876HKpu6hTADB1
oW5k38KrUxJb1bmO4WUfuYv8iJSTKHaX0kipMvHY83sEv+wu8BcZL48BgaTzJ3d2dwwkwJ6bLjA9
7wVCamylkNq1ZL8PTDw6i8Cpv1N/q90fGP33NF76q9Ls+6GE2QtmysVXrfYWoBQ/ySp5hXQI5oDb
RZhm9SoVmO247N6yrtP42DiVEIdfclvcCjRTvjbe17i9e1exnhQPmoG6K3IDps5pX5G6U3rrOa8H
z2KjHy5s8EFhm6A8YXKubp0HUjOG1jOpNqnaux6a1mU9BZKgxRAB8rfApw2p7jmgmR3759oJLNz+
8GknbtvvhOznye3ptT0zVcxNXDlyYfKp8y7pJwybTnMBalel0APGwHzqKEsyXL6//fT/rDRrxtX2
y86QCCCmURA/YYVWNwf7gf/rItk+oxSlyA2AQ0TGta3jFh78JlEbmF2IqGHr21jd3uhqIaCUBJpw
Em/aGhizxlKFCxO63ZCXsndrCHc2h/WRPtjYoWxAp8XWC+S7XVlnqbsBtIXx67WyN4Ye76QSAouK
yLCAPNpXdM+Hm9MxZbAWHj9rFxhY/evfyGA5SABg5jIpMjuILw0JCkGYWxETq0+tmR2dApx8F3qD
UiB53BYUZuRdUqbQCMR65UKfvqBkRcCzZjJzAx/N5hQz57+NGbhBnu9qURKBda3HECabkWfPrkAG
39LWMF41hZAFYZQEQeMADoGYGYIas6SIv2wvJPZXWBMPrlRF4mzAhc1bji8xoyS1aa6JwBXckl6h
xs0uvp/xAYKp5gwNht+VXgf1Ug1GfreaJQWge9yMfijj1Q2gSzi7bkaDSzM89toND0YVupzGl7mO
/VBxn++fa8tLI9FwjvJD69TJ2QKgtez5jO619+PvFidYObtDt6lUuQKi6iK/ju/ltxXObGZI1Yos
vP06cKv1td7o7IFx846iZL4CtNYEZlXAQt+0AxPONnXqqBrWr2Ft+uR+Txs1UvoOlfIRwWBsJyiP
Se2YXZG46XzfUw0nbgOFUzxRE8vDr783IOqN+lJ4kMDVzIQdLaT83coyXEycfGI8yGOxM9S3xai+
H3sS2M7kZdfPC4JsC6dB/KkAT+gynSzOt2l2mhz6Vbvayen/QMD+4n+AYfIKzrgTwkDGXE2GKbGM
U+83CgY9dHjk//j3nJCsgLaxOXVs0sN6uQ9TuS08CoC4WmZzflx0xh/0Qgui1UwGUR2AOn3sDvSb
3bkNtVVIrZaKF/KMWcbYesyYncOmwOY493ixx1gMbaGadGUJk30ZGn8/rpKYo96zAcjNcC+KfCXY
La4PtqiNmPzy4sbBxkWP2oqE3THc0Vu4i1d7C6Mqd8XVViKMa5vATBGxoJAjB8mywia3cVVIdStI
1SiS2Rfoan1jjJZ0XbY84olS2oaZ5tYkT6va0iO1zH6iMfpbpr6HQrgPPtezjt7hzxNiEdDewU/z
uNvhIV8eOzpRNnUqN7viayaBAVmF8RjB7kjsdBrYKbFYvtrekqVxOGADWVMTtbCjsf0qzxxTRjCm
8pmmmWtagR2pIwc0mU8yPELzD24NWYhBGFa/AeElGH9fZjpTkFBsDpBMDPKcLKeAwLFy9iVwrHW1
CoggvCo5pjQJhUu92k4qRUKCrN4D04dHBuHMGdusta+rXv3pnlb1yT+JAczVIizs9v6bcDDrPZam
js3HkYXXa6ZscI2NeQoHUgl8EelVYFNCmHmM/Zz64p1xO6rfJc+XxTqpEg3wgQcMkdsdx3agL1f+
cJ6Nb2i65Pxu+SXtTj3hoQEeZLFc+dZai4m/aC3q+AZjeKvikbMrWB4TNM2svYc1RfpqfjcxtOF5
kt0vgD4S6KZqI9vPUs3VnwOaTFIArkuNvBS9IEpfXbKKOnJ6/iDqvO9RySWbc2vqBPms+mFN7iWZ
PSlTajmZOpETNdmYDYMO2BvPqd+QFSJX1wcmh4jXumwBP6+uDmNyBj9RCE0LLMFtR/SwVsL2OEjY
i3PesYlma0VMmSLnqkElNR1XYTW02nAndCiRjYeYPXMQFNnzbpoTqnmqCYD0jpNr+WHmek7YVhuv
niIf70hWLH7SA5iquxPEe+vBYKrob4vw5byNlkSt36vVjUAskeJ2UAnuDYy94kk/3vBOr1j6yqfQ
Rbwg68Ff5DdrKX7UVoP9g7SrkQxYmAzdnki+FN3uOC3lrZfGsIIjOP2V6wavAvIe3q8kzIjIVnYX
s5YKnzf/iZOEtg6w2cW87XtpO0z2lnAZl/97GT+eKAOy0KEn9cAjgBYJY0HjoDR8jSdBd4SQICCB
lmQ39ku+JBmHJyKZIQQA2Men9UOXR6XD/olI0w6T6rSbHekjQY1KhZRhBo5wwll6rT4dHLj20Sbi
ALerGYO1WJxuIELq8WCupk4SOoCqfvlQb0O+aOF4D4lSJ7TB4DggmHsniR+ybawY+E+ZDFQLPIF1
3gbbNsOHMM9f7UU+HqxV2OvRcVb8eIOquMzxDqh4wPAuDyFb2snz9sp/UZYo6FWqbTOmvOOBlntW
GyvpyZlK3OKrjou4nB1J7NJ6H8JYnY2OCEoLKPGP4iTZG5epUbtXT4u91WcncqgelF8EOlm1RgOx
lP9esXxgsKjuS8BcaKIgTd+Bbeob0jBhYZSBujFEKc0aC1/QlpRoDHsJ9yFGYO2rQvSspVqI7Rcy
Fz0QnJEQvbVUdCMYhwClJuIqW9ySYSD29hS0ZtrvMRJV4ANRmGdhpv9dTp9rE20Z+rW7yMH3f5e8
Rfs++YIF5VeLou6kVEChLpYTXrepLu7tHK3fwEAmlhiZ+lqVZ74CpHLWjzkwJTQU//UjEoHXb9mO
kbpggpXs9oB+tzoR0MEnNVmiqzTR8CF9Y9C3ljn82HxDuHUx7nahpPoqEO2zvIozFEU5POipsjgW
TDp1G/KRCtAVms1o1B1ZXFBsTqkReUWsDSeBSsJA6GgRXwrpiCsZnqxr9r4m1+s7OUpT49Aer/JQ
8852FZnnV7/APxC+QrPYWyfLb1FLnLeirGGe2iAwsoyYu/VxZZ1tQcR3mp6xwmubl7qMbmkugZl8
1UW/bXNkg/KKtOwA568dq1l1Wbo+qayYogsTipSPUgYCQNWyAk68lV41mxEMFbHrtbeTlbpV7COX
DieIlGxgy7hTq0pj9LCZ1k3As1AeniuEdgCsRCJvL7TRwo+tao3Le0QAXOn04N8Ir53dQuEfQm40
CMuBxSPnCsQivrg8/PK9zSs1ITDei+pWC1QGheYSefJLlP2cgHAW0vK7tQBWXXRfYvyo2+j01tf+
9pjODV9D1XndhKGTfxqoqI7zAJL6jPNkD55Z054F8agfvXAE3n2FhuUmJyWVO5c9wAM7QReuciav
yJi22Wm+xwYL8rq9Z27RuJ5aEcPaGq9zm1V2crcnwXfjRua3CeWPTrEzgstDvlM0DosgqZckbkPo
vVBRdRr2t324yYwKBETgATABxxl1uuOD52xXlv3W7wvsIK2jxCZMa9m/9a2A5Xgvuj4I8w/kNuJe
04hI4NYGQb3T8rdaFBznpweZJq9iVamNkN/katzsCIUBJgX3khvZo96S2XJKln5MOsYZ2JUZkPRt
C/UggQORDYVj/5upbhwEkkMHQHiuRL98wCgjSRRnq7IlRgq3AaEjit1B4n/Z60JCzh4309A7mQdc
hR9jXW2G8CxnAsjC6mx7ANifW05UWPJ6o7V4pEhCxm9myAGB9t/Qo6ih04omEyA/px/4qpvOYra+
wZR0IzP7ff8Ut7s7ihShJm2yQJdfk4XjDUJcIFFRe/Hn8xd0kNbG3YgNe1YHyRl8zErsQKjZ6FX6
S23Z9S2Zs7Qps/Gr1BaEo1wZDFUwpL15P4P4vD3PSuN5aaocbvmzWtj8/gGYKhESfU5M98sJbZlb
A/j+BvKbOfzi1C4H2UFBTnUvSWFAg4Lyjz0ggshJDPXTLGM3zgW35QpRcb2yM5VksB+6eWlWo7I0
dzHsK+SMFiG1fu5QjK+bikwouRlgyxbbkLEdpr5z0lQbf8iTMEUgF/RDavirTiWwKpP8IHovVM3E
ZZtTdu92THXa76T0Id/TjJgWbNtMSxUN/S4F24OA4e5r2JZPPOb2II1b4Ts4VktgBNpVNjx0DfYX
tEsT7xj54K6GiMQJR8a1MGqp40gUh63NAjSAZlh4d/zOnXerIzdP/v18gA56L1j5rkxz0C/nFzO9
6JuEYnuOvazVfTNZJ2SBwG7kt9/w/yUDqC+1Y9lOcFDC5IHtReuFLl8m/rYZNWG4wlY3Gmmh1S9A
4fty81fvw+IGUxiI1l26Pmpql4ElDdKHQocM6I5s8fe2yzDBGOEEM7Ti5BcTY/ljnEWrYsG1+K7Y
XIHX6RcDUBwp9YUlPuN+LZuA1ucXoqeRoD1DtuRTGpTEYvE9PH2MrU2V6YDgQPBD66ZdC8LKHAvw
WNqoUNdUL48AQm+3h4DqaYQDd8fJ5PG7wI59RXalpyKNkx61Ugo2jgN8qe7u6FkKgLBNYFnMdWSB
eWEPq9QMfarA6i5DqV1jsZHTYHG9zWHja0EtKa3FUQc590TPWz0EZcwC/B1AqmD+SJe3Qr9GhEv0
NUZCnpD0YixsIngZ61I912p9tMyAsEg29X4sOG5y3/hHB4ssJ7sWMMJ/KQ39G7p7T/fZkMDBQqz4
xvpaTXvP278r6kJ4CuDEWE2VudMsc9FYWv/fFcupZvXUz4CLH8zOtRpFIscv+MqhNkkuTKotz4lb
NziWIyJYvIekj0YrEjrgJYdwnkv+DtMM3Qjf8gOyHyAu8zByjm1LjqtXW39pOkAhp80E2O2zH/J4
3IPdrCP3P12P3wvk5NsLN9R7tAc+3aX3yGH2MLjAdtJvRiVRWfUoFCQzW7yOwUx3d4rsI8e9FTIh
fD7AVESRO2+OpilUIKGYlrfpKeCqPmDHqn6kkugvxXu17TBEpCZWRpF8GerBEltg7oC7DwAcBvAW
0NGZKM4gmg4yYQfWvCv5ZoASeTnvTJsyd8nnjuE7gMUAbJvASgBayLdjuWc9HRA7qLoq95uTupxi
U41S1j8XyPtkjkpHRMiPdBnj2B1KkyYkFTmG27OfYLd87+0Gh0WsOjdS2G/ZESyp2drQLZFr/i/B
sY+TzSwmDCxgEhyHgb+4L5ufb/yt59MPoYyoH9SoPY7vsCPVKmjaj8dJ5PJLI+z0RR6A/CblSv/9
N2voc8ibi/6Wylwbb+4B1dyJSRH7xGCt8NaHhg387nV9zUsm3gdNA1LxburfwasOSMnPPK5TfIyk
h3NzBD8TUCdxUU2U4R1ZPp9KwD7/MkfSnGBBaYA0r+9tUv9PB3Xcc6fIomTNqkVdlXopXl9wNsqH
woNzySxXtbmxmLmuepE87e6NT4JFuny/cyen3ODSAyEbW2+ta0hES86vQP+DY3w9VWrhHrBUtbI9
fYhl8wgyN++5I5NWgWAI/vnSAmwxkt7VUQfrqJNIW1KMxlvm48X/wNtPdhdqzeRpTt0OQNl1Fcz/
9O8VztsjGC4ScSVPpHyfA4JOFz6ojmSo5Ugz9YcehtiEu/mf5741p8lVzk7SIUWLtXmBvVHb2t/j
tFaWrpG1oXj0dzlTSbYWo3Lx4pg4CpAY9n9uFOQbwSzKg2S41hGX+2+Rc0jMns9mKc1rfKpdrJ2p
eMIuasU6Dd+bvwGD23z9NKK81+nBS5PqIQvmPdGt1shjc9rdvxc51cB3KqsAAjgQv1P8D0xiPuaB
b3FpCt7v6fYGbxRf/GLp3++OkXGUJgvsGf9i83Ly8Zuic8Qsjg8+P20JuL8X3mN9edmqjLaEjYN6
hJ/2K72J/zhHneDuJm2DDm9rkuUqKp70et3i1SFEIuZ/WotyEFBGNKs2dUvrau790WOKzAP/ThnL
DxdbsPGgK16MWxk6cxxoC8Alm4XH3vCAI21PczXj+djMgfmnbYmEj/2zCPvoK7ZeiTdydRwt5Neg
D0I63sbV0W02104PRH9mppfTAAwlAJCUza3hAnPjef74mfUab2AKh1RDH5GCoHDSlyHC2x+XRSVW
Ak8wAQgt2YnrjcAROIXD9YBvF4Zi3dg7EkleZn2AYHnbpwgALVuiGSqsGb4Iub2hrXH8+PIQJ0JI
3WGokjMqi7Woq134MwrOqXnOcb/tYIrEdP7O6aPrG4IZS4MvuQA10VNIgWuEvdh9o88KXyKdoxoJ
1UsjaIfREseWQe7/6SucUUGO11JikTZdXB5Hg8r9a10HJB5Pg0SNr9m9Lq6F2JRpKpoKVoqjejY2
Y8wDL/l63lqezAJMDhir90KizLaHUbdDvS/M43EH4w7DNXFMRsxJz13R4x4MoUGdIEyAD/H5KTn1
GTd3RqJa0SQ4xIOMLKe4gLxRbqtRrhzWPvbWIJ37gPwKHrO09vBAg6wlPWuXz9lMPtqRtX+bAWdd
ihI4DLz4UATVvHMHzbTVob0CnXgMMbow43kSjyY7shkeMRN+WRg+v1bnqIZ/j7hilDBQssYrHEF/
GQCU2g3ifkUSi8/I9lkfN2qSIpFwNmlmFC9JklYpOzeigCL1lyMTo77pXU/vZG7nhp+UcqGKLP7d
5on9oobmobbHTZVweCnGuJFSiYjgWVDNAZaYt4d56o4k8WByvVqOhNgUP4AfWUzjITFS30ganUoc
uStioyQ0UG4inpzu4NOakjDV//1+zU9N+GX3eVqxoh2NEQYLixZPutGD7o5unH83qZ2jW/kIC1X4
4q2gwNe3liMLFIHMH+8Vp+1fRmEWEToeDeqJD0QTKVDDywHH+40ZqZ1XpL9P+KQ7HbI3TQdA0Kv+
UdOwkZz85gSh2HEkwo6uhN1pMN6diyKjii2mttnnwL4zcY8nBt4BbKfBqfULbQ6EyzUwjGSDzwtp
JlGy/Q+YjYkuGIzuPqQ3zmRpoxcSa+COaoU3bVc14Ybceg7i2KWIqtwBsti3EbsIo4Ln00+QnU+J
/QbkGJUKedVwt/XhzP5DY9C50rxaPUA8CJljESufrsEfNwBMU4D+xuUPp5G/l4Wq8HkceIoUyaT5
F/I0iKc86XG1/NQORftzmxfeswxH4vvo9F6ilqnUjv1+dXKRGJDdm0Fb7kSvTXkg1rbitUW5n6ax
WfIoH2LCwAxCh9bHf/K2Sy4SYZdTypcy9inApvCK8V7Smw0JF2PjV0HDpseUXVaFqy6h50asde0s
qasJ8lGhkGP/9vnPH/FS2phhXeb2dKUmc7Ydni5yo2YYdSE0I46Rz0CVsWzt1bcRp/flURvDC0Vs
d8DqUcJnH8FVmMrbN4G0zf9jsJAZH8nemZccB6/Goo33c79tHOe7Jzazd0teVkKlvhf70Nvpmy+S
VurcH27EgT6mteMmzjZ/PlwNiXY/9Pt0fvHBV7Eo3UHD1DRfpoq6FviQaCHKrjA0gbzcraifvRB2
mQ6zW0hInUfmLokZjw4SRFXsQvw3cbULxpQ1XZqFgQ9ckVrdXYX+2FnbML6Y/xou4LDkayh8nbGD
QzrPxhhFeWeXaNEadgGhEqMoiU+qKMCmJSt/KXi336CYB6gHRaIH+kDY4oh8bge91XsHffY1HXw/
h3KFLuwBAXmwBAHRgsoEkA+bwGBYFyhagmwbr/XXEUVJcqcRnunPty8o24+GC8QGW64NO1tTZSit
S3DzzlHIJz3dTbFcwOlPTQO78mF1oU6kwCzyoecGtIGizWPGBcaO2lNo47znWZdjHkRHEQ0qBMcQ
zRTbTUNh5/OlyjcRrwYhQ4FslkVn0Qth4/wwdlbY+7tE5Et4CpkcMYoMf6lVHhXneGWkV+c7nYse
MGwuhDPArCkMVIV3X3llmuFrb9H4rhebWbFs6bft+nmEN5lImhYBA1H4Qkw3B2tZPh07OMK62478
WyIE6j71L2FDjrEdQ1o2Em3lG+ybH2MKpvwNsaTEspgzxkGjXCLaWBMil53lHyjVRuYmyge57Ppj
GktQcDT9KMsQ2H/7nd6vpq1wYaOj45SJwgKTTTGB6J07Cxel8/zRjEZcdGwk/DgTZBHtjl/11H7o
5LlQ58eJnONZYVsf8/bcVI5spW/i+IjICMk4S1K49e1Vr5bLtX8xQOu7bhaePIAlXkZXp0F7k4wN
iwEGfHHl8mCcYaGJUerPTorRQ8QqOOlqvZDe5ou8Mv0xXxAMEuwCzhsfCeF2IU6DJ+RYAWXued0r
/JuKCx2mzL43GgtmP+wErFFLZtrZlNNe6bCiRVEVQBXESv49ARdzaTojpsomEgOgFLOQweGVMMam
rr0FaxDcG0pSo6mieMBlXPVkFp7GYQBYa+bNSNnkHh+APSpG2nWABdcoYgGWMM3d0IHiirfjDZcM
ofMJDRtBeEuBL921lMRkudHzla3At8wDCQonMQbugbxPlSHHRetkRyFbsCTHYamBeRngySW68EVK
QJl8YRmeSNnwBZ8PEq6BY75+MRy3ANkW30Eqyd/0uzLBfKBL+U5MB9LLlFMBnUq88fRGF1h+IjL1
b5vVMKhGfrGyTJVFC0awvZIQvU6OeaxQiElO1RoekImRrEfi6F/GIH/4lu6bR6wgFLC+VYNJjkbZ
BqsZvNxjTOIauVxe8l0/1zNtTn4PU2M0WHUppFq5QSa5shIGu21YZwEed+mC1zQtmCklfpxrAe17
kNOi3wNeaCz6Oh5lOhWVhU/jMvwaRSQRkUjDYcCU7HicdtICmVgMObObF9jiGjIltPJ1IRHRv/Lw
tVaToA99faBTlZf+jgwwQOVdoZyXylYVOLl5nxwvwI20AGCVlQEyzCkyQaFVxSJ9E/4JSb1neT6w
KPSKbiEKeHru7vuMvZjrqETSzjgxhvdpuhHPWir1PM2rfVH/r57ERne8odM+7KcMdo71guWi9rBt
cJsPXZk7K0f4wDcAjKveukiJxJaCGP5jafuNS2FldfmDN1PKTRndBnQSG/I6gN3hy+DusCT2n+4H
tQcsadaw4pzEfqGcYYdEwyO7G6h9JakQLF42RTeW5GLIiMZrODo6TXtvLLj/YaZayOOT9409Uruu
PCEXG1nfygF0QemMpRJKqGRL745minkvvJJSe9ZYOJcTTRTTCEi+7D2EAwXunfp6HTfeck4PowOz
ZDS0tPMVFcGkD7E51w+igwT1pVKs4l1m+R45lfXjLfTMKFEonRWKaaUkqcKCM4eVbedfewwI065G
de7g82bctbIrBYNfAJF1/cqbzniSfiIlsRBxhb6fs4m4EBndwlq4wLMPeOJgu20tC9SLBHOsAn5M
ah2pCV9rMu+43X0OvlHhSAOb5cuC81suPlxvX1v8QYuiCnjqPbk8aWLmUc6k7UBjNB4ouu8iJa1d
l3nX4At6UNC/irCuP5R7KG4XEIEFmw9pqjEtLCvhuCSlklaJgj1KlQ0Ttko2UQnIaCEbxYPRFnGQ
IDAMV1U0vMhpO1OOKoyxZ8yDRYgIGjL9Jz4vq043Kums7WrIkLXrN0Z0oiSg1Xtu51tH2d76Wpyd
xHl/JMbD1DJiL0NyrHz8mZa/BZeN8pDYobocEc4WW4UC11Pfq/AIr6TQJ/63v2HdWQar5tFxyGSV
1MgM1o7s0A8UPOwEn2bhUwg5J3uW2cQoY88jbE+0Tgfq5hOvxJ7vltfZG9mLst71OBiGqW1062iy
N+t+Am3QeoPftZbX24BuE6DJpZ2pACsgx/FkDGfGDBsxf35mOrgWCfztPPljQ1TrHNQo7lGXnPyR
RU4eLVdNHyHollgNCwUMbjA9JzEj5PD/J6mjo+yreu0/P/byp5iRn72VX2bclwxJEVhYqojlRKlD
5LlaFQ/e3hh5gxuc+upt7tkdRNZ0T5MuJSFoUwRYMumV3W1vR39IhsVM16Q95P+zKGJ8A+GnFEKN
HkQEvLKyS+NoJPHjfdTDehiex80f3pPmeo5PbmBsFvqBDPAWO9pNU4z41571PI3eGB07FjdPeujF
IPcVVbIsy/PE6+g4EcHli0tLRecGJGk0ZcgzdX+afgIDAGCim3fkhWCezoFdrCLS5yN7khy8sDwL
BncQ+Vv73VlzFmnxGatn/GV8jg6HxcjT6f4ThQHIjtFbIHBVzFfcD7owCz0u6IiEkzyUmTc875u0
I9j3M7Lqs/834K5+nw2l92+QAi8lgdvGk7rOuCg86829RsvSGHCzxEkdWSi+ziGlTXpbT8UhwgaF
c+ljhPGKVMM9kyIK5df5xZL1Fh7f2yF2IvBo5q4gq0vTIHJH3kN538fUqUGImOnPmjYIMh0bHQp5
3MpvMq1rtADk5X+cHvVthbV7VGGyFwz+uJkdYDbDAj714A2KDSeTKBo5DZqiUj18J3/4lvBAfk/+
1Vde8EndWdzd4hsFHzIuPxzJL86J84gSaghSBbGkhZKRoXsU57K6jGpJQvqF7+pkZX1KV+SzQYHf
hJII1uud3Li7j8jYjwYqwj/zhyUd0rzorjNhLGf/JTycvV+AeirsxB3LJZzRVeUN/BUFjArm6Hrx
D4681iugkEQsLZGMoX8+ezhxTdpE4vJSdiJ9AGbniXgkioDGsTX4TWRYJFd0bxckdpFXmfO5OFYh
86W3JtUIjcr/JC3cTMiccE2d8dAAy+ubs8h+khuZPRpqZodIhK75+ZWcUT40xd8JzQmo/MP/zTBM
SEvPLg9KfgGbeHY+O2cBP54OZb669yLGK1Svhjc5BzY7oOlemonBPsXqyfcYEyH7SNyFbeTHzXkw
7+aOxu0WbHD8mS8rR7jRIX69RfxxdaafAP+cvvQnyFuzt2JeDmvPniaxhRHQx63UqSjn+aVwvF/q
HlGMf8IRubmVbO8gPNoDdI3kXhZREqqxwwJTilcoKi2Y7PwbfljMmMUolfsgtlgDzrcYMaTA2LOW
YWJvou0SH5o/c90rKW5pDu+8jYx8v7hGhDXTedp3Ey/v3m3jn8Y7U2HuA/JPFEo2XPGEsstZaOZP
ky7iNlDuVgOvDBn6MGtzG5RMfYeUVmmnq44NGJsbqM0oofMUjhqihP1HxIdh1MQLE+Zp9fk9iMpx
0TAZK9bSDeRwiB9+WdsRrU5Z/+W25b0xY0LC+vDOFRBV669SNC7quZBuHfyqHFpkgRmBBfLyEEJf
OQkNj8WchFUtBVH6NA4u4hDVbHBUP+Je9CR+EUrhyVE+2CtJPbEAZynbds/c7Rm8FeLtAwMOj7nN
2Ur/oifBruAfaK6BIgjXq8B9Nyb6JMt3045UBUgQM7ZZMYOOkSiq/xlImeqF2dVPXxBOcRLwxRWM
XOmQ8aVFuyH07SJpixeupynprKe0NeO5AvOevYtj9pFETJKioiRDfYkGdZoTi1Q3ssMma0TLbUFH
LxrkrqmlvMJvaesuGODlZ0/XYXh4bjd3a6wiR5EzWsWu/Or5FFH8QtJh3Uq8ynXcWITTS3aBildN
oUqPrIl3GyEAcRFEqL6Ui9TwaqLx6ysL9XhQPa7ah0deuq3iwv3OHMI2QTIcaAftGpwu270gMyil
FH2227xMz+LbnBPtiEDMY27LdqnkPhWZaR40kGZpkUjj8qbeBBC0h9YAjoi/pHip6QqJTX2ZiUsb
zithz6OiNy1dRuYxEE+6qrfjUsXM05jyqRvuZJb+bWr4A23tI49TVuLrhll5uvaHn9F9t/9nYqgx
W6jIApa6Ykd/cWJ9iFXhR2eLHBw94dNNMGG4Rfnp8kpAZpI00lX2I4nKQNqHfe55NofmF+MS+GwL
CvHU+BMGnhJZvEdOXC+ytbKp8LbZ/l0Bqtw+5N5v4FrjQ5G3HhImG2Jcx4/T1eKYgQEYobZWGNW3
5nzMfQLKZ6ZewkVroxK62AyIt2T6WeIDYglmEfJDIUmPuxLnQueDTIP9rqxus70tMKDGirvwAEsA
i2zEW0CvCIRY0ost4W4k44Fvw90+enUVOOHdqbhKfYz85S8G9NiNathEP481qHgLFpAp5I2ZI/J0
Mf1w0wu5J2oPEUOJZOs612KuywX9E1fhMbIIZCiC/HaeCBr+DiuUvfPR0LbB6/G0tK2sc32PGnGI
UGIbZ6iEg1WHjXxde+4cJDvjWg6mBWIL5JyYSLiGpwyINudWywqQY2NQ2q5jqDXf7qTIVU6hiOKC
er9shnFxUzQZOeqEHQNec154jgFGT2C2a9HmggiNCiBMr1tzO1Bs/K6m2gnqF1hL98jmlK3SB/mK
Qmc7vI0BMc4hYpQsj6KmpD7yveYEi4dDSKQbwGvIqBH1XRSWR5K26UsCiB2GiC5XDdNN+00Qc1+F
itht0a8SC95rAZ/r1Bu0wQD/KI8MjN7GMAQfSMf9V6e3ucf6tOBi2UohJxvlBuk1kU9+yeDJq4pi
yOlPQ25/KZWSr5yOwAi0L2sm3/73UGKmcl6ySB/zbFUOALpZCyvDwVcYrtyZoPOUP2MFkx8+g1pq
DqhdQX7XZgn9MSob4nqs89t7bKdQEbmgxUW2VfI1rhzL42qXeZsN0QwctihpguqDC1cbaUGo26Ua
rpT+28lVQC5FRRS70Fa+o97Ulw6/rhX2yXd8d+/V80uDjOpe3TmyeRefLHTPApKqDdoqtAR5dkxq
5nPFSGp2GMk9zNIlfhdnaKVsjOEG5YtPLNHB6uqg1/faPhramLaYUvd3kwMtz/bL1zvI/LpuvYlt
3CriSJ/U5WMZSKw94KC26YUdnhkxExd60qIuV5zjw/wjZmCY13p9jz3iUBGGLhN2PHd0g5ek69G4
as1wrysUo8YUMyd6qeyGWkmA7pbKrjtTQ3bNUHe+A3uaxrLlh8blx75S3LRIEBf9Cxs9l9L+PsLo
5/8AcmyFfAE5Gs6kuEeCKNc0Kw4m2gLAZ8q3MCvwcyiX8qUjgKkW4qTofjmnZ8XF5IjdYo7RRP44
+DHw8hQRVfnrX0Yv1sjA12+L9A9Mfl8DVoerqtIXL4hISwP1udfdeEbTPjc/60cI1YMzsymciR5N
O+qIVsYYL35/c0/WIKA88RgEVhkEzaSaz4fq8cKmC/9wtyGM3tsqiBVIayqm73z3Mlj8BRpf0g+q
chbVozdcaZnQR4sE4U64xpTCHJD4CrCfnCyRcJhOm7lUnDD/WpNBacVofC9UkAJlMGDpLcgfyeOM
ftCvezdT5LLInIYGT5Xp5ZVtJsvudvCwtdI/Qs0pKEHeXpOAvwXt7DMfpjkyM/TpqHhKeMAnmp11
2LOzaXet4nkn7WlGRoqtnDrMwkrBaIv9uVnLiRTB8oEJs1iyxrczmJYQ0v2vV5WgnOcOPlZQNrJN
o7Yq2XlMzTe5TsjuVz5aOp2cignsJB6cIuhmm8tfaT/QkBWKK9rJ3osOy7eqGLpswfASNv2/D/pR
yXOKsWeo29aNsl9BNvD50jiRryD9+mngJh2lmYj+vn+8Z1J7QmEZjn5nwjiAJmYWMqaT2wglPacO
msX8A/3L2ngoPVCdEi2vaar6yyBC5j/9HOrPrc+VGVs4mStUpCTKcWE1wFe3AYNpFhhfXq6saU0Z
k0zY6l6rbsafXnFVq3Uusxt6B0uo7UbaaJQRtm3wpXPt9V/yqncb7xN9HqhcnXvvlX0AnUPAEyCO
SWcCDyEmVSApQEC6uWk+Ko2aJGkdIVXylh7QJnZAcC3pIoRWO0iC6VJ32O6zxHFDMpbSRXuQ3HwJ
WTofO+WKbRnffj2a5xwBK81wLOn7tHtIwdDr77A5yahI3xsGu2e7Fq5437bMjl5aumOOuajr3YjU
hnzgxKnIEzMseUVx0EnYV0H1/OMF6UYRw90wzOtbwOoFNfIM+sm7wMAL9EjqSXDwiSwc9hdJsPIT
6vwW1W3KpwAOp0p+84bPx72fn1r2Dz+6YNZe+oazotzI4qzYlONxRf3IHBXbg1xU/GMSOkhBTc3U
8H9Hh0Qu2shV8arNhGBxSipuB1LKfU+9c3VssSlqCQJd/y7iydlg+F+m9gbvaWRsK+5l1VITecmg
WYLcOWNyVT0D+gQdb8luiiyNSxK5us3UbvINWNd6tSueKPgj3DPjOldyWfFRLnnDpUI/0/66JTBD
6tgZazSun+Ysk0w9OdiOJXCZ0/O/cqiWmir7mHGxxWsQqJd6OWUCi3PIi7boIJxoE7xyGmZZspW6
1OJSEK/CofBfGhsOI0k4ikbWziQEhIh+DpHUKC0M1tAkmzgAMjePP/C3D5xRxMLn+IbSZlFDnJUs
fmVgo9Ig5IMtcWICoyU/SGnv87JbF0H3BIbBixnxw9mVAjkGHftwL/AImK/0EvY0SJzBw33OGP4I
fVVLP2DAghGXjQkmP+oAqLZOPqlV8zK1j72CO6mC/LQwAJq59S7zuwYxXQYKmwgoadoco6vo5f6m
5lZxv1uqNFFQYhZOnwLnTDgUWLzySVSr+p8H2fbDyqQKZv5yh7hpVIC316KjU1iKXidtJI9z6zhR
TQlCVM1WlS7xei+MUk+LrrVQucxauz783sEHne2TDLBpg46eWpeWzMfgX0tHFfSRTNI0mmdz1S3n
SW8j5j/QUeWZcZ0XASzD1rqtWqaRgwUbqtMaJ55LqYn+8jExd0JNzQH6LYmzGlYtOM66LpjZarLV
yfm5cNorr8RdoiJFX3PU0SHWe8DkylxGcuQrMqjWwJ3FMgFqpNWHOQRkDDLGgheTX2eJ07jPPKRC
BZEFjmGI9Mm47WjrRmbsHRHQtg684yBB3Pj2MRzSdisYcK7w3SMumYJwc917alaW9F3HXgJTf4wX
3exIVXiHfr1E14FGhizv8VFc1B67qig/AEWSFQ5jSaK3+RkqlrH+S/UQEEH+3R81RgEaQKHM1vzF
p+ZPUq2CoAdK1ZHZ2Wbxq4zi2LvXDvH3M9NZosip6GSVUEeyriDPE3oViJDZStCJBciIoudnjZVh
q7Q9ZAB7yqj5AlBxO51f9x+FdPjmItdxN4k/a1Dbd6/2MvTQdXuEKuEoo8wN84C4xA+qc+O8sQsp
TAvkSAVMkypBQ6Gyc3OoGJXeATH9E28ZZKOd0xJAhgBQln7rO6KQOuw5xzSBBfuJ0k/edvOulnPf
FLh4mhxk6o97vqsCh0udF2DD5BMpJMw82AsajwbErDUxRLNMsnj0kZ+3Sru8ki0Oh1rHVRc2rfXY
fDH/Ro2SfqmHbWjFHe8goJp62psF/9IofdfiXp3hA6cQg8iakKEAm/Vr4QWJLdMEt/Xs8p146Yc0
ZzDUV/I7ggu+CawizyXqmSF0B3BV54dnpmfKs3yYy2dYct4lTo6f5x8VPkWPv8wKOwRFeDbJGXdn
MMJo/B8bAAqE/sDUm5Swqi+YvlVWVsP3sW+Dt5c2dq/iMUbV/iLx1Q1pRTkOg6hDM9MbSbVG5IcZ
V/q45xASzjxQUC1yzbR8telFGten5B9krzknAyrQi7Y5XIznHcUJJlzONEs2sWeJfowJCL+dWdwM
nrnJlZ+hYjUOqIWNTgNPc4kVpglpCQLxEFmRzSVhIVAJQLNeS9pwc/hh94CtTPoPd2Zx7e0YXc2R
7vZgkFqqT331S2AByDAzBLveTF67WjR0Fm3p8ZvqUnmK9PeQd8pPOAT+NEy1JK+4Ls7iEdCU20GN
hknz3QyUU1TlP2IVNb3zljXCB2uc5+9s/V7J/XmfoPlNOHYQhO3H735PURkbHuick3OPloDw+EP3
vGTCa6Zv2DMnFOMWDPVuJh0PpBio1YMvNbCE1HGahZGzuyCNqr2VBJ+px9vMkwN6Qvr0M1PI3yjD
vS+jPpGTR2eiaVpPxe40pg5tnL5y1PwOy2nA0SeEA5MSMvyKnrOaP6acVGIC4bD1eRw8heZPIss3
Nz7RENa6w90C8pcqZtJITeRl4JNpnhYAzqjMwq1xfPWyKBd3TiUqw3iWkmy8qnv41xNMK8RedAIC
/fMckDw7XYv81Dfef/8QtQ7iIiTSs0Mafl4XGNnNtvbrS+F0MNN5Ef0JqDga94If9qqR5fHqInZT
fp4ssTqQxMFkzab7sacZ5IBBfQ+LPeq+kdNHOkazKNf0nVtVRDci5Vlv2DWY1MPDwuv86wog00fc
vCviV4IJM6G7hsSyVWkCOfQs1TmGLNzRGarK384+Pd51o4blv0eQ2ZGmTdOlXeshAnKcmKJkfh/e
zpPpvWEZZJTGNdSPthqdjLMgXMY+GNkgXBx6CXzyRml2U6OPiKPhf1IFgtP5veaw8fHkdd5nETfM
NBJ5UCiWyYdNVg1lr1RMbm0X1of18BqXc/nCwIktjpe30NpAjmEht3a/HJ72UiqtM1ZJU05OuHg2
elACa68nPe+Zr8fVCFvmb1A2lZsGi8D6fviFv4BEiy/Z03TkxUk5uSpVRJ56SiRzsNIh4wml47rv
B2diRU88rR0kmx5Ow5khEEDxj27FqrDxXevujJpVlztLZJLTgtbVBaPsYYbW0OsT72ttlzir70uc
FpnNKn9SMg0rg1+Czv3EIa5TkHMU2ICh8l0oUJZ4MwiXqq4Xs1E8fVUPlvk+qetQwoyPI5U16FzR
+vmxJjAznmxXBm4YgDX5vFU1T9N6DUYkEGGLobOHVSJt2pHRSbPJq/PZWDHG0iLwMYtEMoEWnX7v
sP8N6LCNxUb96+4VbjRA04THX9ze8z/rVa5RihSkBYh4WE+RqQtNBoiN/Ex5LSOYjOWX8WNoDmaU
ZuzB9sJgQnkUcx09fvlAj2PPlOOzXLkrnCX3zMKpLq0Broni5n99hR2LWs7es6rIgvMA3EDpyQm9
U2Tu43gglxziVBHJJ2vNOBD0mf4bVqvP30nQiGVJSOs4NqtFJ86Qx65/fZshneXxvsucYTUxlDF+
9kclBnI2sQTTxxm6GQ6fkz2kfC6SLjyu9x1BG1a2mJmKcC9qBmfATM5a7F6N682snUflNMiRjIMH
NRDN7zlbtj7vZWQQZXHJOGNc/8A1Q82jD7TpjA3IYz4a5O6rhBc+Tj5JM7T+TxxT7HoXysly74lR
67/6/QKqWeF8CHa0DRSQopRgk0GlZYOQA/t+lG/9oMg3a8XFQLiMjaooeLS/hcfjngPmTGRlgTX7
nlfPnUsmAc5nMLm/e3JEi1/ue5UVIUlS9faNFiunwvAR+oVyhDdrjJhGsblEGmvmH9iQ1n/IPqFi
1u/upe31lZ5/qT1nz6QDlo2L4+bn4bO5Ifsvv04O1jiCwQBFtr8PCFGJyAbcojcWMMDd6+Zg2A8K
Hjwrs/6Qc8IhU31c72IppjGt/e8qyvQeEXMdtVxc9X3771683xBfXE4CNHbaQAvzL6z7k0fo3nFU
uXazgaBEl6/+ppkLgibSkTtI6XvLGxPxEz8A6rP3ch65583f92QnBalVBA3iaal+ZBbg5EeIySzP
oxra+sexmYst8uw2041rv6sxOkja/s5tm8VjQqVmJHu7yA6TIAUDGe9AtAw91zZ785Ok+2S0DEmb
Kg636uUD75GNDrEbuHlcu7YOHTwZmkAWpmRxg7iAeX1SeWA5twJTDuL3myE7pohqraMUlF0SpUAX
D7Ny2JEi36oPTQ47WS9eBqiZCjxT35Y64pe/6ipZJ5ZT8gJ8GMfm6+/8wC3QJpOd7xr3ct1jgs3y
wvuP6RP6jZndGM7/mEji5iBO43ypso5CqpQOs3Hy4K80OgczKn5tePrztkcYsIgKmKBDR7ONdVSr
F9JTepyCcnRy3e/P7huwsN6TPM80fbwULnnuXzDh7GFnbxpVi7lP2y4KRNakrmEZWhmACMit4Ex+
csPMSEI1TMAMo0BnMxPhcAh+uhuEuSvUpEkgwYe5pHZldxeQPdKfBMOU+uf3D+i4ROwklezGLRWV
Y+pWn1Ubz0GxQeytJJ/sHRxQvhKD1Db3IJJXh23GfCQJFOLJlD5JhSQ99k/DuW1rUa2CKqgOi/lr
v4BHHS4QE8pRg36kZUGFEpTmtDTi5C9iirZCFO+lRdfsy/rylwldFNZ+0IHRYM1wyv+571sv0sJu
VAPK4X3SfR27s0wZqQJqT9g4zQ8S4/61jbluLTTO2LPwUFpQVFTAHHNu6rdDxQ+nSY5opQ/oDOoQ
qtbtPts7HhjRfjOIvNb5ELeffQi1EcH+2tYtK9kyIa951Rpj6VppdZo+RqQwZUgg3qEavmVpUojr
KlXEzRXfwFcF/hxZTHEZbLjB1CdN3bUS1Bt2LEmWvDFiLTGr8CmbqEgx86Gutcc6D+x9Aiv5vJ0I
60YlGs6iOOLlRLnGAUvKmp6eCIqVI168Tsr4zEYNa870h6Hq3wEhqJLzvGvRuCvD6ccCoW+K3YAc
rlNo55LT+y0vkE/n9edIUYdn8XIit9wLaXL4NRz99VoBcG9GWeHxRKhGFfbez30+HzSgCJyjxPKm
wLfmyyuZuM+Pfr9zHB3kEDr6EdC8aWVcUumpe35yQB55kqFqTur4amkWBEYJxrOy57q7aoB+yMsY
INJlaal7AIDr6L/Jh0vC0ljgh1Jzis6w0QYVoN2fXtJ48ScUX0IGpxXkY9GcGkf2F5rhFsvFbGAf
QhBq+ppeQyAS+XL27/focvbl69MiEAXsWIrKkDoJR2m11xsrjpMCZ/AyNURFmA+2SQPcv2YjICxZ
n5huahXMMFMeHUCY/dokGkHEybWKa+jCY/ovKrKZlcb9myOeiGnFBoNsnXebB8qva1YDUXjcgHW4
PkK6LXXqQQ6DFrll3O0fgUwNXwvpx5i9ODuiuiduQ7A0JtuTJTtEhInlXjcvpYb8OiznuDrNv378
MMyK1nOKauVp1O831w/Pjv8IUFfw4X17gHANWPAYR6qmL417HPLH8kG/xumOZbwP0ARgSk79jO26
j8vcAgO9vnDI5V2OWtLAUwIznAc7IUfsEz4SY6U7xm4K8XjDSJ5UeoxyrvSTO9/ZuPTO9xspcL6L
6izI7POLddBHWZpQZ3VI0wORFdNXPV3AdRmySv7B+BPQqPSKXmDRTemr2taTet8TGa7uGtdX+Bx1
BsiiWtoJRFq8nxrT59xOJdPGuRHfvIIuojME+B+zyFAejxUK90dikH3Gn5GSvuwqKm/bp4dBMA3J
D7SGLsqiiqJ6eaNlpmZvtF9nZu+hJtViU70edhirCJw0YK4S03eY63+0sIBvit/99EylVnfwFBjL
VCby+RSdQIr/FfcuCEYSXp6NWmY+xHSRnm+dtzwkWOyI+LM6p9ZAB6y3BU11e0gULkAmdhkuGyvL
Hu8/NiCfVCU16fnit9KA5QOWG4CIvF9mv882+EoMgW1yDUyOBpMOlma8JSfLV+iRouWdEnZzMcf7
vtlMAWPKNbs3ooruUr/qI9IQwZX7/g0RDkoTKnC4zWdAZfjk2B2kuS/OKYsgtvseiQ2n/6K97YyO
IofOW3g8JWbVPGpCA762ONBIdt1OYJA/ZlSOUqCalRJqUKRlmyeH+ZRLWAF5m5GYu118210IpTqL
lSFZg0dlMuJMj5MqEVXE2FMyrttuhRKKrIoksU+QgjfD++ZR53qeaPR9CHROLlmEHn3DDbNAKe0q
aVJV/9HuCiNkKhJYGzxNVKk32a9MbeT17iXcmzcNcwjz5Y8NerEXPnyh2l1q38irUd+KbJpaLF1L
DgFgQJThbJXJYRn1v33yHC4IMUtDeUcVYej10LKi6U4vgSvfU6Oxut2VErVjHqFnkbWQJ2rC4TVU
2M28NSSGLIT6YSfrEI8dleBvoVAo2IMtLv1kHYf1zd9A/IHZYcAaBcgDQb9e/qNXWm0SgL0p+kiS
gDTe/osElzL7auw5VQqtKnRJoC/P3TOxOBU/EVWf95Z+PMilfGctwjD4K137EjsfolqpntHLLQak
vmvQ+ywDSO8S1VoMDSN7svmr3NSg7teDpveRcXOl/SkrHYRiVkKVZSGJt6fyvKLEiZfAoPi4BYKS
ShD5U/c2Z3TcrceGeejzsELFQzc7oKHKLUZc2RSQDeet0Pgj5QkxSQnk2zZeW3as4Yq6wwjF3Zim
J0INbhHRTbOEYa4NCPec11ZWozu6vBYDXyov7j+SXnyDURNM1nCob3fL9Ict6Qu6siN/jG9efLbw
xXhnX6xR2ohRenUreF+iTx0a+AEV5IMI5CIWbpRKCk9UOVcgrkiFqpKaYeihC/nfQ1YODJJpEqgX
pVEqNvQae77LwiANMjiRXTyNEYX+g9IFPu2Fj9itHVcOwsmQ+W+2VnAJGZoVnHmjavF0hUBViBMt
22cETBIUWjT/A79PcIYBNBSrJ1z0GoTc878pJBrzp//nBGWaQ0uVV0bQKLiXJNAzS4KpP1CcQWyM
BBOtjZHyiEIlHTNn+C6An7/dBK/AXG+9zeEbPEGPNVR2NRs4Y5wi8zXM+Y74D8KGNOtxtbX6w20v
+xZ6K3dUTMTtNa7hluKwvkxS+Pu0c+xa42jJxzBM7NsRvsvC+guo2Jl7cPDhCEQQ4+G5cu/hWFX7
2SoA5o0oPZvChynaZb+AynT2NJwUzUHVEkFI7hQoY5WTOnxkwAkczWYPNe3LpM94TdsEdRoU6ihU
BrUPbuhrJBn8i1OvZ5d36Dvkwjz1VbKCjaPxZ4PuT/bRMg0agPT1DSoeCO5C17eyCX0jxt097ZFA
e7EQ43Rw4Dld3kgZosBL9rWfsw9aUFpYTBMrKcS5FkHIpprsAO3UDDyMI9kA2UpKDvCbnhuEltAS
tPli8KwTjZq6eHk08etaPVSrqRZm6PcltTMLWErgyWZ7q1KNS/mNvcfoXmP6rZcOgv/CETbw8bPI
DKGhxJnAvQIS2qygyUMaOmOic0hHd0AM9f+V/0JIDFbHjgm6xKhEN3H+3MmVsU5a4JgK9QLnVhM0
TYcrZi0NuD2eKBvOlTgXffQIzJVoh1Q0g/6TK2COep+bLHsVRF/J+9d1NwhrsrMHZ3iiM7iYtPQW
1kpqnZ0DNLk/avo1rpcG/2yuOpnkPtXL515twkUE1XTeE+GlTD33G85AaMY0P5i2gpfqq55yyved
RkZcSwfEN+GOziZFMh4K0KXC8/Gk3wRNb3cb/sI+dWtkn7GDyXxuPg8JIDum/CcEA+SH8hA2kKWP
MFUiiBxKfOpanJsNulhQ9P9TiwQa9l79zWVZCyU9V07/NZMd987DZ5jtRfJhkXXjrVH5oPFzzDdc
+ej+Zj1+ZcTkLW1HpRzo/OWU9AnjZ0CHdv/gC6k9O6hk97aWkkKfV4Ng0x376hSOtZOpYMxVGD/S
ljlzxBt0t3tqdX70a8uUMHPsvbwuPkmSSQdinjCb4LttYy0us9YguICXYV+3dhdb2buqxfemQ75M
AmxUlCKepCMSIbv0D1mMxMPHwokWoYDHX6Mg7JHoUCmBXm0J6MviJFCDGbCYKnXAqmtjGJg/QQuG
P2eKEr5+MqcPVNZt3fUYn/NzMiuTtENoebvwezWIV1/vChBHC+9CUmsgg9oJtKI9MUXBk8J1cQOt
2IK7cT1ndhDH4yam9YyONeQRCLqJ+MvxC8+1gVdOyFFfjVNE1iJ0zmw+MIz7WJINbSSPiTCckNJI
L6uhVKrFy8ToNEDp5ZeRgrd4B6co7lqJ5lPIY5G2e+X4M+8Mh1UcZixwIV/SOCRdb2Xffnmxrdw4
C2BmCTgmNr+N9Cp5jURjQjrKSuxeO1fLkxSgrGiO2vGPLEz5rIQ8P6eCVuUBuV5fqjNp1lKecXp9
mgiPj0Ie1spVcvZcaivDtGDDjh618CiPIbUzXVe3EaCZ7yDmf9gjR8JCRSbqxXMBlS7xD4W2Fuuy
iFBDVsrgw87kxCPKU+i1Anv6pMYMHu2/XDzZ3A3oRrhFEcctU/2loG5GUOnKGwi2CSPbDuZ5nBTg
zvo/eVlLJfNE+hQ1GTCREdrOLmAt0ZYqFRkfHiNAEyIc1U1h7VJjia4oFHnOzhzwai/bFIVyo2PO
7pvazOt/aLxEz8crRWFkUuPM/H0raYtQF0K5kWHRCKdpXb6O8tWXGgjDfsYE7vVFBCCKj5AkLhzE
7xUi+gjuQv2btD9eFFE7UzKh9Wu/ru5OXQ+0FeKbsE95Qp0S5xJV9RG3QDEYbzAbA1BsQYODF8Te
QWrUiATZGzHp6GnogOIq1IxZzK6zTz/WPGmJLKOl92s8dhFbraJd8wJdyjqPF0bO6v33oHAc0Uqs
SgS/8hxk6jBYWJbEcYiG9COBb1rCfwr7j55Aoh6ZJACoNFXd8Mbh2QutoYyD8omYLsfxtWgqQ2cz
rDid0y0WQooVAQSomodUhkxU0UdIqKaS3DE/IZDuLgcy9IUjI/J4Sbu3s5uukC2f7YK4Juj7Za4E
zNkgB2zSOSDooZgPnto9960fNEdWLEHWRTrjGvJT4OUCAIhjD3CFJCCPTWAJoLIuJDMbaJa2IPUU
8wxlM8BhClIw3HtBrEtHPPNic1YC7+BYqJP0FPtA0l+/2yAhdOF8TcuSQShbqUbY2fDlUgjTw+gs
dwXUwv8QNoJiBdrRjCRh0FdVnK7fMrERduhMvtRkrU5LQQPf/FT+lvk96tj7Rh1tx7f+Couc8Wxp
hkcm8UBC31RZHgPhVdX6SawKHWVdFWtDj1eymOusFHhJBGWPRAPdMNcOAcAuPmtSZGRroi50cCkI
LFpNKqSpLtYpzGlCKCQ818HFdf4s2ZvV/t/bzjfcjQBTnRPfbprvdUnSOgfEy/WjPA+XR3wEfTIE
6GtmPya47T5+QU86sXYGdeIInQqqn9v/xDU+TL5MSi64tnJVOcplvSSgCNOKm0IkiSJ4fTymmFy9
/MHXdIdYbV2e1HrtVRl88WLAHiuP97PHme0v7fzZ5fVGpFLU5XVgtQBmLq1s9CPOTYq21axBLBj8
hcUUuKom9utV3fGEAd4dEvTkRDYfkLiqcK4songpUVoaJg1ZnuP+ls9TU2nXFO4r07Bo/rTgRAzm
C1XCKrFILOrtFSrOaNI7N7lrV/CHNm5Yxckrh23+uiavV5uzIZhFzYZedKuzMepbt+KWVkLmKGPb
SYLkAdjXs6P9E+1kdto1y09zi5gWbHps8cK767/JamjI00ZDDK9nFVbJmCrmX0vqZpHpxhlCFUp4
gEblULZCy1J1Lcem8dNI9HNcHHsoIPT9sjtpQnj81eHkfo6rsSjPeyuIqMFrIiY455+aS6jdVQ5/
273ofo8lhlWnbQMf2wAm5KSkVnyBXdCmvScoBKlBvGR4S0a/EPIh7yCRp0yINKSWPDS0KS/57XSe
3/rmJMjr2dUZV57MIT/AF8hlghWO09PEYAdo4IRiA0kANV97WfiypDE8HySo+ZJ4zdScSskVyDi8
4WsctrvsZIaAZGYTg2QAZJnR7DXgPDBQU+2IjRF0ky8MDAY3TiihafY/FDmYV6H4UdUE/VfaSGwZ
Efs3sUne+OFIhzY5z+AbLdvBIMvPMGslhujIoYsQ/SWQsogsTC13lVTJUreMdPwhxVK8L0UkCS+I
GRO9uugNANsKIs3zRzpre9OnKIFdZRZ8v6+IFFkuZmm92SNuqR8AJOhtC5NhHj//8+yszzOUgKJN
gFoi4MzEKLYF5Tc9dVfTFuzXVcP6QzMBEAjvvIrK8GcRoD0+Fabq68cjmmmtHQcq3ZkahR6undT5
THprTU45ML1+mk3OX9Sc+hJMAICR9jn0pKfleFOw48uLzAqdFQuGY0OOJDVz6Cv8kdvx4sJDLBGI
v/pI4w359ntQ3xCqs1WGG8nMmDSHZ5wngcphzgd1dV8+K2R+KhioiVCDyVyNKdD923196jkSdn5d
OBn/SdILFVwVGiUUUA6HcWh2LOo5W3bBHFrUe0FenGHmawZAE+t1DilA4dih/dMCvAwiYG+486TS
5VzdjGad+uo6JgRsZ1zrJFe/jKNiVkJs6lui7t8W5tyRI/sbUQKcFiJdL2bWBUSmKc4DhrbVgAGf
OymYRgs8mdsZVVuM54yzVI+V6NqxwnpPutKICFC32l3c8wXyZ9Zft0isGvyyn6izWK6B56+dqBfS
AHqKNt+Fb92HNvirPKunr5o3BTC9neGpuprka7kHaCt/PSFXp4VQHaNi0dEvFAp0N3abQ5eLhHgh
He9yE7vROrhmgKGwgjB3APist0wsPVA04bxKQEW9AA7XOsQaWj9AldoiVoNfKN2uOD+OTD6s9GXM
v5Q75SufnugMrepbz467KpzwwWNz9QIo0nW7d8HitjP7w3n0Zpg/hDWkXOGa+7Qe8ntq7vDCEaoQ
b7EcLYecbokkMsPBlx4P/F8yqwt+c4ebWtcQrdBbMscIuCia9RFVPacMblLqb24O6yjXZ6wwVZsa
BEsPCThHM3694BDOKHqUfGkM5Ks9SIlwWAgPraEEgBq4fVEme39aag40pGUrGTBECjJNgD1m+tyW
VbLkJS+23Ln4kNNNWwbsVje+b+FkZ/83iCQlODfYOQodbNTbkcNelfzARffhvKlm7oJQ2yRQcBtT
5KHDCEBEaWvOmJIuICl1yznl244hEEG4XC44baZ5KvO1O9vU2iBuKqV7Yef4eRWvc0DehJFA3ox3
6AUrMIWHMq/lOPlFGLh2jiM90O2D68GToPKnWBswUxzdLXi+MGXvWDzsiThmU/rddZJJW1uVD22+
TNEcFpzVoixC2EhDzgMoq1R0bOyXCOBioI/R91qdAZHG/RWi0I651OU1BxeVFgK+KtFs8gZBXavb
gXjd7BWoC8ssksUgLCbigupkhFfP3issX+BxFxFoMbP3O1Wl1gcAHIf+Pv9dZLmQW7inZLxA02YL
7UrYI/R9uJStyOAQblKwpRsgG5zco5mNnw0ge7flacWV1Bx3f5FYhu41mZcjPQDsb5SLYTxzvM8r
8RSygQo5O2eVABupoPyxZzPbcDLQdrtFCnJedcxfuvu/g61ljWSQ7ZX4OwReBqMKMZRA35NGTmCU
KjFq5Ot54EIv9xlr/Kyz0NRzdEh7DXkXtWq0hUcTbBTmEuLxsf19HpRXmOrrFMd3+HHrwkoHSbeW
WG2ROYrXxoQG3omXc6V1ddOASne7HhU7ZnLJhhGFsS9+Jeh+52MkrkUgO4WF+9lyP+2GNPUVmX9V
/eTZKVJTeCookZy3pViK8ot1W3mrtKLfQ6l2LUBdU9EK+ZToc0Vo3QDDOGas3OwC9TDW/IND2MYR
LLUPwsbFTM6HHW3+/Os9RvdjnlVJpXVIOAQaQiVRGkQM519d5NKRonOkE64uW1wce7bq6lTyBvg8
7M3aO1EI0GBbhg+Bj09K6EFhPgEhbdSoj4noO5E0WPvChDnstkSG2HW2E8ynMreWJnh6Y/1fQQCN
cADGunsN9u5tI4U6RdsvYYPpgDz4b+cGIx8qf65mZcA8e5cHhE2OFXPnXRMrb1C3d5l08QMrEbzE
+2JquP+WPDgOvFbly8ZA9ZEkbZYGFWhAJpPnIKAD3BpeVrii6cDHnCQxiC8dKmsahgirWIMqd1EE
gNUYp9ZOl/EutRI9+MhAFj9Y7DdJtJPguryBI5fbgGgx2HRLo4jQlN1ztWNGRhqSR8rHDpwa75hK
w+oq/8ESoJ0iFiBCIZDSxK8ze2aw5cXrC5YW6ssNxFKi9QpJZ4ogYygRKl6PJbR7iW3XLB9zmc7I
y4gHyQb8zzFSyVYML2AAgJydCNyJXrWgaUfjOApJL9wNmORSZVzM23dciAyxomxOoIGkHy6seaZV
QNUhBfGqrjkgPfaIHzXc+uK9Kqu6Pnse6HwTjAPf9LD45+Mfy3iZV2oMWagUh6dupp27isOU7H+o
kF756QflYhdfhX1qXG7qhz1OH+ck0hoUHFOUlziFb/t1aEYCHxTXMiBbxOcU1G10ctIroAKeRN56
RYYjIIvM+uVyx1fPPWT/619HUGvLejYjb7Hvx0n1SbqkLiWtAXr1QmQuWkNBSTaxrEl27qS+OTH1
FpKj0Fpn5OIKSBmkokQLwE73wmBCtu9LS8goohU6aouMuP0eu16aBzRnJQMCiPCoY+x8IZvvc5m7
zsom21ZJ/leISijpvQWB/cslP3nnkHLD5gfpUc9S7cLB/y1twOrfrGER9/bb8pE6XgD3HZOdtRZt
hoyDw8WsK2BYDcLbcA30qfgcI/NlxGYBh5X2rv+FqC48HNOTnUg2W3EdxT8l58v17zh0Qe6SKLsB
uyMW9C+Tv/fSgrFu0XAQSA6HXoHcQgJuBzQez5ey67tMs3qPznG5KMGx05hTMjzJLOr+zEN4uhKZ
tiJbBCPKOBg5JCg2+CMAEVYkYEzgkyu6i4NyZvl+awKio1l/DnD/j6owoKU45tWJ/13Ui9+Sr3Or
89BMCgzJHt5R6s6qP8K1hV57RzfCVjsYmkMHoNIiCDbvKEVAPlnBUjhdo45ZFSjuAkSc9x6ojT8h
mVVSN/8T0i/dtQdThw4csJBbsCyc5L9PeoQXXKfJckcjylgdRHXF31tORHrJmnMrVqx27z27NwaV
7Nop6ijOFizv2sXPENdiJn5CRGls7abKma6CKghiIGuFmRday5h3tsv9SZhXm175a0/kKk5775MT
xyMJCe6H1uondFEHmcs8acqV2daCESXLWkFOkt91kM4WPpnNRvqT9HbLjwwluqQcLNmepUPhfVhA
WPeQQZZiR7/BDpZXyQhPljRbPDsweXwRpGjxOyMcFzAhkSGmPQ+bz5KFzax4E551RYHJDIqJsJ4s
ZTk+LvdVjxoKXMGwgFPNA6IBndBLOuWxxdlzwayWsw8ginibgg6icB01v8p3R49HlJRJuexICAVV
38na2DaEbberxXD6MIXhp1Ar6y/zX8dULDoFI8ojUehrY3xu0hysQjwBoCs7xo1Fpad7lf7TKT0x
kBiLBSUj3VRHSfbqcRVibWWEHq7vXhnBmcX/zZmO+EuqK7WJz90h5FBLQPQ3wmCGSZj56l9WH5YB
VBxyerA802igiV2hiR+Xy8qsotKt9v5EY859IsNVZGS8H17p/iko6zboQg2++Fz/bKU6LQJFRAGs
Eki2r1XiNrN1qBKLREy0FoIIVUSBLyMGIK0YXCKdu3fgBw9Mpfh2DhC3H/WRitWT9kU0hsHhTspg
djWlp5rP8pqhP8NO9T1OkjflY6Vua8yWGuSN7wOpbLknkDAwjOOrJmM6vZSTuOaFQGQodWl9l73D
3gkIPf5RB7mHABeLTzy1A0pWNW1sIoMOwLLcjkLL2k9UewRbKzsP8ESmOhHVSFYU0I0fxHMKfzny
yItqPFda5AeE9yBahqT5fxQde22QuL9e6Lj5tCk7YvTrJHuDjVNhTFJIMDbedd4NEo2nw2RGALPj
7f4F+uwwJ4EFuaiRxnNcipP2ZQ8y+dalFHAv6YEfDxhVzXHO7aMtO/i/ljwuR/3yjP9SorsN4xe3
CVXdwgxsDCg+bbWTolXxhe5YiFykoZPqTOg8LsuewTiM/H0VGvnX7tBJvtYGC/DLAhv4W/XwhKK6
SBrvAMYAPr0cdUkOXxF+BZfBddC0M8Ah7hQVCXn9FGdtH57nLNNjtu8FMYeZ38dhMocI6JvlFG5a
304YLw9ccP1VfK5VnVtKon+H09K0FWUMx5Nla4g/Z+X+Lo/1DGtFp2fgQd2hqmCLZl7ZZVLASiuW
EqTJ1sSAAamN4Fc9M0dolT0dAoP4spUOaxM+WELpjxgMjPQ/OrPgx3KXttdt4/YSCFJt1cbGVX7S
qG+9r4uk6GV8Z+9ce1SsII89/E/6fxfFbQdudApZdoWWIvEgT9dXR/Ej+kaJPhmc0MvJAluENMKM
JHRB3czkMDOo7lOY8xuBWs+An935cDKIsEUpUaECvK3mAMbaI+voEmug8dBuyxmAAaOrVDfbeBGi
a+apLS6L0kvf800Lp797Lcl3S6sQnaZRy976qHcTytggWmX4ghqBPvHARCwvcPlrSln9LL7hLw5F
Iq2R4DA4wxsjp3y5eKgi2C7IbIhUHJxNyV+W6u5xIRQotAKPc4/KhKaawqzTFJDwBgmdcX+m6xNc
aFPgTxv6Pl/y6uaayWdyrpM7VwHNIrth+smOWNhecLUmaxjtYE4Ueyicf0FvkWRAqFCmVZPTNddh
B+QiKz7NWeovSPOOmdxy5PHCGgR0282O8jWX1UA+tmpVzkBw2scrtwGk9E1fVqAsT808+su++8V+
Tl++SgpIvyb4QHVYxCSYD0gA13tLL6E09nbC745OGvDB30oxMfaXoMEy6uihI7KO7L526pr9Sx9Y
pRsj9+5LXjJH73d8d027uMM8uXC8OSkudEux2QwplDH9rBCCPrp0viBQVukQO88tzLIt/3Mioypp
wzod5sfd91rJTm40JbiFxIa9nyBDPAoX1CWp3prhtc8D+2TiiAuLhZKRfGFgd87asMd0mYtnVz+o
zuAf8HsRXnQRzvZhAvJQQVWvzpt6FCG7L+psXu53oEYbcsGi7G7C8dNQusdvoaxMj3B0xrfhR2NQ
h+dui54yi9C51Sq3rNot92lS73oVv/e/rfMx5mhSjXewmhE0V/guROsUaLdH6t3VE0BhV1F3Szp6
3mLiR8HB10PjK5cBkhqHXW+Wwr68KzYhdCxMqxKYQvwwgdMASf8krULa2SCIBbBl7HmxRbb5vQ60
iZs3CGO7vU3/fSSdaokzlvtN6Qx7prEYLyUNnIon2tHxlQX3Cp+VUWBXlYWADjNkRMZMjEXnd+yE
yQdiAbSVRhCZhTKIWdxzosqX6g5GhM56ShhZiyvSTWuGHKvN6dSaf42TxSFqVeloF8vCgj+wVABO
JtuB9Ww5zcgSB8kAkfadqaOqb1sBd2JO9fm8YqoBfFJdSoaJiES2nmq6mD7Oky3Tcqr+5YmblGxo
6DOE3wwbHu/2AvNtSX/pTJ8ZdLTpdyL/MWB+TtVc7IXwVyTn8YJmZ+LIgif/0ovDn1XwR4wZYphK
COC1UP3rhrSv1NVS2OtUCTi6yZV+ObAYp19oLikGG9U9tmuxOm5/YpjyWpIT1f832bA3Md8JyS5A
nVDp3n2MGzZbVVEZSgSBo40Q9aXK/1VhmhkvLJ8o4ew9hC99Cx6ecDkfizZq68BMXW7GTU3IKeet
s/QqTqT4XcGLAxQARoKoefhNr5lSDJsI/5tovNkIfVOnXw02Zh86k96SR18iHPPT4Cw4DojDt5dE
RWZU0fLC+ooly1CpQa6X+eIhAaWe8ZaNSL3BSGB4ZLR6x3Fz9gh5O+zNSkrwIA6dtMD8Y/E5vZE6
1Tvwi67wRoTfiGJTgqLHpu4xIwRqKRuQmMABf8WIXIOVYgX5O3pHi0s6thUc1tOkj2VrRfU+yAd0
JRf7NPbMMD6h2m5DXap5n3l91xAd1mPJm8zet92PURLv9K+R4p/ByCFUI5/PjRSvdHViwIr33+37
TYTRry5OTN3Us8PUneiLt0OCxiFUz7NxSbu1dcktUh+yqmTE+t9fbTg5zzK4ovnOUlF3vyyPhD3x
DTBV7AvZYZa8Wr1wbmRoSWzeMPFkkKGFnzHkx2r1GZOXZRmPmgoncoqT9zLxN/3jIm391DFwRc2t
g0yhDsIF1yy0N4/VNhEd0rR03eMskCHshNTq4Ls1dIVXOx9XEWSJAtK8JUi5EUdxG1PWMQ0kYxmL
TK/BN/2DehyEl7Ucd1B3YHh3aR9EV7Fda73kM/aze2NEQvsN1AyPsa0GPp8BuDT30TA+KO5cvHk6
kWZkwWSAa/xWOmJ1upJTx6L+iNRjdSc4zQaByOLRcNTP2fjfk6qKHIbjCNc8Rcl7n7s7XkQ2dqWi
jA/c1BP3vidH2fKNF6NYkTP+fWleAdSwlXMONjPpvcKlsE6DAehWRGO9THuaRcmEQMJGBCRAUsSH
m0AhmaX6vQ0lVnXCfPYuX3MXcKATXSYNuNr5angRQEbC/rELNIA0dIubkiZIYJwFSCvTorkKbXfD
NIamI3u8Duv6bPgPUuaywTjj1nj86p+M0h1P60fF2aOxGHE6nFYMoAvzYXhvdjgwlRfKhm8p80Pb
AvaMkB56ABVMFjRmNKPyoDgSmKTd8z8PZI5T/u47cQuMLCcvGDFzvMYy+TvqMSdrhxzjvaUm8oK6
yvIcWAUjWu6z3zpRwBRc6KAoWRQYKPETh2SwfgLbPW/TtJm1BO9Yc/76C4h7yk7x8aU61iA8srsS
hpUX93DgANxkSB8eFaMWsxC8/TM2QgI4jR2We1X2fx2uoZk08s6c0vQDtD2JvjQncSd5OOqYQZyU
cJsco0VQ1v3NLBMcDccPuM/J/Y0z371UrPvZatUusK4cYEHgx8bubxQ40OJnl7eMBn9GX1yozm7t
Yw9SAVAeip6rsLH+6Cv4YOWCM0fqqEFN0ViT2nSQ8O+fbwuov5u4KNAuNKv85BkryIuabApURfdA
y0JS7s04auYSpL1nwfzWKIWmoCsQTpiIn4ljSuodeCvx5vTRiB9H7Ltt7xLAi4kHCmanXDix+NyA
/43F6bAv0JCUFTZJIvRfroBbaFPjIPCXOUfPMuSYK1s4/+Gh/HepF5XsA5hqiZNSU0HWt3+ljn7p
bd9Rn+sPVY0qk4ex0I5/twyH7SLlwmy7DH077bwMpVKgTEJNXamLsfNScMhYDKmNfK2qUqxpbr/S
vgwb87AcKda+DDdZCgtUv7WtO+kPYw9hfSHJFwpsdYSxxAkzDn9hY8nqMKx9/V00acqr29uyvVKX
BRiVKhDTsktI4USylV3fNUopXFbqpW5jOoJfLOr8RQFBvnNRgLrrDM3/E212sB1KPgJix9V19md7
0LUTTyoXa/nRxK4ngKfFlO+Wmbeu2/4nSLrbba2H5Q2oOkT40MbJZOWMmhvS0u4eDOvHl+vVhkbQ
KL0x8rQS5tSpZND4+A6pLCnVf1RQ3Cv/Lk5EG/Co8UAN3bHXyJRgiLO5QZxIgrhr/owiRftw1TOm
cEk76EsBSUATA1IkrkVSZ120Oq68h2HR8X7xranzgsJYSJ+4WHCkOYrvubNDwHfslZ+5w+piKiXt
X4IxQaZcWaReBZ5x9CJ2SzlEohgGJ4qiDwWn6IX+UI/1iGzxhXo8uPEA0+Vd9qlaII3GMr8IOHsi
ve5I0aMbMuXCErb0Hy7G4J2NPLPLVLRhDhzNz7MzIeWXGEWGY84icx3G74IiyiqAWO1TnY8Iz5pe
sklvQfozfnDvDiROPIn6ZaZ7/P5/ZnUy1skJqvHe6i3BOUo1JGXuMjJWcMN0vskEx+o/9aetsy1O
efRrkPIkdLapRWUPeEZ3aN5zgtg1UJW2AwnQUohjPpi3ym8D8g+Llin8yeZhWn60Q65txljAOEyK
AZ3LB6pIiUiKeEQ6m2dUHYg6R4scCZLgTbvj1mAR/GCiaClq+35FA62pqdrfUaHlKkUT7+oxjJXr
nNAkagLXd6N9B97mcaTkSi9xnMFiwi3M8VcEG/Eox3HI0VYQMgNRqClbOZyAkE1b1/LRi55XmdZN
moEEbGobuxkqzT7PmEtMp4SXPr97lzMnM+8xuEYQDmOtdejrWW+HofbSEjzFa1iZYmPQ7SIwj9FS
210HaQCfyRnBx0nl+3uUypukn/8tZnnCrjJgiuL0g9jDkWLhGzqZYWqXVPMB81qJuCZlA4vmy6Qp
hPDDYcSbNOkMqe49CXBcgwKMxIXvgxu1cvO+GljhCbEd4GrmRA+UZ5P+QcISc6npPQ83dmlF/sGZ
F36K45COQPQE9hLyDpeErgq60b03raNI39Ts3nKqEWaJPioDohpSoSW1a29JxnQ9y5Y3OETQKwUt
DHgF6P/QSRUDCDYLurKXHzj+hERoKIBgzBS01U9Y95Xqd5aJegdDfRvOIv+0YPu2k2UfrV0zqnJh
aIDQJVVd51f3NKWarLkSJcOKpjrCZFrJDIAkLufGLQjT1R+ip1OrVN4FTx0Xg2wOzbJHJf+4kv1l
l7sZElhYfhNg35Z3fE13fJkKng3k8CQ4P7Xz97a1UbO8USZpqA3S4ibcgMNxMEW5tfBfUoxdORgU
issIg3cFd4dG0CDwfYRl6vDOuK3wVLTy77VX7C7GS4WoQ8Qov/tizNoN7XPqcekHEzbTlWaVn5DY
wh5VpZ1OQqYCY1WFg1z/LEdt2AoX0lqEE+aIl/T5/aSkWCKZvvyHMERO9uapMdWCMC7cML17N7mK
FnNj3RUojxC7N17b1SThsIaQ8gpp7a32PWbKUcuwj5QtRqzYgK3BNwVHSLpDGGNyyhjwJatz6mDn
YvVt86u8fool1Mp0mXGd9Ss6KPCGVDulehomihox793Jq9B7c+y+iXnMA5fHy8RGP/h0yGpIMeJN
/SbQPdP3qVyOZwuh6V+YIMJj+tgoQW9joPzZz34YOSu1C2m2DIdbpbT70Vb4BpI60EagVAPSo+UL
Sxq6Wpe2OpS/8eTd4HDJUTpa5G5V3m25NCV3y9xRgj5YG46WmZ9B2eVsQajm7jvTyLzZDdYwkeMT
yXR4YxJjOHLZc/7GTQjiPTEyh/VzHyv4kuBbIaMqJUUAUUcTM0LnMJ4eYl9J7mjfJIw3fZnPsrZT
jHcZvEcQQqJPMxlqyeY3gh5toa115PTkV0mxTWUBNLrEtp3rvPYRWMlKPfySuwFDHxnC48kzhsw8
pGRJsbLsG54zh1iHATdaHa8JAtU/Tas4IpHPgq1DOwCNbiNxcVFBrfsG6FOQmZts6ahuklmiZGqJ
2nSuOQSKyMVTWHSijwzw0C9+lvsEmfhaOhpOhFUxbBZsDPRReyZeVnR4GAbJ4Y4etD1F5fKwXSe8
k28RTMiLOb/WB4VnbPMGAeq8S6CQLDVqgO2SVCbhQz5Ui37ijTVgtQKk1WP1chIs5ynrZlX7n5JU
cC7vg05nbIzMII8/YoqDd7qCx3AfoUbwniTB44vUljsfrjeQ29gymAYV7HaCKfHcnXiP+y3oXo+9
8NXU3j/B4WpfOj9lFiUcfqMdFQUTSwZWCH5/tJYHDx4pX0r5xqUW4Lnwi/YhVcOs7rrmy/khjXa7
ZV+K24NHObJ2tXV1iE5WES28DpU/Hx/bgC6GkNaPF8dB86HM6AFkYsr+UlGPfacy/dzHV0vQP6Z/
c9UXtl52Ti+XsV0mm97XcdPbs/nzzk78fIgD4D++G5MfgMpNXSZYuF5IzUy4sgNwFnvsmc+xoZKO
Kik3b2OTU0Gr9npfVI2J09zLjd9HgMue7T8uD8DMRqMP6TDIuoPBVUw4WS9e7kfqGHqh/DtcPLxI
ua2v0LWF5zUw7wiCx602928dLYGkOSE4aRVqueRlFFM1PrqfFhM55xgPrEgDayMmudbqpi+5UcjC
qzHS06UTzeMBEhhz7CMf6vNAxKATqP9F8YKE3b3COnOkJmlQnDIUOGfcefNcHo5cltW+LMe0CcfP
gEcLgUfWmMcDeUsAMRaNzlcDpvfTco+cFjB9qKGfOZSbsRtwfhV4Imt1At+VfSss2s3F5eF/DvUP
EfTgJiIvmYCnnP4CmEIerhAqe708/w0o8/9uWTNtZ1Dk6qSqHhkOP4zktP9p3oBmIe8OiNOe3oz9
bPOwIlDlYg00uITndr2l7oRuiZ+8WDaLsnpFh4ZOS9QhhJJ2oDfvYUj+Cke1n9jfBc90uq4lpAXW
hK3ZmPGq63qejnreAUze8pRJHa/UnpLBPdxDX7d2LYjldpC4Ckz+8eFbzqLX2FgIzBOkNDse4Udm
jAJ2JmaVm9/uy2a/dZp2wc+TkUtXeBnYte4ub1sNKxyzrS1A8k/sCI8yGw8rsRcAITDx7/MjlQHe
fjICVWcDHSr6ynM8K8gtsXJ9csBIMXWm43ghJsR757XW+VTEAHyf/dH0PgMrmMYcdcnv+uP3Posm
//hcQLfaC9qoU3w4rFLY882y+hNUP3bYM7JvOUEGbpMrBw4wovNZqmaax7Af0LY7vaGkqTSJx12o
547KWxUqIT/hg1zs4kcKvakn2Q6l80lnpjUOPGszbYle91s1ZZebnjBPeWdCNbJ3m0XSXBC/lNdE
g8FuCfjkEsjaojAF7yF5126S78vK2MtqlCTwQH0nPWtU2vtfIG25I48/6bvyTgyPdTis6xLZ9s0H
/JB415/9QcPYlUOEQFqcmrLaXX/t0xrAsfmYdPkppAYl4749xNtMunO1oQ0jbFUnV3EtB/D6FxNd
szxDdcfACiqYZFgXrtVGa7WFWcsG8253oE71VdUssLov9MMZ4rtxrx6vYUZMfhFXd3SzK0I+lYaO
NVs7aYz/d6cIsScwUYRgMgUZBv2RY/jTYgG54P66pzSGJRUXzQ8hSqnLMSR957fQh6/JbVjBEkdm
L18YQGibdafOxVpxm6BK6AMJRCkWEjvmOQl2mi0P59s6kcIHKyhLakWsMSCuR+6YcJ2k81sIlI8H
ZN7Z+lBYO8ehU2qEvs4hed1/HJ492xEFSDOz3R4YRxmXr2Eu3MLaeXICORNPGLkHMNh1TcVzGHck
kGx7ScSvs5SU4CxuldrNqXQbeMpo/GXOgOZE3IoDCLUa3B2sAfm3wqwmPIwOAcoO2Lf0EpShg4Zm
PApFMiTka64arvPxbmBuPnUO4Qe3s5DedbjH2vWvc7xlnSAQCbUJxvERM9bhCQ+5V/LnbZiFx8jn
yZtY8uXHVqN2yfurK1OGioPT0aQeTQ4aq82fxakbqFV66/sEM8jfJLrL3ImOzzulw/bGscJ/aR7Z
aPsI7Dy211xnk5lBH0MTFjOvPOSA7x0NobmvQzGOHK+3z29D+PYUHsC1nkgWBXYYRDAPqnPViP57
GlTBocX2kqsaNuNLT4b5K5F6+xtLYqy+0xzUUwTQkeeG8gAsGKSfybMRrGMBq4P+/+JPn4ythUjy
7gTX2yWITC+hn8LunIXLFuzO+fjcKqUIzFGouzjqUW8GiLzCF63qJ1d/l+B8zppRx1/gWeZ640RB
QPuem0wUbymtPil7yLXWo5dA6s77QJTU1PVGZRA+A9NRqYhYrEUIzX3V6jq5Ieb4CEg3We1Ddfnr
1DpuW5PdlYBTzQgPwnGPvdMs63KFkATvCsXoetIbk6vW9IxDADXGZ6CkQ8yjDaDg0xCRH+hjIW/D
cVkrzkuqlJIM2340scKRe1I2VtAuRcbTCAc5vp1ZvIcfN5R5R891C9WoxRnnUhOOhVdmyLSVXtRk
WCAgwNwPTMWODW/frK3/cSQmS3uo5hGdS5XdmLc/CbhNBnr9j5vafwcETPt1rQvVa2Vu00E7+EPE
8L3hemN341cUPStS85LdklF1HYURVJfg5QHlCaAcEU+17+6Q6SsCojuA7aM77ymHffj6ItEXyy/v
L96lItXWR4cBlsZjhsn2KUGwpV15kO88LyveN4uf6FN2Fk3R8qMUUjwuLhibsY7BpeY50p0KgEP2
1PP3lqXHkW6e3Suefmps6tnrKhdn7NidXykJwH/Qyj6dz9ncfxdQQ9FoE4Sdi2xzQvMy2u1Y7iSn
v7gXmsUR95LOK/cNizhzRYcRULEic269pBiI5UF+mhMCa8MbDgtUGr68Zko0oJ88QzcdjENxqMzf
xVUv6JkI8evcoWCZlp+MlLGV+T6BCoWfLbIMPLnXpxJRX6FEQvryseVwhppSFP+dyZcNw80K1KQL
QlPs7HUCo9Gj/8ScbJ0ufxIOVejawKP2qMTZmLavU9yA6mnVvLMOYX1TGq/szk/LY0KpnY5gJsjx
T0fjN58Snw+jLsSDH/FTWFtYmzxO1nvkJ571XYD/z5frlURCz2x17N1PRbm63aSuGYTQBLWIRn1m
LCsooQnix9n3okXQXbSj4CcfEjzAsBPzgV5dptOGTAmg92oOr6IUXZ1EwvTpD+gAuklKv2EGAAKd
eAO9bdgsbjQFHop+hqWx9lYd694s+qipIC9QvH0HQYg/UqwrHJrTkTkiLmPr3rdnKCuyGxjXeViO
TtztZAsZ0eOUXISquDiUDPOY/iw6OAfNqo8g9CLTVOTFhlrdSc9mUzG/LS2I+3p3EFYv9WwMCzcE
czTFhfYpHESAuXI/fsgbG8k1Rvt3435ulCVt9QEuYy6scp7Z/lrCb73UEbkhCvPONhvJsE1uydHN
6YPTVZchB8xNN/VxpCNW+Ai7V3FOTXniumArmlXcKLnpUJsvz81nZItgtlZdFHn6h4Ldo5TZoPXI
Cju44tcyzbyVCX34gVVxmq4h2d9rJix0Y3CVy4/lIuPepoxhuhGvB/ckEAYoHzFBZN7aQC60K7/+
iQgEHfVGZ6NGnPqoFgiqAsUvba3zuRSONgQUkOQX5yPeVggqPEjpziPyxxx3w73y19C6bX0Cl4QM
1RFaUGpSZlOUcQHq4FsWpOkJy5o75t4i6S50iWiwKBbJHTmupvCg252qPUEmLtZ6oMlDtor/FoGr
ZS9m1U3qUGiQgz2mYZeaPqPZkLJTwmCV4vVJSIGyM1plkto3cTIWus276NxoUaIVIV0l0TbHvC0a
UastAric02pOs5jjvHP5cKHIgT2WoeqFCbOYWgIVZqsTHHdO1H/a76QdKW9y0zuuM4LKJuvAirou
mmjAGNeHgDG9x/4NzdSyLrAMxihaNkOdkCGjFZnLKEsDZ/TjA/q7a7HUqNyn5xNb2NzS6SNCJcIH
GE4EMnj2uWbZtHsordAuEGsBiiPMZVUOUF6/UnfYSmwGDGr91MvxlDSzjzf831He/uhx2iGmphgb
6GA7wlSznwvpk12O/d5ENh3hY7T+IX/eoL0LBYL863ZsQjDcid6UKUGLbiv/TbZaT2SMr2v7Q5jF
d7/9t9D5HIA+Fy5TrQ/0NrvQ1RKfR/E3quEoxEk+1DLf94g1HGsIB3hzNL7M5caz1m7p4uFpXyU4
UZ05qlUd4EhOm14BeSVFiFFqs0bFWxF9wqNrtLu5AgzxmlFCT4Np1fvrD9gJa4lzRx26vT0tQrq0
AxsIWLwDaaS0sZaH+PdWcnaU9erffQBDQ29ACiD33cUlCLnjKKMQc3AZl+GW09x0rTv6C/lU/2WN
EgXsDF0P5hiHhqSy4koQOZLcIp4zvaLvblcIt7FyfSO7znibdzfrOdPGaZBWyerQw1Mzjft9Qfd4
qj0DfBfQn4thVwEYRkdkD7vmAiugJwr4XoJMszMl4OZNQ2cpbTiYRMTddxhc7SDQ32iO7IStt4ns
TC1kFHn2F6l6oLJwTuEovguFdpkuNbyqe0YaOGwWaOR5OLJuyZTFcpNAZesRda1f0EGylDGyKWHN
rHcv+OH9b0GJ6I8OCoHTib2AprKVh81s1fKDDnMYfkxNo+/Dye4zTXyy968qN/MaqKS5qPKOaXu6
WNXHthiluY6Lgq++lGOah2sg4giTHD+X5PSVXQKTKwkwcCdO0mbBBCZeMQeBTHV1VA4CST54c/1X
fIkicoN55eO2NCu7a6pMNdO254ctKrPj8bBKimXzUK8pdXyw1F1klst39ZNwEKpMyzV8skMh1A6j
YJSneU7ZHFU1lHD9WTLr2iqShbLsKoAmRw1DxbcY/DtfmclEnBcLOSt+eu7VyrbL+KfW+07rAO3N
hN1g10k+DwRk3hTkygL89En3d3P+rdWGpRIM98pNLcpXazV1ffNO/1PGvje3UUhGI1NPZ4pHB8+R
yaXW+wBbrd0oE3Hoj15rxDvnbxmkWI5DKujZuwlTAiU0yDZSkfdZsPQ0IRCOoEQCFcrmP5Atp5nE
RjLXXM9SYEwXVz2Vgr/LA6RVOZ+LkIHpwVpzAwKSGWwT+NhnYgVfCOGRFewxolVzg7r8ZWlIBwGp
rE577PsNhObLbigBA7nBirIuIFaNj77wv3qaenGu1PO9ju4YqfSTa6XcqrITtGex/oCLY3OAt0Ea
8Vr84UVBsUF+fAWYzAkulBvnrgyFlivjnC1SD9AOf4yHoiu9N2Dmi0cQUkt6pLevEq+GRwC8UwIG
2DZaR+V9gxDze4wq73nwujFiSomesrdOoIfm8vRQz7fgbKIUHf+vWzekVBGn+yHgy5hpo/zPTpbF
iOS5MSKGYX18D+uqSBiBzy6WeO0wnvWMKYyvWZT62jabrh53+aldh1h9c1kukBCBmA/J6MhLdRPX
WlS571N1fcgQNyKH5X+zxEXnzLmeZlAsKN2JXz30M+bB/KuYsZYaw8JwS1L4d4OwunXG+VcZmTtH
EYzeJVDLX+bElBFsT+mQIxqKZuc1LfcrXvw8qQ/xI0AdMMNGG5cSBNsA0LzBCDq4yZW1+ilb/YjO
qu5OEafGYNiq33Ovm+h1jBEIsVjkYMb84st9RPrYXaIOl0EBgaLPwX9lDTmEniW2kSZ6Lv5YJB6+
NeODaU0lOfGRQxAWQQzPqr7z2Gy9cM2Eoqtby2d4l3uZDu4GFbHd/F3oed0IMmWMoXVlisAc7cJ3
1kdMutlfv6/Y+9hXLiHurxO5t/WDp2vVI2tIoF9X3WKDQAb2uTfsYQ+JFVXEFoqDTmGZNVyiNy8P
7xfmD+FPNXEuimaiqGVVT57P3bj4L3TPIsqbqNtkjc1G9QhKVaj6+uUjLXT4qwCKJoSlDDtML0QC
vIToHZ4xdX3T3nhmXuX/izAU6+pQ3wewJ+tqHZbflxvPbd47oPjDQFMT7wwif5Bg+DF+XKRVl4Jl
EKVYJfaAyT3B9kqN5hAcLg0/xZ5kUFDu3lEJ3P0B6TGKZwagvFIAo+mhh0AFrEgBArkVV7bRBQ8y
/8hzAYktkdM7Kn3L0M+YRQhYpwn0rv1jjnZTADr/RWYImmFmbQmMRgy+7cIrIlUnPmFeH5o0CykS
5CU6TuKlGjRAQp4L1dvZwySVn5pFy0coKmaOSVqYOrQluVwCITH9x2kb/Lg7jN82UOom5NRfVzcd
oIgXIEcw5tblsrfE2ANYVX6TRDeqWMC1m+t+PjSyCbj/KfvzXzxv3JLo1OhlqhCMO2Drwskk+atk
of/Vu8f4vsS3vaGxnWdcvzo0JiD+IQkGVI27uuTfTB8j43kpbt0ODVzOxT7AVJsOED+6nrTSAqXq
5GYzWEhKlUamYjoISK3ImAnyxPv+19PlldiMOyjyG8JJGQReQIHfLqZFQ2huP2JU1UFBpqgMNiVZ
/w/vZdFuXIsBhlkGdSyPoBqZRGCrfHRzqIA+w8FNOtmD3JPYWFma3lIE6Hsh6dKSq0F1atII+Nni
/M4CNhNw44zB+wukSTwgD5ABGIUNAlti82H1PdrxM7G5o7wrWPy7Q9+Mwqk7u9s9RC4s45fF14nR
XjYd9XAk/QECeCtd2D/MGSb829o/5237zpV9bDXdi9Y5zBuYjQWcvVOgtNLNOY0MO1MsHJbia09v
kmdELmxqTxAFbUsOjvGca9GhxseqAGOqSV+oroGhN0XatIv/B/IH/aEFEKXuvmgQohGTYibeAb/J
1Njj4Zqm8xsl3WNThYqABxSntaALE0pPIlHJxPvItNuk7B0sirH5X5eY0bR4DsjEi6aDk59wEol9
TYUFbxe8olU9JtpSZXSIzRcmz/MNfiL0lX9lPq4P6sNGVPzNvuV4GJrb/uTOrm06U7mi8nNC1fDk
iIO+fj8Bt00EvD0P78sEdPX8nF2vhmQALNCB0jpwNbQug17Lb9Mzc8epA3xyjoJbpd+O97oKD0a0
99vo6/v1BHWFD9ahx2qr0LF15I2feXgFfmCWTOO6PCQKGzDBP7E8wILPPAkosSj70xkIBdn9IiMt
s06txCLJO01N795M1u9FEWiYXbNaH2bmfxmxvGOryqto1K/hdJRDzcQBIcCSVj13Dvt19pOQAkNc
ZIvh2he4thD+Ul6FjTvUUzTbV2pe9E4op6Urd9N2l2Jb5K7Mi28IqJIAvTKmSOD/4CdVDoh1bZ6d
xXYyBYfjoWfZbqc3R3PsrOMauE4ZAkKvrJ1CGkEEFiBmp6DT/KLmrQcAjmBrkDjzlt/m4KBIoJZ6
i9sV/U5p+Rm7MLszL9x0kfS33d9SinqrrnPgNYRkIXAgTjRznvUTkh5UBqcO5YfiNI6XyLJ3q+jk
QgX+boXYji7ev+zxbm0Bg4pjEu3oC1VRwMKDKWNmcXgNytcg5bM7Ct/Y96EExkFrqLC43jPQcYWV
qc/S2qopq2hBV/KzHAA5rr9dB8bWViTsCkAam+9eIRiepQ48Rzo7XA1dauJwIi3and2+j2g4Odav
LN2tqhmQAoT8N8H5Dc5qNIfnOMn1W+/skHOzuvvzT32gnRGsC08sXPFk1QFTUEiPBrKFlgOqqBaj
bJMt5LSEC/nlQbCshnUOU4+fMxWRfBQgoe7wMYBwRdR/VAYSA8/8VjPMGwBPH7We6Wl6nWzW+7Eq
S4LaMJFwV+6qO5oNgAfcIf8IHDwYSzfXz3HUx7jxTKwT6jurrZVCB34xNwf+4q3P582UpPE7t54/
Twl+C9ZPY44jLjlFDHrfNI/einfOO6z3m/fSjgJx45OsBbCyhZcwRkL2s097XRLVMNiiEA5DM9zL
07Rh3xa0i00sWWZfrqbOvP7Dkd2zMR/iPo7ICgRAy5LHecNTpsGObtIUt4ZONcqIIDT701I0TwRN
T9Nc+VX1bvBSkUbuuFH0PCirnwq+q6rNP5YnY9IcIttlUHA/TFPz4C/0w8UxqC/BotLUf6ctXFAd
odCvP+ELZ24N/YvedO7L+SjQ4ulsbqkestUfDIHtOVOhmH7/6swATVDcHgBR5wk+xAKG1UTDMGFI
Ap1jI97OuUMla//BzhqdL8sYW+TSQ7Dsi3OK0TnULxaOF1UyE8UO0YG/Vip+sJg7phpCVAe9/LOD
ud9njeT3UUyFupQFUbRt7Bl2IZtpKi8NWyKw1Vac6QWU10jdYh3+s3VNGklXlJ7lx44fKLKI+tdX
+eZ4JrJh76GZC8hbyD/jGFckiHff1aF7Vx0yWrxW930MB4XFFgmSxEZ6ko6Nf44xqmhQLaTCnhMw
RMpo0y4gZw38Q1qnprH2NRoeLTipw6bin66AAFzYPWa0V4ZBbZ51GhvSJm8ud3P+4+hBoAXtJ2n8
/bD2DB+bkYThm7SviSRkBKExQS3Phj0CA9YGFtuNoi/xVdlRiBuWhx2NhYkG1C4kbt7nRvPWZZze
W6Sl93UcRI0JEUr6qx50zxt50BkX/f80Bq5b9RZfJ5NxBSCBRP8mGuz8MVU8aXO6oXBB7BXyQfaL
JirdmNREpd/5SuKws5ee4K3iatmNdrUf/aff4Ubiy5dLCHtyG59H+Sq8U6VTheQasVcqYw2umHg8
9mkrN49r1sG8wWELxALN3LlQe13kxk+ACccmO1jMzxbJ/LqZNOb2wznTAZhw0qfQT3BWO4rnZCQw
znl7JpBnB4xChoQP+b8jdYcfzu3DxLs6R3j47GZhiUl5QhjVe7n25SYgU4wP30dQ+36+IWvDMQ5j
s24/0/2DQHlZcHIiS1svPAd+keAnI2GJXkjsCtaTFqyssSN0WnQGxVjwgLXLaAAXMkDKmlL6QI0D
t5lya9qWanByqmBrKPFHAG1VCeY0X8tUo2xvfod/5D+9ovIsqu5Lpu41nPsOEpjrB/4yUDfYOM7E
Kg7hLhay8no9yQMMgiOdzQztjARLqIGgGRnNWkVyA/HZ7F3RNg3YS3R4gt5iFkru+Jpcx0fNSrx5
QTKbAorNnvF0iKbb6u+nWk3kVAivGodJJ9EWdMtSV/Fwpnt/b8d0EAgDkOlV4J5pnvm6iHfkecw8
e+fJLNTXdhnYglfGNxl5QEQi99CAUgyvL4AVfjPEzdMcKOJQT7Sb+QqIGJTDlhM0Oloid1swCBCL
KmwAzHoqwYdmgMhyiVEdm9lDK1ugFK/6ztziLmfOXgYu4zUXZiNOOemfsl4q14ExdS2LLyBaDACM
estlsFlUDgeqPJDmrHTP3rDifS/gMe5ROIfNshbxH1Qrw+mdaqclyYYKN4XKojEGAzz/Yi3RzE1c
PgAhNhJveApNl2WzLMpkiO4iomOOQbeSnNZo6ScVtOE1DSpBfOeo5tZweQc7Z1xSNthB+lOxQWNV
U5xcHS9JcR3hsdlJR9uLcPwgFX6PgFFqGFQ4uoG9OV9XSxT+z3zqxao0lcEL9VeuuhhH+bOF3bkZ
Zyla1TzMWG7LeMK7eTSOUnB4YXI3WwvLlcvNNlE6UCb/CnCJD+2rSOgMTB2GKvbvib48bg+jzqb2
UYeuPy5TUlM92nUqo7xgfsefvWaPgu81qVuI0OpmuHtOxwwyMqMOi8oRMEQXzuJTr6Z3jBrd5Gia
c+ly10/zY21+nqbODp8/uOTbrKGdQZh0eIoC09f7/bA9UVtoJqdx2pUZec1NcUuyb25EN60jPmzf
SRgtVn+TTl0JXAcgYL/j/VPLpvffajkKlTppmjJakz+pYSwulI5TNDwLCwMBx7qAD+Gsh4EkFhdE
oIFYDCywtoJWIjCbmuerLuA0m3+zIMMiTdLv8/jKzpzfYZs3bNo/GIjpeCNTYSF84cdeVnFhBrQF
ogaJaXKSbdryzCu/V4NmJKYAGqN1gafMnx22Od8gDrMlbjnH19ncyiavRub44iNkc5GSZ//WUrNn
Kz8G95OgRy1MzcexjYIK1FB5hyjhU6oQfOEphGrJDDbfe2luvo+JGMjeK6w/2PAhhG0E21aPrkUi
/aF9/eCxA1ecn3O41+lozY2sro3pjKKeP+T1JEbL4dyz6S4k/3UmRoBtUJ7LVkq6JcQXoGkCd09i
bA5UyFNkpViDd8KCnmyj3ijJpuq7BUhQOJOLwGBNlAmMTYuPYWxKA/njWNvml7oOucii54NXSQAn
XLrxf1b+4xTvFqorhBqex/LH7edykuu9xvmpSq9X7DnRUwbbKGhxWLszvEWoAIGB0S6o/QmJRhjD
BBeAZEHrkIKDJDZoHq1xnQxSUmcMWQqNZpmxEG1KTXcrt8ww+DFhl7FcOEnkn3GpP2JwWyypQOqc
k9PCsF7h+LBW9gmlpKCu/zURkS1E6NZFuoQM0vk5yZQucYXNEoCPx69xNswn2UeWZcCedM6ehwmb
KyHXSb42Zdtft27O+4OsJzD2caxBXcjPV/joHvot4o8TYETS40VilJb/jqDK7zwO9ogkgeKWhB1x
8FedInuEprySZbf/7VD1VzKBkaEdkaaIBIXfLKscVCETCI41x99LhR7LlJt6m5kXh+0qmW6PweB8
/21JM5e9YAKl2lTc7cfBcWpsGNfugLHn2J7QY+YDBdVKq0WocRtMkcnUbcNtDWUFgCi4Kq3B7zZ9
zD86xgyTEgnK+IS8UQaU8d+fLMmpxSXwvbW3dYFzQX8Mpp9VUORSkKt4TGnD8vVQeb0ZWDK5LSrC
lQSXeyMZ2W+4WV/pPpSdcyDZ5GcsHTR3fk71GlN25tRmWHDB45xR8SOeCHOlnXEYHuOV+ki0MH5U
Y9AfmAALJcY+IwKE9Isa66k5AebOTfNb3SOva1SDUtsXGmsV/D/SLe+C7Ehrg4VW8AKQPjVIPhBZ
nrO7Gssjl/paWLjUBmx/qq8czZeyOO/9p4UaFBNgDtKZw3ZhF8baSg/lHfu8TjDn67PXGAaPa3I8
obilc8n4lMe5n6xp/Zbq14p2dndNQePB0J3BpAduK5ZStsev4oYgHByoD5/GHb+/LxY4gKlC04La
0Fkdd5UcistYecagVzA+A+PgA2PLNJmFfFxHW2g75Bcxb1Gf7CXAVzfYe+O+/9BDAwCn7mSt0nyD
fAFp674ZBG/oJEeg3+Z0HQv2ukZg9RFOenszhJUtT1oI6PYy6OXyxlRK5U0U1FCUNJtOJ3OVgnwP
jHATFplikjpjbnVV9PWThDb1Jj3UI9OfzTUbVjOp+8HuUk4HHYDqiJxGfv8Lwm2jmqukNWA6iAQS
kstNJfxfzcaJV3Cp4RtWUSpWWw/EVOcVvIT5ocTsxGnr+ImEEmxxq7terfP4LvLSksrg0cIw//Xm
JsesQ4Tyold3PnUdh/GszBMfRlS5RmFgQZJE+tUcMlrf5T9xhWFP9lH7ww1JCIhM6NdzV/wS9mHG
qB1Eh6fWeFUKnSC7HhtBVtst1Q9nZGeHwOK5P2xJ15OR3/D9eJzgqIEjvU8dNr76jWGMGVeAUiJA
pzvquzIXZLB3hfnEJWRSQarEWzvaEjKI8w7SFzHJvvOqhCM91pxqK7r4uYarW2A8EIEGjkh2m7s1
jHJCNoIEYqNlcJRlth+56lN4S6RbEaoS50rYE/0Bf7NZm5+gbcrarV5RWRD81XTrMoGIycCeuOX0
P5rVRkJhxVhAj9Hr0A1ywqIKIandycv7ckIJtcRCph5zoRSjVl/VtLosdSHfp4araQnUvVuUlVCD
ABWzBDYeeU5XdH7wsNVNAx2sV0UDNk+Ypw0Fx6yiV5d73L4AfGGiQkawV8DN86NA21DEeB/Vykto
jgEbkZaFrDkDDN3QgtUrU6q6ma3YzwuS3WFtzMPy7EZ3ldLYkdXskOUoz7FYcVcJ6PdoliomGRdV
2O+aWtcIHzoIkMdhIIeCknW7NniGccFpfA3H6ha8a6e/En5aTj5kZgYwmj7VHStcAm8V+F+dyPDN
CJZg2KhSpt11849cuEFSnvTpvqLMgbNF6d3MkK26yy/DTrZeTGWWq5/mEFCq7qxZHbIefOeYDXqM
HcXaVkI+bcp+OcGt1UVO2cGKn5kWgieCMCu6xpjWOm7XbuwV33zu1u+O9UxvwMBZDV8gez+OpZtW
bagfs2XmSsAdB92B+5qoAas/ykovKDILV6EowG8EQNc/fy/7pjn6WoGJ4PNtCgUMj4RloHYsLvin
uYPUBQrJM8lp9Yf4yg46vvjehGg3xJisqkrZJBaPmn7YpK3ADC56SI9lbLOnC4zXDbqvcRCjtgRV
hn4sWAu/XvtDj0fTAapGyNbn3fMoYWEqZ4NaPP9l/4bnk+KntWj+iweJGHVHWUvKfyO3Olauy89X
m2ETSfepgvkgPb588H3gQ+C8N1KYlwctMORhxqaJ80B2yaFaLBXrHaw46y4PLW/GzQEJUK01P2hV
3ED7Mo8kOzNCjBcVb1BiTMTbhsRJ9LJZEoKxZ1tGt04DhGA/m9iuifsqTKWbIanSJJGn5qFeLnUJ
+ArMrUvhK9ekZc+WcQP8yhIsRi/lqxpba8oBd/DBvUeqDDv0n29OB1QOu+GWXqTpapNXc+GKRfCf
9B49sYAiR3wt2aZmnz8/sxLXXfLAmvn9v81iYjxNoh60wfz1TOFzZXnDq7nr3OIgjoxglzwo/OXB
kaitYsjap/dnMh9Aq8EYBnvjMzJZleyRps9jqLsI0eJptBD04AIBMC+/5XxPZXAJRbwVsqZA8zuE
/yh2r2p7bCC0F8ShBcfnlUgGo9wMBlxosSZJi/3D/sfN6WHTZfFYFnZDp2hKwRuE0XfX6mrf4G/r
370Y/CUa5My8gtgjEJ5TbZ5t6Go8p9+h+VVCtUwC8WWjwqjumuU55//6ppwhoQ09AdP/3IweZpVK
0f2nBFJnjMsugKT4n2q27f/sAP+o2greoLG36fqGxcmnHzBzeb4/n0DOFMEwv2U03IK46BsgjC7X
cfJkmqmTkp0DzNq9AKTgkf2+qiWfZ0uqRHjcnP/iv4nW47+Nn+0KKaZqCRknc8h1R+uI5GDqcSU4
tzcyMbYC8zf1znBbRxMTNNUpWk/yEOOf41CNMmHAMuyQFBrTxjUlBCjc5WeTjDn1fSPMgtXZu0bs
Yp5A150gpDEyghv9jMUIbXmTGxSvGz3E9PYD8JAT95+SOptDAvOPv1DOMW7rjbQrZyhQZ1/d1YP/
A7tWl8sMKC82MLGO67eIhinS2GsowwaQC0xjsNFSdq5UHabLywowS0N2vmKG7VL01ai5x9nTTaC2
6IsJcATginnzrrBaYSYFpkwdFzZE3YSJHKmzAix2ZPXkK9CUrUphm80CGMVZcUd1aK7n54zHuZl+
8rFZbJgODgSlf/TsmaxEs8lrS0mkhORpRbQdc8J9g5MOnwLivxmdgfwWSgGjbTG7P717NmHmiSdX
A9oihVQmMY63nISt+KFgTNvVT+JYV0hc9pP0PtgMpLbvKJOLWMAVJMM+mk7hoiVMhXY6SKxivDqt
lDVqAlLzWEOzgmb0TGfGNM/dE2/TXZTLPLFCo0QL7NBMSsUWizBoSlIo+a3X97jbZnIgzb1kvt6l
y4G+QZhPwlEwtEDARyNP4IBPNPhZ2fjf0pPE5vXnEEpVJAJ5QUcesZ5jmsobcbJyIbNkz/WWW+X6
a+4PCR981AHBz9mXR9uyeH0UsPOLoCUOBArczKU5DXyE/mixqwY/G7SuD1uVAmS7Pl33HYX1GPae
L4480dFblX0fGLz8L8X746Fx82pGFarz47lSeBUfS6bNJ799q+mGiHDDWgAOLzQHB4OHmgEGfT5p
Q7YzKh6lXe2UYL/l9PlLxw3g5zRQkwkamSzIiA15IObMsAyiO1tOVY8SksxKjqCdJ4YuhjPLJ7Ba
BDoHiPmKZOS6Z5YZHVKvn8NCqJJ07ay41fq7y5+DyG6KMnzmW7k6LTijgR8NiuJx+OBXcjU+Ua7V
PeDuKqVkIZb5zdsWW6AudHf2GHjLWjp1BJBXHBnvKZN4bGnVzAs3Qw9ygTyGujP9J+43GoWFA2HM
IGGFkC3MvXBJrHheslsbHOfxTfzkA62KXOt2wWElFZYoYOQDQ+eSgYkUCJUIZBg4c7CsNcIgzdGi
AJZf3Iqj1Lnn6HMYdR9I08VGlhdr+NBldAaOE65eI4sQFqvNnw1n4YuZxKlIE0Tk9jOzmrLG9Ntw
iExWboBg2c1AjnyBoRF0IbH++PMWn/ISo74klFAf8ahgigYApRsDRvJ5yLTsqrPxu9rRajE3A0B8
PKWZA6C7WQi8jg/k4Z1t1mCGbaT9G8y0CoKam/QeXLoaMxWrWJhxATf6/a7V8I7CtEo36+V3PXvR
Df+jwBlgeysV9b5wRvzmeALsSP+uzuzwB8gT0VDd5ujud/NqCusN9i6Z9Czhf9/q/HLYvJMOKWJ1
2nrOMfv86vAd5OP37O+aALtykal8had1zJKKAVsUI7DpPvX3PxDdKzIs/fN9/EYTDuLy7GEx4LoC
BCApY8O4HkeF/nBKs9J7yttxwo/5XSaS7/58NrlI5rXJUfMNrcTuUT6uB4Ivc4dGJMKACP+4nGeZ
MyeDxakkS8+jbxnpfuk04iDhnBqCujkDlo9Y97kebAyB6nMRiMprk8avwD9jNSK/jQQEGEv4yxCu
M7BHRRLse4+DIKi5bkXk65pMBB+cEj30fw6aq8WvOmw2OsC1FCqhjAFZdZJrzwjfCa27cwr1O7JS
W6lNBWJ8BpDY8Uwe2ziVXe23meWqxSJJHBT4Qmm2XvhsOSTvTh0nmsHzlP+A6h8DFWdMdZSaYQp4
8aoqqu7RSOnxjQssA4gnpaiM00Z6XcXZ+Qetd71J5K8SaNNnSQPBYprr54c4Oer2Otz5p24ishkI
QIioQ4QDLWq6qL/NwBXgyi55Ia4+G1guG6WueAApaETIZAViJ70e/Zn56cUypJPtJ5X1R/mgwSkc
nMZrFQHD8CkqKZ8BAkSR0C8Bp+tjY0cVw6zhtlcPCr7MoyWW5ai0OH8RWG9einrDeSgUh0IPYUn6
ZihNyzZCk3z6ppvIQiyfroEZv1bKd8tEaYPn/eOW5frZ+4T9GR7J8vmoG6rocuLgqBVXh2jiNz+e
NwId50Rpl09iLJnjKG1CDy9E8v8/YnTr3EedhgMgJEMmU4RHaFTZ4J0U5BbwLWpY+I5VK1DJsABn
zwyP4jyYm85TajWfyhgwq+DGoGwoCTI+2ZPaChnlSHN+DEoikpWjZIitwZBieEnDOxu7kRlib3tw
I9JsMc+NBO5n4T2Sco+DNXIjO9PAR7V1EluaPDid8BWBkPC9nt0R5pCs2XKugEMVi7J0/SrNkHqQ
bHYU6177bRDfUbTJsA7A05xQC953EvIoxKzZc0rlW6cDarCPSRcUuqTA5Qv0UiDf5BVNQCl3AZvS
hA5N4Obf/2hz+OjTAiH7wYBTg4dVfqutweUcPSh0FyQiksBH1kGtQ6jpHokxKHKWLS8X/TCIYNVl
XHX39gDHn2LgamfBIb8FdHUrigqZxBcxNYZJVmp5XOk3drT4l2jDnjVJ+iX3+tDW/I9n1VMfAc0b
PxbEOEjyneCK6xX0hOet+D2LO2Fc7N7ilAqnHS/+E3PICS26zGDs5NWA/ZSQoqpXU6v6aZRLDayC
jCTw56llZ+xbLRfWb+iOR+5hGNBbw+fyeyNDdiPfbWOx6Xyh8s43Lpegk+5z50r59zoiXgit56V2
HO5i/d6T7cRhu3xu+79ylfDigR5aA1Rgg8jWYxYBvIQJ5x66YIMT+1IAyKxb9x42NLyo9w46lStW
bRYi/kdneRq33vz9+YtmumvHaERir9KOvNWIwJ5aIADY4GXEXShxnKEmtgsVKnDIUWsZ/A4Fxoab
zquEC7Jb8U1Mr4f4rKH002u5CwaXLg6dv1nwNYe3N4E/V+Dk8Qi7eMIzooNFXuvqlnX+yPQYs+rt
efzSPAoj+24qPazQOLM1enUwUCCBPM8EwIxbK8j7KvXcbTX9HpQQ/APqdU9VbIh+1+bIS8zVWtrF
uFVKBBu7dmbi6/Zc7usqznCLqIZdjGXUTAKT1G7ZC8iqCcYEnasiVdEiu+R4OV47iglr0kOsOKWk
bK2ZWagLEs8o3PGhsaHyeV3T+OwzWC13oQ5R3lSOnNRyq1WwW04RpKCUrdSc1c8nkZGt/LYXaieS
87TeXF9C1KQ55YbXjmYe7S7AJmPzk5tctGrDbmDG1TvY++wxm+JfSo4uC0drC9ftG391lmwLaxYo
dF3tDBzCqknlXTpB31gQU5sRClOYS5Ju6mxXohCYjg40BdlMqXpsdUejzJkaIjXawhB1KEGFxaIl
fCa2AX5NSvjZR3foimRE9hu+Enhtycy5lin8i1TPPn4Ayr6lZ1Mfnw4aIEXC/v3yiE3hztmItbCe
7nIdvJ35+r/aj7XvQAJ6j8d4qXeMrz+XoUTo7DeOm8bLgkg/+/ESTBz6M6GnB780aCMM3IU+E4xb
cjmalmCMbBXJ9T00N9OraL8t1HfwbiC60UdVHfyN94KZZau64LccRfyWujBO1lNwubvlqo7oiESH
+p3XfDmDSUmfay8+UVW88Heb/dS28ZBfCapyTxGLGpzbXedYJhko1thyIurRFrprJbC71EACWf2m
I515uvRmhMYcBwiJcJX5xYUsbe2KIcJSyM6efHYOnYIyzvQnNVbKbmFr6bZJJxYxNIOa5wExdRF6
SYfxH83BeNzkvdqWcq7ISvJzELJMO826mvyyK8aeokvSqWI0PC5FwETXwuOThIIQ/zZBRC0ybBde
MPYTDJ56jCveOCPO6ZzNZczupVYeTQ8WWWyOjfTu9mFfM5PJt1iGqzhCEwbViDaK8JLiba72WQz6
QnTD13ilCfYi3dB3lR8U5EFu4eZiP4rtzK6XWC52ZNskmHHE/wfDpBaZdaOWDiYF06Oil2GyZz5j
7bLYgCwo7VAKwpo7s2NaSKuBSAbLXQx0QWSvjWGBHaoWQ/M1xKV8zJ39aecRGbpoRc8P4LhN/8m/
RJq9DDgohrnk+QDdz3H4qnlLaJOnBcbONHKbrDfgut9pjXSBRPVRCxaaL4t12f34vVZAGtebVmSy
NLYlrSvjjXYsmc9KAdgd3ZOH/zGLTsTltjv7a3tzwE4p2mQm+eEufP2y55C0SS+tNX6qzppyghWl
tdNtDa0hGeOvrBXgaQmC/Scye8bRmv4vL+UaKqUw9Kr84ipFutFgR90wuKT6RYEUUHLMvI6OKMf5
UnnxVTlqUuDQ3XTBhtPgWLWrLsG9sZ8/v4fefgUplVEx1KI1INuaxdzjPpuXB0qn5W49B6mFIcjU
BO17ov2JrGNydmzIaalWBXsHd6zv3PctdxnoSL8+6cwGZchTVBosn/J44bMfp12ppWyqO15HFJAu
4jvLdU4ZPZIVpPlWfG44f7un9x0B/KqT4uEQYd1o3FONXIPzx7qHQOWIe9NOVBdorvSqnMiLkv42
qo3rc6UoiVGUHRgtcq5bcYLt5v7tqGOMvwNHhoj2v2qoSlZkOVBU3CVY+vq4rFUL1O72iGTw72hl
Q+HUXEozwx7S1PvljhDfwCJTYGv+hf/THNUVbkpNUxyi021oK3pMRsKDxVOkMKw8e7uHD7HCKAQi
q7S/fAlD/5AY65LyjMVrgHqlbLaszkcFCOxxLGGVHxZBGt6N3yvWYVkOD0P/5ruZc9cLhibhDXGs
jyzm66kh2KlQGP2oJBkY/F1UkF9gI4Lgj/l7uUtgv5mt6YbewCQMxjQkTwJowoqt/wBqMfWAhT6R
iqKvg54t0r0FNbKZzfKSenPuCg2MWRkfVeSlpNR+qGZlZeLZgD1MgumNAYirxYretNwrm47VcXDY
a0KbKKhMI8th9wuUqpfI1RardFGgfUNsUTcmfC/U181qIW+B0lCRDXvZXNCNbkrMjLkkTpokE3Jr
Mrb7ZYmgfFdGTEBEmxHl7OxDnWsURa1rXNKUf+c35Hbw1/54FRo+OCrCiBcdFAb9hEMwdJDk6ba7
ad12AZlJxbvvQK7MEyvUEO9JFAxGdWFlknIpviZW3s9bJofrpCvXCcug7gA9n7bYQHvkIOBPOnAJ
s3Issi5XO6yMLV//UOWn7sms7KtWL8MgjQ88dfgWGgmZDAx3V5pgM5aRZgweCYrcPrOrsVv1RJ1L
CZ0u0dFoPRVXeq2YRLsbrEMWAMnmFr0i+drmTYTRCEQUTfNmSEYEoq8Aur2mvO12bYIL4ycLO/kt
lr3wzrJrTOxxroAwp17uct7fkd24/5m5U9Bq8qWju9WkELSTm/feOYhy9ORY84PmXGiofJZ60ZaL
jcdEpnvPBbfOEMEYxeVOjD87Yg84V1PSXNCPiIg0namgxxtyw5vDuDV3TM/U61RoyJsuOCBEaNCy
chYIXeBbRmaSl7/8AMg0quKScG4cyCtyNsJ/tHDJumuI1vczcNJdRNReeQMPq0N6bQ87wgPezcdp
/nJkYVMh2Gdcz9UlKEjnreuxC5XqXpz01d1ES3ouiqjJO6mEqGwWU3dhNnW1odXrJFdwTNh6VpWD
32coOZZbywqVaxfa97ZN96xNhf//5gaHVOrQYHkmB7v4fX4VzqcIWu3u8v1NcOxUg3haeE3CzcrC
HESPQAdpb+dFa/O3oWUEMTGk1748lZw1dsVYLLeclXjF3wGlw4+B4DbijstFNFjXaksUAjD6354d
DyOLeOCdYIkt14jtfnBhFBVwh6vU/bpaBP2+SOffJBbHB1OJahxD2Bvz09GBiS7z4fIoUYtb5hpd
E6ZwZGuMVbHQrtcXjOpq+il887wck6OtHcrPjXBWzxcVoYxVr00Ie09kEOWCkmnHn50+VWEYg7yR
otxW0TQNOGgTIp1qjtNFoMGrHxYFD83oQPzVn948Hbz7MO6L2zniOGDLEC/Q5X5DCtusUtuSzGVb
qv9PVB5s3/JhLjP8/lS9E5pwpteaEPlMdOZp9ss6Uqxl8g+2/HsQ961iG9ZoArWV5UOI60Pxkzwb
O3AvKUjvbBQf5ndIrHOGHpHdIw6iEQ0AuHvauuHlsE4hF5bjMDiJKnzVhZudnx6C8xzGzdapqYrp
zV87/bT5OVcIEnJLc+s/qfSjdr63gykBel1JwpGlp1/aruNPPJRxwe3OcyUms3dDOLSr/uvQegZ1
SvdLwmYkxcsfVUWofRsX9iiHCTMDFNgm4Ij5yOa6Vym/OG7Tv8T31hf1m5nLjMVFQazUf2xk7Gbf
Iunng0y8Vol48wi1A6WsAbux/YmIMTa+T+AsOVkkHDxYfvtySgjbSpTHLnB5TkhEqMklSGKzd9/t
xqIo9mVPnhUDc6RQHEo7C0wmhnGnYCbku8CXDODgvSNpaFkxNv8CCFwNAqbEqjpbWUaUsvjResoz
QJbQ+KZUEpkfEOPDypHNaklpbeEjwZMH0mtwnvN1QEPSiBKqogM30d+/WSr+ZS0qDNfkidG6Bfr5
g1yV1lUOOGFpi0bn8j+dhg03Q0E0OUfvrE+EQixTkODx74NqPXPg1Ia1eIftuICfWr/mAQJ2UfUG
Z+Vz0K942rtBVwDYevhbqf5pzfrLFPqmNzG23KElt2QC/TEtOwITQd7WcR5+dA89N8r7xtlzT9r4
RDRgYVsNZZePIPdFPUy/0YbtOBPfswhTB1QVUFRCBkeH3A9wzJZz96JS/R4uGAvZY1/csi2J4J0j
L1Kj1oXIpV9pYvzW4zutxbERYaEnkDzGnAq7jM+Qxb1imAkqmP5/vfsIxp1OvMa/GgqhWEYG28Vt
clRsTl4o1/PevA+u1DjzVEIWGOR+ruFYcW6f9Hq/TvCsefR6P7RKgBkQzLheJkr260MLouRHa+Ws
FQJmiNyrKlUKCrJGdhENhW8fA49UU9QquOBDVXQ3m0Y0ah1Mqo50W/FLlN8y719XsEu8uXaQAeTI
XWDEbPrws9Va2vLkWjSuW97V4QcyLV1fePE4PfQzbfBdjIRKkWLO1vHHTXJHEZJg7trH7Ae+33//
YBhOSUqdxiXRvuPTpZsuc2fftGpF6z+ao0zuN/5o++C5h9DTWBD8Gzld+MLWc12uV34M03BcxDOF
lfH9N4xJqOmMunngx3DEIgSuWoEisSQg1CuZ5JxRpTMIoqUap8LDAgd/jw2eUFG0ZMd9cNeInTff
gOIGP7IWfDU7IyivpKvprzpCwwLy4MYQIUkAmOygDYsg2/gW88EGZu1efcKWjPpcq+hkrXLEcLRi
2qGq6Z6XVCybfT2nbXph72HIgMiPvrPZGBoxk0RBPzTi9iCrVqiSfetgGRQpyR6geREfqdQRnfzo
a5d1eTyi3E+Vns1aryJUEzFqGLT3H+QroAJmXwOhrdpLDIS25cUaHbKiK27nu7UwwNd8X9XYL4kD
jUvEA0/Tyd8Qf7mbWf/l+dppXegTd6MHYiU6UI/f3tsSTve3LbJ+3ach5YMba4v9zAQ659YGHODo
2/i+EUkya70Yv/pI2sVmymgOsYr2ipTcWp3eEfjp0Gi6wSgn+1z+FO+s6i2C5tY16sNNarcalgUB
zgLRrF+fYtHvboMxXQNhkcyHAYdXZNkcwx844olGfCk6jX/pSKWAMaJTmoD5FUu6fTCu3OkRE1eF
+Z69vFRfz60HeV4WoaFK1qGy7ceNv/J8bZQC8wD/YxuLHnPWHIkLdUwvEB6VjYChkInfFfMhiOm9
WUnJ2ERCqJft+3kYpw0+urVxzlfNlSi01hoTiqPoqLzm8238NGWK2QSZOFbnHbE8PHnMBetjEuLG
dbMVU2Y7WM+YQWLYfeozMoKBCC9Renu/9w+8oS/EHG58oBriVj9YZg1qmlNmT8SADYA09AA0l4co
2ddueQQ8h5YtrUn6qkAs94xUwfmv0CFfKYXDkKNhuvu8UL76dzrCj7tyAD5DEBr8uK4Lx42iDySZ
MH8GXn5pbXoAx5RnA7jtUS3c850GtfKdKNsoNjQ5aSYi9ArKgrunEwlOwDIj1fJspJp5Ga0npCl6
3/6wEvzJxmzrFRlzofpaSSjFlo6I48ryW7cc1HqSAwfhSDrn66HS2cpJu3tH3UW4DDwFthAHTumC
dkHJU9ibzArHk7rA02bjKACY1Luwrkno7lPYIgvb1aUT3hV1LOODcq5L02GthiJ5sV4n4nZReTd2
dvO2prMP2k/90Hxy23qzGuxk//r4uTy71dF6xJqZOUgb6Y+7DCTncVM/3EmrL+mPK4COk6bEHpWZ
VOqm7GBqfEx63CN1kj1rnfI1iUtFW7knM89yaYn7LtDPPluOtOe3Cq6roiPZ4KrKJaE9L+fK/MLC
TSPPOmL6OU+TjBAbhkd1blVyhiygOz0TgX05Rh8PtYVOnnwZg+gPxcPL7jpVm0DwO2hDOakS10Cr
bYkiW0qZxETg6QFMmlJo1B8PfSmO9oIFRKOSELqRc6OV9e1HI1jZGjNtFOvdR8P5aRV9gWnNHIA7
lEpHpWWbJscVxRBeP3c1xIQTrpQvxBzzxTJhvKsVUjTUdVPjjxEgBeywQ9vTgmtMaa7cNHs/YLMT
E6MTiHKXV3VcJubEfsmcmHGeL0rmnVoRm5I7cv4YQGX5SJ2xzzuhiHdRjLuj1q28LRZWLAjAHrEx
c0dAiqWusobZJYbSBPaSJc7s3KQXbS6sBuvo2HpsGypJ8FYXxWOgnzNZzeBkmgrVtJ8dz+cOTfwz
py0dWjAldhhYDavuJZiMOMpD0ig3rpdBOcKZo4uzneTdS1Fvb+1Fcitfg45I2F8ezL1xBGki/rMj
jURwg7rRN+Lz7ptLJXTZEft8yzCXi69gojDUGgHC3o82aM/0kWrAQawQZ6UmhPOg2lHsb8dfq62b
Sp14hFwPxdAYvN0/bDJune+yqTXVYvy6xrq5zaFIC6LT4/W9JEYnvTMsTuE/R90QOiTbCpstXmQV
4Oj/KxASwVmGObChTwYo4dawY/IRAppkOVN0Feyqj5xrqy2nLX6LAP78HQugQz80MHDvpeVG9i5i
4HiKOn1AuEZrjQc6p7iNPGqSfrE+cvbCixKRHGXaGf5spIoA/Pw9DovLmmS1q/eg7uVXUMU2JiS/
hEQEd+voobNSpKFx4GbIKHnecNFjRZCEUGfMDFBubdBhI35m9KihyvI/Tg3+AzSCXNMjxqK0LZli
BkbD3UTcSybWfE3ZM+85+Y98x2QywneK4gkIxbs2GUxWS+zmP/IP8WRE6FO6SmF3FMwQFFtN3nQt
p1J8/kfQ/o7B5LE7fD0au+gcgAr1aiaR3S8+fanHVI37Hv0JA7pRohKyDiGBRDxQEYgRXWBYDdr7
Trm4ke6Zmi/sAAxuSMLqVjMuGxlVeuDo5EZkUZNl04qApfO57WJaT5AIZiKh8EtVAqPcfSrSBIF3
inV2qWQkCCF5+6Qc4J5VQCkw9DheSQK/Br9jujsyb7iWvSdwFiScC+vJDpwJBDfTgEEgHPl7eRg6
PqrGF+gd1zXUwhl3BdyKoYtvnCb7juvc6X2AFFHTm8b/nHZVYFafKoTyy+NkL6DC15keeTfFnplY
mLQIMT8pC9C8eNtfmEFSGVdluSWw5alszC8yInLDzbM0yiHQYsVQOtHjik+EcgzVeNljU35spx1L
Ces6vNaU9lvtlChlsIKP7ZKVbKmGLKRPNQUNVQnWj3hPPwLKz5OhOwASCDPZg/ECDfUasvcAmVGe
/0XHgRACp7D+u675k6TxHS9XBwYJyrU1IbG+mQPYZPloy8skORu72+ZLQlUfsbFINWJGVE78kCsY
13L7F1glI3Nu81aIx5xKScVTSf46+0yvJn5ePYj4LCqKdokMwT07lQAE9xtbHFDqx9YVt3qeWT++
DIpDXrs8f2D+b/4qlSxVfGIKIRa8alQ4sVAfM/QLKUl0Dc73sZkFJUBPPnOnEnn3LJ+oDOTZF4XR
nPg6VKCKOCG3Bmybn9IHpB9c/vVse7xjTruKnR6yJxjo/qFBF8gCjc5Oh1ZqZvEzDz+yFxTt8v25
DfCRl3zcuE/qDb0mkLs8T7NKBajGRbvQIDia7UsTbCjXdYagU/XYyr+456XXFuWj9MgFGBNHrCVs
AarwSVBF0E8PNA+805HL+RzZrzqKIzVI7zNJRI9Rab+yU0ufeMnh446kWou9Sli8ekyLNXJYdUq8
yYQzb7f0JF5Xi6wKnS5mznk1c+8mBD4SmRzhE6b4qzbQyyAqhJqvMtBETP2pWNkB+V75dMnrW+OU
wG8C/o+icT/ZeVZwDA3mHMSB2IQer4noC87mJNkGoRq2lBOsKTNUl9PCCm5n8PTgTh54dM24MY6B
Y+o06cQV25zbIJd9YMDe4uHC7l0uKgTVr4C+ijoZnYjo35L5g++uDMnsUIOMG0Dp5OGVu4VWfYpx
t7dOuT0DSPBHwrQR1RwVIGYKmroQbnmCu84eBUNoI9Q070+utRSLDaxdjtwY4n5bXtvTXFrsz3t/
qb7kI19tYyGVCgKj4kMNEDRTIPWsVvxQKlkh95KbqaY6yOh014tKSjZznYP5BOD4GhwgIqOXTmPV
8TVY/rONU1Hg528t1ReOov1QxiXMPwAC/Ww3MRy9u6wyPNYcxcwU99vlJMgngpvtO3yjr6d3dZ3O
BmgY5buwVxkE2Ex4Sqn/OI4B1xQm6hhKH7NqNA6OGx0MWgUV0ffCIM1zNzfSPhE59XKcuCGA32uS
lkhjq8Pzwf/iXAAc/Md8/o7umqQubOkjzGNu7VbpN1p79x20Pdn+QifZt7AvtDRhxj3a9q6o9knQ
U9FJkbXY8IAMpwkV/sUg31Jusvm33Txd3Z3C+31Ru4l1Ai/3XrdOrPOJ+0aiz/zcJzq3MazOfq8Y
cRcT8hAEwI6aR3oZ3sppwqDU5i7ljtte68BOxLEWMkadyrXqAXWArz+tM7tM/x6qb31WgVjSVgAg
KF8l4iMnJ8Pj3GTMyNKL1U0OPdRmdxVnpWm4llcXtg/r7fbq0fz98Ow2HqtfVZTLBj0LwbJXHNn0
80pQY/BA6tfeVa18hLqIOvjgzusPgOgndzWst/1b3gkbvUKmRVRMyXNAUuO62D+SHoXRxBU67NGt
Km3wF+dLR20YllKjFWBws1mEY+NLMtI9MJVOwqO5k6HoLbqYbbZs8Uu8puaI6p+gyZmJWlpwzSZg
1S8KRzLO7bwbJkyfC9J9R4teAlyGzQsgN6knQLldDEeIo2JzujUlCIviYDLQXOllbklGIyTSmRjw
bOqRbCbRB1Vpmpfv+Q5YdOKCor3aPADDccxpKie/dwl28ptjn2A14h0blwGGn+d6MtZDFn5ISni6
jVjze4mfnogS0gJx98XDHdea6UFEsS2Y3a6a7vnE04p0zaI35iolWZuKMF3DYg3QlkrwHwIGCg9f
vNbetFd9UqjfSDkpM8O69t7/oxG+4qJx9eNBKmMHn7JjOrHF1LcvafF8mUbPv0hXV0VQY38iiY+7
eR562JDkNVI5HfnHyhSgiFBADS4p3/FTj1WHXOVhOZ+Z2Bf+bh3PKbc1DVYLbz74bt3KOazQisOd
QImrnwUlYajwPVkRZxc4kXMGBbxrlWcRIBAmQ/QU6L2LosKN2vWeNtZ6lfDxYDD7H9uygBzrIgNq
6OGSvr+hcIkfhFp1LBltaVzVuGJaTA+Sqb04ylLIkRhIAyxqx4wVTy4vo97CKsCCArGaqSb3mgSI
5jRXr/JVBSX1knjDpr0OmVqcAhfnuunlflzd8MAUVJL+MdcjuFAy8TxwoDtigsMwXxI+8yUqLBBG
sRq7n1ombY45ubUGhtuZkC/sIrkKfkH9szcSbSpfoeUZMQBNMHwJ8gYrR2FCCAW1HSx/nT6p0DAg
mA+7YsWOYc8/rMNG7J2NLywRvjYal+Ix8w6YJ4KXaSLU37EACZuGlh3LTZJ/3Y3pj5MY8SCtvHty
egTYzer4mMf7cM5GFbm070VCXxMVHu6szdZUNwQU0MWr4+Q6y15mZoTtfrHtXQIJXDO0LpgMkGVa
zIGuUWenUij7qKqTgEfCEQTOofVSulmXQHWzMVlbvBM7Kd5F7dvNB65Jq9IrImhtxhHAQCMoBuLp
cHgwW4lUeJivfZVvWUifsqpc/AU17wRwwYDMBm4+KJKX3neQ2tcm6lvp97clk3x3H9y5zjanJyNG
XNNMuqQe5mc+uMGgFrzoLc7GXJA5dToK4o7ulRDA99aUXjl/m3Y2h3eQ1FWbqYPO7mRReOLhK/8C
VSivH0pHvcO0tSvoMo0oVpia90jIi101m8BJCsw+N+cSDDBrOktbxHViRWR64e4vuwg9OUeFGHF8
3gFo//SwdmHdOv4xCNZ4+Kqb8Wb31F6rluEIujBtoLLmnAEyE18tag5uqVMOKu36rw8ypH5pfuiW
EZ7lZTuOsourXU5ho/nRa8HIn2Q23GJRdmVFqh3WpXWJnGLgToBDYTD2i0CUkmPV8KJoiniBRSNv
p8B+o1kkz4L5N1tK6PrrJ4+49GpRoeohdJFFhKiQFSifgHikTD3/HBFqD7YKoJRBHgpz7kj9xvEM
BwsrF2KJhBK8w2PCtxbiwWQEpIU2S+325zN7AA8fxTmN8tYqqekozhcMRs5ionSXd4Y7IcJnYtPT
L0EGTPZQEk818QzkUCyDGBGSy3h0iShno2SZyyqHEboYfiRF03zjLB9w2e6TN6Qp6v8TsMF9rUSF
pe+24N1/oaMjocFMuf1rv43E4KmFqfXHzokNhC5lMWG+ww8SW4c8uMPyj17aFny8qyGbzGGxJuZ2
2p4K/z1kTNMkQubHEwuyhSD4RJHl5N6sYh558xx4v08FDOuG7FDa0vRJPhmy9iz3qs/cQkRbS4Bj
JdI6jJctxYOWGbd/GAGB0CVdt+B6fDSTHYLj0NYskPBZzzUN3dJunBXHCyk7iT5pzm5AUoIRIHcZ
UUSN1suJjFhUC3YE+0irZ35vBU48tRqU4Yiqf5LpnTTseKJrIeUHBWDj4p1EiNWo+Ua2DnlU/rBA
JMisGF1Q6YCPzaw17PPGhwlx3f6P6l4a39kStH3MpR0eCBYo8qzokwfihvpRhp1HiMC1JJNMNMmz
0WSRw1yxeCM86n3sjPPR6VUzmCLgbY4FEqrXzefKhElU3KW6QJc6LKn5c+/Z6D08WLeDXnad/Xbq
RvmDeoPGOKv4UdPlzFJ48+Lz/65BJRdSxJJ4Vh26rACNPrnbCDxZwdxV+CDpa1Zq87IkmIKG2jK0
x74hlj/kRDa24fOMkGA2D/6sFlMlp9JSMToeMPmeeVHrT9pByDvM+ASSc31rEH4j2kFUTvRnH7PY
lelNcP1lR3vsC78TZ4MDcBVS7ulgAHQ9FSa7DBT4LAETqdhyeSeG+XrLvgjiQL7JXLq6j1vyuPFi
lMQva7jPXwlp09r+RaEp+uYxHR8yxHmN2V6mVbUTV+bb1M5qiPWhe0QGP3uv+di4K3vwf5iofBc2
3+XEW42V22LxL1GMWuIGIN1lnzpwFC1i2VZNsO7L1FR5an9MNF3JdA+Gwoi2OLBKMIMM2on6gcbq
cnedXcc/CjJC7x/k5dhNfGkI2VesYKN9quDr4Uy/atCzU/8Kp3XlizWcm6xbtbg8bLmdxgPKgQWJ
1QiSFPYeXfDhzDcxg4Hzkk9TfPL9LuLoPQxRzrQDKn8BdXXA3PUrtZiymsnmFrJig5xWTjTURTyg
SIHGaGjTOgvzy9PpkPpmVsWwag74xmHQlwWw3Skb4snq9/jHYVfIT5LtS3YN9j6NdPK4wCdtaqsK
8RmbJPEVpVr71lLOxLsBWRXgERhrsy2nwe1uc3pT97Vi+5GAWK8PxYae9QWgrQbtED3Ut8MwRscC
vA6esrOeyQEoZqO5HNUCxuhRLCj794XdsptbSCURBBTfk6POdZjMYNVYo///DFaT4xWkKA00YNO7
35QS74ivXtf6MDZrdbRvLq1RGmXMuFx324YIrW1Fb0BYzrPSJ0N0fO+hGDN9WGHLgtyirdiwwG5p
MWaZJxgiOvkV9X23mG4dK4Q0DyWTXLiY+qcu53JMThGM+XbNcTv7ATu9uzx7PkWjGhHJhYuZqCh9
g2m554+Ef56EX6A04rGI8loSeLYw2cFLVX44MftnHoP2/5piMTMUf/xFipl6ZUXYpUEf1J7Tcvcz
SfZd7vtBOIiyhm7XFVCICi2sVEm1kiLr9bEOs5WN+MxFMeOZZevM5Q7uNdA7TdWhtAeiJ3J7KFaa
Ernsy1XnEpHrRqTPLdw2nfqQlBatk5h8FztDj6HW508Curq70Zpog8imVscixAbKErbVAHPy8MsJ
4caiUyYci6LSaB+hbe3tXyz0wCPtF1pughOYJ3nZYLk0SJ0938D+Sb1ZJLzFVnSBBBDCDmlidLN5
NzvCPAHpeaOr4p1E2nlnGfNWvDd2WpSGrfsmkOzaMabfIQrbyl4o8hZHV2yXSWhR6VvUF95elYOr
v67R8AxXTZJXq8oAmnb7zgyosUdeM15dyfrm5Nhm+wdc7RI/Sc+By3RhCU5Yp1kd2RkxaiEjr2BX
bBo/yyEop0+44yFNZbzwDtWFV3wJ4HSkq5K8cRLBql2WMEcevTK5e9XiLJuVs3R3suCDQUjmbWTs
UuIXl9o0dWYmrsbPECfUKtyyOGBvu7MelGv7p8gJEKVnPXVaDJ7mrNA1kjZll96uwQIVu0sDZAJO
wXdA64s8QB4DuNy9iET4BYvUepc65wbGAlZom325CQLfNQAeGVizxy68rF0J9iHpCDqmt4VRyIwK
+kfwzPpxZBy4LH+RFBvuqivTOqzXzeyPsKNhTQEGo4L/UJS3Y5jQRx3+DwEoyu+nLxUqP2pRvb78
pdg3xjqWGdzDOZ4i3O1ZIJzDjbfT9k4aSWgFU8o2HRHtCs/g+T3Skb0MS386SWSaQ5nkWBqgPBp0
nVsBQ+VSAcf/4nmKFCYZ09ECnHEaDzZQJy8VmPSCMyqZwIS60LpK558E9cVf+d18lzpT5ohKf6Ya
z/678dKiFkpoPAkq6Sh+Uju0z9B75qbD9n4XAD4bxS/dhc3nKc6LNh4otAztI/5QrVmYPsxs5JrE
FdZxUmj5Ht9KK5+ms8q04p90AlfN7CcWxpr1XD+TwRU+jQsltIk3SZG7Ej39MjVf0SDAEmjtZA9F
1ZsCAEctmbNhs8w71Bc/p1OQDA5RPSF28jGbuf998SawpqYw6ATA9xXvcPuckC5FJ477R113Qxhw
6Gk64qlsydhqpIBXHyZ45d6emXuP8U70QlEJ4xoHchFcyE5MeA1ZTFbzMCrR0IY1dIyEHLaPPegO
G305uMVNzs4a9rMqBTQt2dV07Aqc3ulo+i2yuOpewpfQwphWufXQBEk6BVYKlbAbOEYmu9RxWds/
0vQuQWWIZJv/7Z+s/RjSJ74yQ1jKA9lw9G6eOvSJn20q7KG6S7E0dmJDcFITY/rnyBiRRxh4cimi
eGZBS1SJpNTYTqDNVihf8D6UV6snpn/igrfFxkoP95w+6B9JlgPajwc2I99xwPoeorwBgqDkZSQv
F8k5ZRUbLSHVRnkWAiQ1W+GO04VTTTJFpWV/t6gRS3nrxDyS+38Y0Eqo86S4yARAW9P5vIOpcQRn
WTEA4w5/GJtjI/3Nd4z08oOhhaYD2NJq2tdHROLdauECN73tKIeUnpVz2zBUdqOedfd3J6p73Snn
26XNLTVZAVyOyW9hkBJeGFcmxsh9bGMZlo6RGqBPKA8YyuBnYs3t0idAQ2h/mMeWcMHYJhDltNnL
YU5sUz9uB7i2zCHwyz6xz1A4Zihos4GEsbvEW97yU+GMzYUR2NbERFPKx4h9FuVOYkGaCQ4xnTdb
3MBifCOA217YJAbj9IPo9AwnR+sS6jrQVsyd8SnSdS8NEFm+fiieziFvfmNcqnu+jZzbIEdxkpcY
eibEaRdNMmJALhVPToUY+Fbq5hhfLvIa4La2AxJDljnYfYHfcfOXbVDsm/CkrBuwUuZ9gn7DfTay
YNqEo85qDYwVVFH/hQAt1GqQLV2OwzLLGvP9unbZOAHoggEFC++jsYwnfY8A4eOGJNyp/wqvnFlk
21WWTkIJPkGU1ynsVZasE7CBgTEAcsEABhMxU37Tl9RuXx94sPUoAYRvo3yVRuFxQJtiMmWNvZV5
D/PM+Wie7yLyQKk5fAA1hXWvNL/RRtJwjZ0BcsSs69nvahY/SEjwwFbsNizAtw8T351fhwg56gdi
l+zm8xt7QMpoRVrwwiHjCOgK/N8NYEkpWsIuAFrzdcGepRYzgM+hAQk4n767xzRhcrt7fSi3VcJO
y+N8YVXo/UYQWCvrVv/r3Gnzhm4B8hWTzrEVzMIXoTvpwKvFXLhSoAYDr94LjgmphylxQHenWrZS
wKk8B4Y9PUM3bjt/gcFaVSVYGyLLgGk5JE3quBF8T49E3mvgqL9cG5XWEEiQ+B3dORguXPeSFVsf
MTQXSZs8R1+P7b4aCKybwV9c0q+XEMOYOjFfZHOa6v5fVRPFRY2frLYOIg8wpltbqNKWSWAOd8ly
vtanOFTplqGP4CtZKJDOLgZG3TEp5C+AOSUnJ7LCvDjgGerDhwSJUdenyRPXAHBTcar/9wjIdwh1
ilDD9GNMYWazsXRn2SSlChjy0/iu6oyhM9NdzwQvWs9x1RszXIqts2zs5eMq/tpADrgCkcXFgx1N
Gb/2f59wgfWaWyZfcnG5ZtoyQ477g980xi+DXuylDvgmQKZOboKKAZgeb2w8Ynh3L+Lp4OgPNOKE
QQVnshx79vONQt1Kvdb7kxlgXLrTtoBcMSdi5jIt/rWi0Ye6qJ4Hf82sK3Tgt1/yBryvFwAs0HM7
v1KLf/4+vOxq5SyZkl12vhhXNoETabtKJeBqm6oUmlmB3Sbli55tHb/OS7VCLPuqMos+SaPcRY8a
/2yEWzfQbl7YplADPBv+QtP9yhICinqx062yYCShXqvDNHhCC2eju+dd3B0ga1YA/kejryh684Vr
aKcd1cp6c7131/UM5N3+OZMIzIbj0uUbILnxVbouvT8snvSW8Zgn76mdmlJRDDEOjyPZZN0trfAw
Yy1hiba2g2HvLUMKE4yrND9CZrEsqYs+JLhPI1R0Ctg/jsfRECyI5Der+KG9xJEcY701n1+q9/Yj
YfKulwkNfEhLDoCsj1pUWokU3dQJtxh3CJT6vpSK4xiD4s2rgZxoSf10tsu5oapS0dJd1JmSaG2g
m7PuiumbZCeM7KLx27mREF2FEMMU2xOQbV7JW3HMkpgwvZrC6VPLBZc8nSy84GTNefTyS1A4+eEX
w9cdlyU6HO6bBYZkoDmgrxOXhwBGwQ1nIwnl1KfOROaFYMF/cbNZXmOTcmOcDW94HbGaPw3YtdJj
UUbD+rtixRkWF0iEaeiQJBsOx8qgkbXIuG/g/JuE+OmKv7UZ6uVwzaRUqYvrP0AnEw4KMq11c+BG
8xU7zwSsS8AZUOIgxxo1AJrNAXuVrCIPuqK++NAazsr8CrZ+8sWnVa39PxpcU1szn063PMOdh7dw
1M2P9ozTFjfITvk1ErkETqMx4Fgu2+4B63sjGKYKWXYH1mqOrKu7mu6bm3ux2aMpxqpDpMCS1lJo
6GqZBgXuH6K8YTP4qzCkBx/UDCmzRrXIwFBVX2IeD7yVkS1kvIDyuJbQmBhZ3bX1Gzl8nUaBVL3q
WSNF2YopxDjAbVzTu7VZFomU8XESz1q1KFfsVnS+6L4tQxI7W4ZaCiZ2trJXlKiJNUBwR9QWKOZU
W+KcYvIKPUkm2JvkKM4S9BkGrkpHP98xJds06jYh9LlL4T2iH+zuUse+2m1Y5KV8IbH/T+sxXsdQ
w1piySobro+BYVjslW8raCabQpce0BS+9PUdAXAu0nIsOaxCbXDuauyeHitdok2yzAp43QSww/Wa
h0DnzMk3d2DWZBptYs9Mw0peSLSSoaI9jx08MZXAUrP2wWRmaJt3UwDn+ZzDDYaaweLzwKn/R6XP
Z5jQNZzO6gEBppucY2OvcdpG77+0CYOSzV9RwRZsITdlf9GRFx9AU8zapsDevwv+QBa9NDPp7cnP
O3F+2MKeqCrTX4v+fPe2MF4Ub6+bjbhtZdAEbnCbUe61qGLqjd5bPy+A3cETrKMqVc48mP4UlOQW
PykrgSuq3N5msFMXdFtFWeRYicHnaf9yCQHU65Ym+BAN7wZXA+nlW0TTgUw6kgft/6+ASRlVeAPx
UYoGrMG1GFoxIcb7LuhjOfnFYdrFMmZ5oh4Eh3RXDb9G5N1jMZteOprKM/v0EoOovbysfupn4hB4
kH33JAT5ZKt3lalCKISuo4BzlOwBarBxTnrNG5huu8Q+PtoloibGUpfyOep0A5qVObqK+ax755Xn
XEoq7sLGxW6M9Jb5RurqE1/TBulwSsP6th4EBaUoRF66cz+5TEctblVsQ8kATIhbR8tOdkCJMWnW
YgDl0o+kfCT4xdFLwm1Pn59EbsIshae45l4AFDKOXj98dRBg3JyDpsTKeQNOlOqOMFM7F8tQpJ8o
+m8SS2S50ZJ4Q/twQHheOQQ58SnkjW0lGVpzz3mOKau3YlN2Cmb7ZvD+n+71Qzn1FJ+gaMLaBbhr
Kqvq7jSkQJuj8CgqqVYyl0oIzy76uqHL8ljMhXSIavOtCwth4S9fKE+sxiEvkDYPEkXUn9p0hqYz
ApUyigXFg9DQg0RHnCd1jyVtEeGWk89oVcZHyeK203l/9OygyZ2KHL57+dbHVUQS2k0wtBzx7Bd8
rRwOJbpl95wnQDE/BfJaX/o2l/3vJj8NNcJMYqpL9dmxDYOEcKf7MSWiIP5ZOZf1uDcyb5qsdZ51
e6BGLEi8/Q7ONpHNCq8+vCa65RekFbvpw5134xQPbrVTC50EDuKn/iHbRGJGrNK+4NI2w397P+Xg
xHGz8YaGoRYGsLdb/zgMzVnaJN5cxtMTo4+6X2V27cS++nEPAe6lqNNhCmmK1aaJDOnmiH41f8Uz
rpwOSVrBELfu20jXVDg5iPETwfiOOThuncA7XGZuuK631o6eSI3oUGuq2VwitEPD+Vlt1nBM6gJB
yQA+OcOdwcVqaS142wMOdzQA5iJdyeEOci/oTj4FQnC53JuPGuyXz3mV+gxbL0OTiRPE0b2Xjgyk
GHn7mgkQSG5hR4Vh0Wg5BY3FRcp8SxMSylg/3//TziuD5ilgUJ0Uwnumj0WFeXc7feExBLV35J0o
kAU72RAzfX8559QKqdOQRX+FRVknjrRwzr4rIt+jmZnngk26CUEAp7icxo8ke11SigDtIshpg3nv
9X6WKLo3RcPj1pm22Jhia7xodqLJ+JfUNVCAVeGcewmxaZc2fKmK1/71g85K50ArSuhwKvUy8TmA
UyIFJR7WJsJTKGK3NUv9ka3qZ/w9S0K1iiM9axK5K3inL8KUlDWoQzXOZM/kbXpwtv/QAMHdE4HE
we8e2KsPC2r5asVUOGoi/2frEJ9/3v8gfkR9GszJIP5tk1fmfjtm7cCqPj1ZJHfq3BWERItecA8V
PkGrEsrF6VBTVH+V6Dsa112O+zxvfoGjSelS+DRl7s1jWQEUw+iUSUZtafjbIuGMHSCfd8LPE/t3
sSn9sACXecExe4A5iid1O2xPWuN5EPZqAo+VchlG3yDaNkRXzEcNO32OzdAl5d1MDoYhKkqm4myB
HOlZwooMl4t7K5QDzfjDffXXOUK8zEsv30Cj7YKwNLJ+bloVRNAh+P/g6cAal0eXm24qnkPQE3Ug
hBp5H92vW0/be8/ebtASbJV71Xg5kInfjCFR+xElMskrwE0q3v64maNhDI/osFwAJzVu4haQ4fRE
JAeVtobmyzaswvX2uR4gAcXpq33mdVh9Gi15BccBfoDrZhJWSim34NbnQlqfN+O1DI9/NSHvlqfq
gepLFvS+anUbwheO5gIUo59PvS2SjC1fBsLfXVZlIy205fAdP80/1vIewUzDJvO613Ofcj23TnqM
SQrT6PYoAOmFyfui+e2dqJcf5NU3q3MqqDVd6W0AjGgzZzQUWn8aJMIEy/c9QBxo9w4VHQGTq1zD
XyY85y/ILC4VwjBzrwjCk8PMH8KYn9hC77DhmHVZwXuyG/iwB8tEOcR8QQU9V8rl6vT562eUtrRw
g0Brl28uCn7ea12OMXZNvhw/nXcIvMBsi3Xt3vqnHX4t0y6UYQZXSQIIGw7QEa6mXsmIJO8Xf9LI
HNpxSFmWa/3aKsmTMTVJKf/nsWcsuu/CnxMpsz3IZn7X+tkrK2QdbRi3kiYOh9cTAbNYTrm3rP0+
QjLfWKFIuSnSW101mAR9tSqC2DGOQaD3Zxtr0m9GCmorV1wnZTNUjPvgbUNwyASmagDAxfDTd7mw
j+TRnBa+wWd/wXgmjEgLal055lgobaPfyYfy9rdqI0kgCOKLTdyCy9X7lpvf8E0E3zOVeZUV7iSt
pBXa3zYNi4b6fsl/owAhw64esDTfCTw1WhcFbOAzbgzgG3IxB9sbQn9Zwd4BGSbOUL+BQwvWww+9
T+Q5RpNMI1jilF0Uj0/VXBCCS3NguTQJRf7DB+XLtPA7duW7oD8LMf0qLwzAkslL1CqzXi6g0BGx
Ye0JqtySkclUGMOigKiw6/r3+q+8gRUk32oHX84wAwCNIVjymto8VPVuphMeq1tZTNzbqib9l581
dlER9A1RwZB+nXTmQsOp3rNLxc0E8si5KFIIE/qT7Tquri/+FEQeStRmkjSQYu8znCELC+iYkvAE
F/CajIlKH25bZHL2aUTOMz0GZbZDnIBNe262mN5PtcMEcxvaaWS46/7lJ66ZQUh8ZUGIZkyGllrG
VdXKjzHo91eG3CsU0koUzynsTMYKkC2b+f2IUBgzeuo8R8qmoKbsJvp6nU5OYlyXZ62FMGinZv+/
Gi/8CID1+xbajnwfL9Oe3CCOgNEUFUcP385QlRmQJAP/RqlNVa/SXpb7azLeGQq28ZKT0Wef2EJr
GbHlrQ1SZR4PwR5Vptgh32YKyK6tgDkGu6kdjWFxsmkyPzv5eBFn1ZVaNPja9v9CHC8xQT6LoBjS
h7DvRqQgnVFVhPNDtMv2NSGotYU8g2y8FLR2axnUiVEGpLSSGc7R8uikHNCN1OYQDNSVYHlnT+jN
iSqrAmKKcl4z74vX+AVvy0DA5prKb/G6SbQ+ZwqgBLAlO6I/4zVRtPqKLT59VRIR8TqeuVo2FYvs
/Kz77z9E0CIRvoKJWNZrbDep5MpEaw8e9zzrwj2tBusPHdqNDcqjyVJRJL9uOG02ljvCvrrFlnIT
ojLeW7KUbMUKWTnnD++bj/r1XWiRH49FGmBMK8pZkI/9X2Ik/2FldkANVZF+QRn1MOd+zblk7nMo
og2ReCqMqOE76OxUEIts8FN5/C/heXJo09H3gOEaolOJqU6LoZy7/USMuo64grHhfvpegH9Jspri
2j0VCK3MgLiL2/UfJ9h/u1FMgNrW/0CRz5dHuFrUQdB0U4F9L/IMDia2DmeKPIzARihf4I5Dqo8z
RT66/nIx1HBvxOTUXkEiwgw8rbtPLw3luXch/j99Xt4xwywoxG0D+yS++cZ3oVFsuv9+ID7517BO
T7zSwZ8d/CpgBnBzcmLrPSX9+X0i8+NweDLzFgrzRCIu4VtpyZjQseVHmmCERNw8n8MzCt485U75
IETH9HZ5VP+Eq/2TqsAgibBWqUx5lyhBv6pinWpFTOYnICFnmiAUpEyLGf2+AQmLVKF2HWS6+lTQ
4d8QG9yp9Oz8Krh0qQqojLvF8msUGGBSkJ7bzPaBUzs4leWMEwRS3C++RbsNXscTOxugE6u28ilx
hkhXC15AQxdFPRO/5B3K4FcS8KcHbDDqFGEL7dQImryzG2GKbjsuclf7GoGnxESnOr+gZ3Qo+IUV
WZ+6TW75ypfBbmNXl8pe/Tz/A7rk9wXQgkXYgNQLXtRx0wc6YDKMYcnjqxDb5zUfVLSNWDp0VqTI
F33MTUw0KCcM/6dD2LOrlQStZ29b+pxrn7RyRbqBMjykA5KLiJk8jKgeahwent6uCKGDSxDHaNYT
jU+zc2wtqR7LvkXevNXeqX6cBa5VpEj0d/MxnJqEeyL60hh/fBOtiwqY9AJ2LOPq+MowsUv5IcR/
V4V//rZLRJmviG29v05ldyPN+c7p9vIpZ3zz1+6p7eLdgrA2BRc99VogaMYaNn+YXNlQeoQiTOVP
JJrFnNYmfYCBQDqiO/mhGoNTV5N0vUraZsiwtuutM3POfZAOb/uFiq4taro/IQaEORH33KyC4D3u
w+lm1cMoYG8byJwqcW2mgCYW9HEJ3b3THdsSdcZLsj/w/GpPHabRmNwOSYgqfazc2mT4/LjRcYrT
v4f0vl20x7Mc25PBQp8qdM/RrpTviQU+vu2JCNhnt5UNKIGvEv6mNGVzPat129OnZGgXFEd/0Wzr
TU9/O3qNjtphw+XGZXjpnxh/sPiN7X/L4SO5uZV1/uXzHXMSyTt2n/AtG4X4TsRD0sEJgEAhbVzD
ZI3Nix2kSiWeZj9yZVr7mze+n6ZNZoRGjTz2Zt05szZRh450yWKmVHRlJBUxcHoeeXgdto1ZG+FG
zYTGatvxgDKEjPjz+vMJwcBfkWFiyYAaUtXZbhY7lo3vPjz/h52/9b7Ruui3w9928daDtCkO9rUd
odta0viBkuf1F02+pxu6yv4KgH1B5xWIwvPTMNz1SzOgmmXsFoOqeItE5h4V3iwLRsK8Vi1P74S4
SRu1aKjdg5CnseNHp/UB6VvvmC9jvbBXh6KmTP1kBlHusF6MQs4zKBHIkA0hDFzaMBrBaw7qo8Ry
KQdRN1628YF+rP7xC2rYVmy45cQs5mKJ0X/HLM2pNohLn0lCfSGgvRoPvSsmoohHrmgQPHQRiYuN
iOwYzzSL1qrPip/hsWQMdHq1hrH2ehS+qHQ82EIlGf3Fztfp6TvqlI+KFcqDTl5dsuOxhePC7NiU
dD6H7IcFjETfYVprpfjwxhaSGHxZzu1fERvoLk78J/p6vGymxhN0jEfpxAIQSnSAPKpeq96b9gbc
8bKxs5BfioUQfnZBkGZdjOOTL6kECvHvleFHxL+AC0JWzI0s9j85hywRIE3FJ9obBq6knL12R8u7
b2Z4MC0G2K8WVGjap2uzTx2Kfs+wao75EPAzA59vWZ26Oh1cmg99siQ4jOu/OPEnZWIJQbivLaca
eflpl9NC68Epol+UMB6/qgLTflqf3Wm4e8917xcif81YeCT0Pk7DzPbtQPea2sbBS4ZDliOPoAh9
DqOW8ivIiuwNooBz4KDy1n6wBUKn8kTo9BwkRKhg3ytA3IsTMA0uMPV2jXYlSdJ5Vxd2XoKDMhM5
V7AXzvnbCGoc206vebd3X6RxC3plpf3GZ/C1bC0TVjxmph6CLdEt2OPKeSk5oz2aLYOsdYK5zwvQ
0cbzKZL3Zo+ez4jHeWTVDJIaUkcU3oBek9Ke/EmG9Qoz07OsLjRMhZ2c0ASSCM3tPL5LAXEIdJt3
nVLayqxsY0q/EpTeRl7+HFOBPXjPQMx89o7RC4UOGnAYGum/yL31+ujPf3Bpc0XFP1Lcv3xetq6t
FwGWp8Iw8rJ3CJsFRGwGTt6P1dyQEJyq+Ek+dhY8LQY8MRnJebfW+04ZfQslPkJqrIJPoXlznWFe
tXFmXSfekeXN3k73ZuXfp3b7CuPRpluTHtx2z5YAXYlscjNtUfabhalrwu3zpISaMVoV2L8SXAtk
uPYvMUQgXV5qKxubP/eiXE3pPCessw5GVWcNzzsNY3VYYMd827LAKLLiOgJ+9lDqxh3ydKDx+RYa
T+tZrOrXqiXAVklULdFwC8MsjiU0BLM15qs+pYMqMHZHjDyAsCR5jJBNqznjMEiPr7Qz80owsMrt
ATfZq0QXXCVTJrJc4UKHfCe4wjrtReznrDqS2sR4cfFm6EJx5+I0Ba2YIYF2l41zL6cZms/qqv34
6B1hQivT0zPHt8PcI4eoEZbL8+Ux11plHNIs4vQPXyCuO3QqiRKwk6QB7ImCKw3FnJPYTKmFefMP
KGspszdzz3kE0xp624OvEuAx+NSHzkaEwAGs7gN21/vWNkkHlD6aF3Rh+t+E13JotDrMj8ze8vjt
D3+V+iMWgthtsVdjYcOzeWxOv2xqTnUYnkB+BpWaLr7RPw9GYyexc5bXri6XaJxIzU39ww4RrUeY
+AqvwWb/w2IUDNQ6I9u8OhTY5Mi6STs53fT+Yd9EfmLQr541w9wsY2VYcsS4vBi8BkjMSeht3Zle
9Yv812Te5P9SvrbniiSJr1qO89KecdZirWXftS2aNWD2G71qKEfImADblj0Q16MxME67OcDIiHFC
HudqJEjbTr+4Mn4l/kgBLEUTYWAsxY8/1U6Ea06aIxqh/ecUZwODfjKwXYJVrrrvJNxUzbh/Jeoe
OSDg76uFj1jVRN6RC+DUoENWvoiSnlxBvNXCEbJ93zmjaNWnDTameePKmemxLvFO+w0l+FMfnTm8
syGNjf0cY7B1twxpKAip0bG2a+x7HRxZUHDwqPwi9pYHoYD3bDiSX9GEWwcAlQXEEYF1xi8WUQne
GTTJJmWygMfKYfW8/u7m9u1E7eyYXhVuyT4UFnGmDsaigXFy2rx8JRip3SGkNVsfmA7jxYQCfvdb
z+OwqQlP5etuimeUYQgElXZMDw61E+b9oUOXw2+ZZVhOJ0ft2dLAQOrMsHfLjUNaudU961ldgVsj
jjgZkt3hcohPQLLD69eBjyqIUOFQSMjEclfy8iOjQSkfciykjb+Fzvyl1j+VsOT71U0Ax03t4waq
if5tj669siIzFAlKI5GsBJjDH8UDcCrqvPpXMC6/eYH8lBbeg9ek1Gin9hs/hgX3IOqtYnahttRH
s33zBxYIWrpHVGDU11Pf9suoQ96TwmNBawwNRD5O705BwxYt1KcrqC3utAxNx/ZI8o/2rMhH1YL3
kCe+6J8aHP2CohNSLOota1OW0f8oa3OmdaEsn+2A9Wo/a37+h9PG2i5aKuW00hQpe3OELXIiSMS4
QIdCYrDJjzdKLi7UkB+MwFu2LxGglZbH35n0IScjc+D1mj0pyY1+LDz5X9U/PEYMjMWjE9QYAA7G
a5xxntmcwuMYmjK8GRzcXxXLQPVHaREbsXKEoeNyqAVj7TjghiN7MF3uS0cpt+LL0pdLf8k8HoKr
PLZPBF1dABOtEVhRCuQ6Hw0OTI07IMseVg0y2VyX+8WlditQzMqGgf0minWa37o7YjXcXUKTp4YK
/8iCL557gQkrKpDRK2op90D1UZPGzDsj6lTSSjtbx8EtnX43+1bXFLATm/mY3nVVe8Y1sHXYLjmE
RcScuKNNh2Vcsgh6Fabu3rnn3kjDWGghbJrYQLaIdURU8BtMAIoWCk4J62MURfXS936qXN3ocNzb
57NoejKhr9LqFL5cRi06dEProJ85IgFpltu17U7QSPlbSL4KFeEJDci9uPiiX9sKfoxWpW/sSOBW
SvGYmQoVgpDur+BgU5lKavNFVwdgoY++XIYgJF6i684vysB0TBde9qwJtnxaZaRAzVSxchpEXG32
9YVJ17NJQKhavsTp9CmjN2/wb+NQPGnKQ6Qh+Tms/Q+kiiQs2tuWq9y8IrJOCwFMSDaVqCXOefw7
5FReqYx+eZql/vvz8afuhrJgP4W8Uhb8QiJGbAQuBcjKz6VCd+hymvehTZvePysJ2nVF+yNp/gjF
2Lm3lRgxfiGHR8OunKm1DKq9UMOcIL0nwHpT0U/IKfNGb77Kao0HQDPyuC++R4cw6AAwoMGXzLc9
XKmabeYUFNn/CA94Vnewfxu+hFfBpyv8xcrWjaHfRQTatZMAkfhi5r+Dia8bX0f94/VzalHToBr3
rLCkdM+/AVFHkQFj/HXJ0jfVW8E3Yg3pKpWJWvVXgzflE9iWPSX0pbQDPTKEwvccc7dH8cDPRprj
f0sMP4BAYRJJWlF6H0BVCxpdBnRDW5LYdDbHdC7TvTPUkY5V8K8xjGy3Y1z2npGx/B05TGeSHZil
ihEw7iqIiXbYFBypDsvoosT6CtznVIP6dpseYOtMadzkTM6I2aUaMoCC5XuGUWOyeesvZgCj2Fhs
PTq6hd6T78uola/vEvDby86wn34rqx6xNTWX4cnijCIRsX3W7/m1/LMrQCaDFaLJ09mnkIV4iYzW
S36f/nNlFmQLo8xD+JsIVGUb/tnrTFT9c0jAihWAI0KLbSbBVn8eeSnwE860ZsDQVEncFutcsBVa
T34JUPCYXeebqjFe1jUuWX7UjpUudwIWFLyiQPDmj+iGa6x/NonfAGvdHa2AkMgAe+L+a1vsSru8
l0aSy3S/T19Bv/yFIRT+7HDOXEYQl7tijyxarDMqhIbBObGopswelJxtm1bRfNFdkKi0DYTsrwZF
+QgQov5xLlJ/PQixQIkikCUx2w5cixzZ1QiFLUkAKRH+FoN/uBFcThGkl0y91m4XH7p6T80AfsOT
0OeRHpzbPH/2AsfMDas4dHzWS2VFppO1XqiZkuUEcmTeE852aaQJ4I9l0G1dfmmJHBxNuvt1uiFC
ZcSUO6w/fWpCGrUQLMC6XWO0qZkFIHxpDOCbPDDReSliQoDENIqO6SdBGliAzOsRCY9hk75THZWs
zpg2tYl9gX4SbrhaBOFFKhfWg792qxs1VSTol6tUr0k9QWba82jUEVUlVfjKrFMtQD+mAnpTYNyD
CXQaR8HcRNZ1JQEf/SQNwLEk2boBn6SYj803BXyXzzBsuYdNMDgT0NE03GOcEZ3bsi7ImAcYdgT4
zrdrl/03FLwK1YAjNjMp0rKouOqe3AqHA8869xFMV/Gz4BcJTZD3Ymz9cr/meFIpXteEbo+Wfv8M
o93rW1C9odkTRcsiz+j7hoKG2H2Osj0me18XsUsOb7OYr1GXuxF7L8khGDqH0SKs3pIlEPFXxhZ1
S8s8Zv9/fGaAuiPzVazeioCx86ASaFc6vr3ckmR9+/IP3EcmqvUVIM5hN4aB70oorNl/0WTGNLYS
4ysqyUdQGtrXnxD4iMLRNjbyJH8wnIa3jKWjiloh+o/IEO2WLFjWNBezRdMJamsG9iO/WgZZJxx+
rV4jZcGUwdhE8gEYZa6c+CXimVP29Oj70A+iBxVnyHsShg5yZtwE6fFDiO+pvS4kXEI4LY1YnbKs
ZYPmnj9sSOJ2CXVuquZdJjRKREM/w7G0bhX9UFMm4sOOfl/9C4gwrmW8wMLjy0izGfcQPaJMU6Z8
DoWK+09wTyUsmsFmx6UKXSqONugI04BBvyaYjiX/49Y1RQdEq7CWI7x3zS7bnphjSftX82YI31S3
ER9LRIYATiT1v5ChhKqDREErcjIrydXry79Nw4K7BCBVgu5olsozArD1S9i5WyczAhCrdUYRNAuj
WH1/fSzqzjUigC0eaSbmISIHmwvrGfq/ofguJWUlNQZe0ddtVy8OS4X+XuI0USGkiw5SokBJOxdV
Q7Fb7FTjBDvEENzt49cLV2qjrH/xm1JrP5Jnm5wYWI00B/eB1xPumuE2/j3YaKLdyXU09hckSxpq
k7+cmdZRM1rWPaC5PH71sCQlbnHPvtk1eXasQMR1zQJ7oXrT1cnQoIUy3cPpM4xLjDhxOIvcTZlm
r0FMUwEvh3/TZ9l7IwLkWoGX7X2zu2rR7FeZzMO/9AYSMK3Ki2jwzOqF6wnnd/nfduvkH0i9HtO4
hJX5MMhfz2F7CAxzMIhoy5jaRnidTdZHbCxbIuWL4RKNiY4s5sZqB4C7oTN6ih6yWebahvUrRRf0
wJPm9F1ewTqFU9cKOMWq78m7m1H4st938lMQWdU/pXFuuQGrUOS22CpmJ/wV6AfwjE1p+4PCn/3g
P9PANRU+UghyDYzHt7E66u86K7UTeSgjeQJdfzdp//QnRJgtwdRzNOhzK8B1+xZhAKXexIDNozuP
I7RzlS3eF5D0FCJTzkdmfRpslNzgZaB+wUc8zTBExlqHuXJnTtCG6mhjscb8A6Vhcv+G9LGE8yTC
IwD80R7tT/9uhVOOdfS3SvTVdDd/yf3jBFrvJZSetiP8wHmzRonUQEd1sb2bUy6dtf+HghAotgjs
nUSf+mv7cD+qKm2ng4R4/B22+cu/rD/GPWJD4JUr53EKDI43rQX4Cf91w0XMm9qio6PcMKPGz2QC
X1Vui6PJHlF7Ma+WWZxqWqi3y0TQb8m66VC/dH88MaOLh7s6l9nnUTmD2cVG09NwrMSwqP2Ne4i4
RsM8DVvwmOmXIum9CWT0/CGiT//otxPGdqgJBKM1YWFO4WP6FRniKbzS2Vp07SLeLiW8uPzzeosd
8t1EP7VN27ZbcmALV1OEKOH6hDR5nU3wrY0xPfIMVqyZU56B64Zq+Zn+7NXhXToL2gWANhxSaz3F
oYCebVEDDicL0vUOPep7EPzJLOHyr/5suVxk46t1XTM5St1WTKf2X4hpC2a8oILaM2JcLYJ4vVVW
MFu07J/GHXNvB+PsXIpt//eNx7v8Vbd4NtPJ23zu8ullVJckqFqSL/LvdkVBvWkKY5GRfBeh8cHU
v/M9Flkbhx45B8h1+aED/3qSPt7tHpQkTg4d+dzqsZsWnj/9YPfLzYoJpn5eb4jyKx2tLs3XlJEK
vI4+U7Vwm1r0rt5GJbEiscnrC6XDMW7woGEsfUyDCOcHcw1K4GNnYOvUcYt6w1ayRmpS3TrZEiox
9I2/d7cdYaf59Ckzd2rRszg3FAZSWmSPhvEHkgr3xa5dsERcx+QXJzbIsKKOlnDakVD/C1VMDd6G
QkfCZfrS1AzN3a7A80u0BxzyHP4jcxxl5naoOJLmhyy1nIxb0auY3JXR6gfliezsoJU5LcHs3iGe
FlX2ljERu3RNtlbqRylnjZJALP3MnRBIgBwQWd/udwWsrhyCalqjM3IS4vdQ3NYZ5CVvahJKuV7e
nkYwYBTHP1f3vbo8+TBu/t+nJwXVLOmXpbjIkKecdkmPlzOsYX99lURlAbmX8k8EWpJfLIRJSFRM
EjM+hKoasfQ1Z5RgY4cFvqRpCFZFjqiYLtXvs5plbkcm+CBReeHWSdDDgV1xhmY2+bE3H98k33mK
ZdHS5MxSs+vBesLB73PqTJ/oUEGu9vjCHpGKZZZP+pPKtPxbLbU5Wuvi34UCnTJUYLnnPKRj0zAk
0ZM0U+2ki1zaZmTBJcqIbutoCccTAIwXY/Xhxfoxcvt7x4VwLPNjLdNcfEbymL+na0p2uzTgzuC2
CsXJ+Ye9OCuXs+3JD7W0YTCd1UW2uCgEXRsroT8j9O3lBNnQjCdp9yB8EkirucpBF6f2/cQtVVHg
d2nmha/XmfT/LuK6nDgIYRIofeAnRfIQY4aUfpHzQ8F7MYeYy+X7RDE1Sba6Jwj3dPb1syiNI15V
LAfBVPRuIQB84VjAqVoSROHtZu9XwCZacJc09BXEAvPhwtgATkCTBbOihP0JX7um2ZRvE2DSkFmW
Kpn5XIapsHj4f4Ts0ZiMmiZEuG91+oa+x/TtlojIkddUYjmGM2pDeQ2E8Y/aaTngRwLpwaAXPk7Z
V5n7G19KmzwYtXIzAbJTaU9XoEY99yUHErD6NuVlzdczGDXxv9l6NhiluUFGDsLeMMRZd8Xa8PRN
pyi5pgxClccE7anrKfoOGWv408sixTNz/eIV1fZdGpomRYuls+e82+cGZR8czp3BiEiBjnZqO3F9
uugGUNEQGWIv9K/IZDyOo18tjy4AoZfSJtdM3JGh/NWuEFFbA9AdDC9UCUEU/etypMnPByPSOJG9
VPdtrtSVZTNgyo84rLP+9kJGqKX0dIBT6mW8MSOIMU0UYj2EAC1hf1BKwbCyzwj4USRgZ0BxU9H5
AFE80jhUR007HHykz3zG1A1uD/fqN82sNtjpM2Z546wX1Be31gfEE/HjJEIPs/azoo/kFWaFb1WH
rmLZ8rk2HEH9TOPA4fHInuSgIofi36r4JfrW/d6fWYkFCE9XlpBzEOAQ1iK43urPZxo915O0RYkd
Che6NhBg99d4sg8x1Pr9TNYM3qYq5Je4Za9jK8tzut4YrJzmAzwDOa/Hilqvd+UEOYuBwBTCVG6i
ec31NgBUu4iUHO5+y48kfnMnAajMOl43HqFT8AhF/WxiPoXqhL8ibPEiKlQu3iINdQATayLk0X8w
TO6eb/eb/j2DRfnmzLBENiOrpFGAD2OMM4KEY65m9OWwhRpTyKaeZsYb7TO5OBGqAUcsgC4NDpgN
pbcuHQKnvR4/mZdXLCjTE80L5y13I7+nxL5Gvqf+KSHRQCf18OGceY9o6Loz4APCn0k8IdHR4jOY
vWb9qg4GjQUt8iGrqpNLZN8t3CVVBdlAIMeM6LG04r7UM3uEmCaG2mszA35LAPa9jnxFW+GgB39e
fuusbj4Yf3gmYsaQxH0VTzS3cuqRlbg2C+xJW8F85KbZCY+KgeWHbK/LFaAfJET5f+y3Gpvh3E+u
aRW2bfbZy5s+/6YCuj0BMwenddfY5zfSRO5xul5sjf865D9/90r7GUSf3VOQdPAURAGMNru8ZNto
pI8QwU2jS028VTTrN6MwPuLyT3LCeGoDm4mYXK7qOnwNRs5AgKp+4CujLNYnM4EeWpyqJ/0065Tr
kKVDP/932pWFUc264TOEJr6+2AHBKEG1GqMrT959PpkUoKsJc1mVbaHvJUiyIdximLU2gn8ScfoL
iWwOtb4YEvgZb2/7AcXfJMAGEyjXLDenA+KYvXObDL9+EPirzEqHjfJ5VM8g3lji4iwnHccYWdRL
1bDTyRjwqVqRMqz7RZ9EkDdzKUAx0DMpadJ3IscVhZ70+GTbQ/vsICqv0UNjY7M+tOUJXtVJ44cT
ydi4jXIspYXUci6ew9llekZN9wWTUMIBR+4tlgq8qob7+hLE5loBvvEyELI6wtzlshW/PXIHVvS3
LpBvlimmXUburMkD5J0LNOhGiPvxw5KlKVq2LJsWzP+LjvpkNr/qQa/AZV9gvk4xqANVdBfIGBNy
opo3BIGv9W9SdET8QZIZ79eMYTSzblFxbDa+Jl7U0xzV2CPBm31FyHksqRvImG4N0f8ImoX9Oe3b
I+W302jIcrZ19bKLF3McxQ1vYY5LKuBYy3mEiJb6EQFOTMRUe+a2bKo5mxzJiRulX8PoxQzMWAPw
ie+fmB2RCSIz98n86I0tEwJxd92tdMHC1xynzv+c45ZAnkhVMHeEHDJ0Bat5LDmECVBTqrcoaXfz
TfbgrW0U2/FtjibPGS696RjLH60WBO2mOyGutY09Mm4jz61+DSU4MZDPEcskTYIVkwKQQVg96vP3
R9WO5Rsaj4dUtW5qBriwMHJV857CEXwypyJQP/Nd6cB7YU2H8wyHDuP0ybOCKD6MF8BmeejooDSJ
/2xtbQ/Bhj+jVVf/V+W6ANsDyidPu5AArts08f1ZHCJmEo8wF4kikvn8cG82Yoa87v1JEY3cHkaa
Iyx1hrQKFAxnfnDv7mudo7qisGYJ9VdKruFmplgsmAvqzBaeE9ky++4fMDd4knHCYkRag5TxJYEg
u0EddNMP4c0nzDV5YIzKf+Ozu4aiER0iMXxrS4JPqqeb12UEPkiT+mhvcSxkpCzatHOZy/5Z/osN
Xdr9xRwPhBWtPBfA+gev+erEk28IUfsF1/z1J1VW8W3M5ryEmO1N3nLonHEBAk3AB0Aqq+KuYGab
5FiOTzuWzw91DNyhJFvH/V7oW94se2XeOL/vqF2sbj9L2EYLep5ruwcReUDoTgJnqFPWxhiZDqxZ
bMMqwQvlfClyd9B62rrOBPNp+QkSGYDImEtPVsiDuKPJi7wZ02qnLlvpvde2Py6ZhHrNAo+/0agM
vUlHNsMuxP9l1Fib2q/vbVyRRhl3dlZW+NiVliADts9L6BHuR68wpHoetIJbBGd+DObfB7tpuUY8
LPAeImF7kCdAckRn+MlFaz1kvJAcBP4dy38IhoNVLhqdfz47yK90eYe3OHUQekFXhi9vk+Q1O9gd
U9bzKFV56rlEQRFkhGJ2ISmDUXwNRM/B+KhIEA+D5j/oYRy2/Qwmq7Ew1b9EdCyK6R3M+I+fTZj4
DRL2Hqx6wUxn8l8ysTV3dEroYI/Alxw4BNvEr16h7f33+6Gma0kmwiENVRUKg0t+Uk3Nepnrkvoe
nu3HoC4uTdcyJMYHCz5JrIOwVXWTj9qpnT/odAFY8/7qPWZRAYS3GNGJVRl8nJRKr70b50YkzxqK
N8RsMBm6o+iaGHOZ6mJ2SMm77IxmJ4kgLG5lNTEwc0472OetxbZzCAXRSHo5k0p0LEFIcuJua4R/
3kuHBHWCFCUiUS21R7AJbznm3e1wK1sJizSzmNhmoqyvPgHz4ZmSV5tY+ZWF4ricpcEE6pR0vlb+
c+PSNAczl6vB87pho1VSD6aYHXsSOw0PWI3yH363tVN+65+uFtpPqYu3CRgmH9yPXycD/2fsLGHN
KncPztZBJszg9/8RQ8CjSPzksgZyzUn0oDwtyjr2Ec4RfCutMIL3KJeUWxQnFxZ+gtyugZgz93I+
wp8BTI7SifolCkpIKjcSkXnVBrQm/wyVatB/UgBDHfvWSeA5lsHAmoSvMddNYPt8bKeQ0ez1wcqA
F2IYgJfeSeRfAX241I7b6GFR2NkRfdU6sJKp07ealxsGCaO4KZDbXQUfr9vBC2b6sNA8jGXybSId
Vl/3/WmnT8BSJKYailF2EJfW+WrFbzD+AprB5j64HM7kYcNENl8J6Ba1YxtEbHjSBtUsKLkdeq09
J5WQlwQYrkGfdZWG4W86VvkA382VGoQdkjFkxRpp8Kui1CXwdGiaqJ14OUB5tkOYWFkWpYb9kvw1
m0BdnV70JNU4AH1Zsi+LEsSd2yLniFCtHQpFyj37bRZskg6zJozUGMDgfWwS1v8BSZIb8gOxLfjK
c6Hj0NtTRhTfSiWsAcw6OUwdQrSuQjBHiNhnNaOH8hXrXjbY30yyiFxuFbXrgoiDUtgags2DnF1R
TlIBkvKP3bDWXFLPHvWr0EwqX7ZpYNJmaVB1s8HutTzf7YLCKyzYFO9TSQRW4E4eFpNq8h/khOxG
NJweR/ETA14zzqzwx2HNs0s6dCU89yqri2ufA5T3wO4Xas0Khb4zrtxZzjfU2RTwlTKgG21T6tEq
sGbgZgbQLdGnkZnxicCnJu9PHwL7tzw/1gLEKLoAxtFSYlFHB8dzcrIkeN0Cs/RtgWdU/oy6OSa+
srImDRYCOUDwwo+2pEXxltLEAZszEIhH22GIwSQLv+hUJklOzj9Vy/8TJ64/+0hwk7u3bjvG+PEM
67ltUv8gKA3wH2pvtZAmoIXtLGjEcvJrJ4/nSPqjKfNw6JpQbhK2NK1i9jM2eVRa0mUCZ0upXYqc
6G2yJnYWFOGLY2JQdp1ESF7ZPF1jb1PNDuz3HPX5fnVmIBD/4v5B/woX7tkllYQXnJc6RLdItYTM
+MSqTDTKKKrsiQaDBSUisg7o02cDJ7wyRwLXYfMoF6Ct/MtAXPcUndYQuYgAbhKMW58HgRtmJgOo
/pxGgK4DL0YoOUOyHGYNUffAl8/RT5fAfQgIYJYfbE4CClq9cL82XuOcIeTJuIMX5dykH7K4253o
r7oxvEQPW1m6tvRam17YZMq34Q5ZRCoZgje5Kwkaxzl49PFXvz3+fsjQNLOxTcyFteoSce3pBDlE
mOoO60IvLkX1LRQsp7Ywcb+sHPz4lMUPbVoZo0So5u2EWm34wDU3vLvT73r1rPSFFIWspsLmPkNk
g0KtWDmSCmAOrVb9WdiFpOkUac5rmBSMcb8N9BbDXGqk1NBwBJBWzVE8KM+6dNs8VypCHWUg50x/
VDefnYWY6uaTbof9p0RrkXssT4uP6hZhsaLdk40gmS9Ra0kfhWirN+jqKq68itZAkQ+lE4Uve8kK
o7Esv/6vhMoANtk13Ak0ebzvC4AcwNTZB/eMyHldNlVHSHPCn2E127u3PeZ2fE2DlvKxI9mxXZt4
9xNe1Lu2iuFbVpDu0EOBS4c47GMlKiBPjSJMcKlTdN+b1CLZviswzTZJCeIC+rvNSdP2pslZxzk9
HrJrb8ZLOEt0rSa8v+Oacwwup0HqnIKPYsMCcnzEmjoNjJVaTFJ3shmgrN3EYEbGlCyQlbAOR4l/
c71ijOBxFA5FZHBWo2JS+nHngQd21sdnYQJTNv6/x7vMoKFdvoXP31Mb0+TpigqYkO2JJnLPwTwf
BbaFvOf5ZN7Eu4fqpTIVHLAeoZbM7Habrt8piLsr5+JL7PjUN+ZWd3JOlrGNcD0smS4C8A+jXMcB
G161U1+GTSFS/mEbzrg9f90ghSpfwvZSsV/MKvlOFh3dOKs/qTSe/lh1ell01qh/6IyBLw7Rgd+k
610h00D5ZhnuHGltgF5ls83c+y7zoSVCyyyO+D1MUoJ51kuPumQIOravjHptZsH3fc/FcMRConVB
+Jh5IpfZLw9GgpnPJlX+KK8i/yxrRD4HLlzVRId2hsS90F4uHdjBPfjOtI+FJdYWssxpGIBKjRwj
cG7VslpQXx7OJMSgckDijhVJ0RxtvZY/m6S2QcqcMV6ZWoCs0bID0wrFdJ5mN7o3Uqhviz/2BxWz
4QCN2F5F/SWgUWSaMtrCcRPPAKVbqLfl5o5mPQ10m/AK0u9lul6CAys2Ewn4Iw7AcQlJv5f9CJmu
5NPUYYsRNDDU2GuAa5ig0+XEW0tp1P/soliNJ0/fn3/PSo47lstvtxGLrRB/8cjFZih9cdJ0lXjF
V0GGSOkBrqNuCnTKsbcndGux6cmIj9h43d2gAoeC7a3fNEKq92RSVPHl+AbbBIA/6wILkBqBaMBk
oY9tSlga2b82yR6sEdLkiUI/su5k6UGevQa53Fvcw9m0nP5DpX1JR9/h02IzGIryPi9l9tnjjZ1Z
pUvaKY3t4QfL2kNV25XkO8ohG91xF2HWnnWg3LlsmMfHHWq70HeSyh2qtsY1GwsseNktHp6Fjvn9
Z3CSwPzhkHc8q/mr1BYnoMziwyQhk7He7tuBa5OTkvkc0XytxgLARCZVRZ3ldbta9T5lTRjmQNQk
OQf7PjOO+eTFqMeTSamuKZDidpUjcqASOooFSePub94uqyFYsw4V9y56w7hWE1VtsO+319ZNFtgj
PoPT106KfAv0kikIgwTxlVN7qWAnpRqJeBZgrg2PFPHXNO/j2DK6fSwmQgfXQpqoxPvh58pdhp83
Nf2+tYvvY5ZpRomvbBsafPCu1WnsbDTxvNh/6hHARySmrWdNDCN4fvGPISImfjcr1xjyz7DAPx3M
ad2VNaV2muEsKZuyeQVBTNslAvGuGaXXuH9+F20qyxLd8mTpGfOjsmo5t5ZWlbIftAAFdF8DEqej
1tj0PlxZ/B10/gwZ42rYIsOHeK0babBc6XKgHFLoYYzZQeNIU087jivfyydQAs2opGbd5Wi3hKYt
a1D1QhSBeYgi/wpJ4wdHUy2xnIm8xX9I/qGfuO6U9pw2mHwqof4vnvaet9HL0Y79ZwhpGEb4onN5
RWc3IB4W5mG2sMzrAqKGvMEI6C3Rh5V9C9xK9blqxjTDsPlLnvSLAZMVvwLvukYMSRe8hJiOwHRD
nRjGEqsGezfM1t+g72HMgbI4yTP38htur/tjd3yaFa7MRfym7YlRoGwg/jH9nQAh844L861aPiBb
+eolRLuK+mx6H7OFNrK/aTYJDDRFJsw2PD/vPhAVBHYAmHj14iRPHGjQljA10IDu5OCtHmrtYYFs
grp0O1J1/OJxFbet82DPTiq/he5bkFOmTtzUhkyywNKWy2pupzu8GSB5GH/pGM9KmA1YJ5yQ/lYO
lm6Q3vqp2iiAwdSuAIugz8lkzAzwjBLNXd9e99JdPwzTFBeqyztWnR6hTumbJmPgAxoia8se8fZt
2ar3YXMf+ZgUYuX2E239Hoo3eV4EN4AIve4SKacFTF4YjofwG8ruHr2qeAFTfWFRriS4WKIwdbYQ
XYj5xRqYHriSt2o2Xg320Leb+zmyZKfQGnirx7+CFoggalGAeIILM6kB379EPBZR+JodKb85Ew9c
AJsyeeAxZpTzAOGqSjnxCxJ69tPfkLKawVKDLt2h8804anY8p4mO8Ie3G5MSF0m+wqra3gfZwHVp
lauQBuKYoIruCWkmzhmzduduptj0hOeljyZRz2ajmfRHDJvkux3jkW/WiCJ7lKyUufCRxOPseGgD
5WOqgtOyeTU+YzRSHF63pSAR/iDLx99yV5+vA7fKQYIH08jqKoBEhx0sIfZjUF56/YWFoztkd1sT
AUp1QMDX9d0W0p+/7g677X7ZQFYhzddq7QNgGq32XJYNatkrKwhN/WgsK22tdQCDoMBaYlD9JlE8
jjPzXvFxEZVys8+DgQbRcxGzRIZAFaYAw4dIMI5q5SgDcb0bJBiAVg6xO66mUSyMwCBjBjrlH6UA
QWiYFwqSO0g6xyrKoW4S31sbxOV0XwKeQbgsSmT1Y+qkDvzVSN7Rbh72FcnYO69ohaNG/OJVu+C4
AyT4WP31OA3HFzBLRxhpjMtg6CBleh8b9nxQGEpcAiDkhfDReniflXU48BCher2s5LD7D74qRItu
BD7AexHKnQZOR13DR4dhsAO00v9CFepXf91kSp1ZQcFKVOULo+H90NOtnI+S5x3PFiT6ihbhK4Fx
YjW9J4/WSrwELzw8tHTfg0bsj652afA8vU+T72rM9VUdwG8tveBvUdr7P6n8oyvWQbQyFIvSUWlA
bgMzV09mnCOeapJudjd9XacbinhEhQo9rWqNUqz2zMMD0QO3DtBZC2s3GdGrMKZDuBhAKOHBuSLI
Xox6VAZh3JsabN0NjfmhUFBqBZk4zibvSWQU1riBTBDbexQoqVnpJ3W2aFANycLftxeumodfqI+0
kzJPwqjcbpK5CRWk43R234gWtFNDzR7PidbtNcs3Dga17hpHg7Tjf6nAiC4ZrQqZaj8RnqziNpWg
RJBZ7oJEFVYxeZlceuV/6nj6kQiBc8ADKln4gA24Aco4J8ZK4fzVMt5dfkgr7HCDe8sD1jxcAB47
x/Pt7NXXIQZ4WQbtL2/+8MvNvR2qk+1+vYCYYW++Bh+kZxRTcKezADWEsYUOIEVNNARxUuPrheOp
s8OZwUgtfOF5z7Zu7xT70mwTwhCAIUrBUJK7bP4MSXzJ2QAKrYk4IWPuSaWTUbBspWz7RE8RHn26
oWPb6cvNl3u8FUx6sG00cS0qeP8eb22qsKVQ+sNQOlLvxSkKfuSahcVr2vwLHlZDQt50AFNyOr/x
4W1aHLpVVJb4voTVI6p6eRWA3GrY4+VWqaPmWj6DzOr/f7XO/BDlKXKsQzvgnmL7XVXzQrEKdzyr
6xbdkTvKziGCgGo8WUfhq20PA2BsSKmIaHK2vncyDVy8a/nQkYAq9VA4d9LPyXEWtCPm0SJwikxV
wAakeC88ufW7XPZVVK5ei8UgyY+UUTDQrJcTS99UFiaOYj+Sajx1FHcJIn4HrE80/l/2aC6pTjeu
X+XzhM4G9ysy5MhEsVZ//EXAUubhFXSqQCck9W9PeadX8eq31JpV4AJi+Jdnstv4Wvxi9I2Bwzdp
QeOyFqW3S+r3817sO5IA3U1a1bMFT6JQi9pkrTh+WascISNqroXeNzHwE2n7D3hyNXDjL1IyFT3e
X4fRI6LO/JKiKFnyenxHBBY9BhcNzp4ngFaVpb01BAmifTGGRkT08vF14T1rscKWeU6qIJhFI12B
nT7TjYvFew6gqlcHwnve9by6EOES7rDj8xzdz5F8Sm46tkNsSaWRwXNrhkhC7IzIM3Ty2kjkB8pq
ksdw6B+qc22PPx69FhpTdZKZdboOlZrBSUSRU59GQ1JCmDCzBcRK/y+7R4KVP4Lj6EKnCBP646zS
WMCQJP/Qem0npYARTq//8U2TLnxo9c2JTlf8dXtq30Tb2FOLeY5SWhazABDQ6vyrIj0DWvJNE9iS
SKslIci4J1hslVK3atECVIlM7HTrmQiZM2JIpYIA82WKLA1IWPxvIlZXXh7QpsHS1SM+/wGU72F9
5j+6uKyU8CQkBJhhs+m+xnE8KPJdRDTlwsVoW8y6f7pjltKwERLSNXRVmILzY9vH1edtAjaTyrbf
j6HUYvyaql/7FtqQ0y64SQXDOgIhuCSfZ3nBpymNIcPMfA7g8r8MrMXhm6tMTMou05w+XZ6zgyHc
Eok0aNNqn3ugb0xSEWn5VpPZbIBDDX7gtcJIzoX1yh1wC9b6rwSbXYdDpBMCNqOp9cboRkUq7FWO
7FdeLxSFyTbVAOOz3vF8r2z2trCiArfDd6TJL5hQRqPcCoOHZUHyzRIaQr2XuikkTOkKF5I8hs5L
iT4bRIlysgD/3EM0UkabMKd+5oR0XZNSSams5UhOtkFlI8rGEPyLwc+qXf63wMi4R0UWkwxnPHgY
J5Bal+0QKUpFW7py0pD5ia0/YpD8fkrxaroxhZ6CV8/DyOGbbcGq+BWexgCJdErRM0ncNpjA8MeE
45jvsjy0m9uPJmySnx5V3ctchUcsHFYbVBu6BMGdKwBycBdkhdomz4bkfsUVxTVvJikkX2ah7wdt
suCRky9/w3rwb1yjRqTHJPF8NJQryxKjx1wSv99dseHPvjVmKusP7n+eYVNEbdiW2BqxWkOuQ1cM
OzeOGu02aRHeLZEyR6lo0GQLNwVNF90nqmQ09bdsshSBgcG2BnukQBsOlDGdn6s/9INEazhhzWX7
Jx/ZIg5Se2z+HdCOpAMzh9MXJirKbPTQHsnRfmlzKXezSOOROHhyrfKC/CpMGA6CBh3rGq7AvtQy
TsNCqUJmZeUAbrWAxAZ/fR9Sh5P0uDgyvfIobftZl9g12BNSYwqaaAUR/fniiZ8udIi92+5UTtwe
CW6hkGm3sblS0vTvQhS1SD3ml3/DEaWxh3/prQ7RE9YcPPkWDdFWMe+025OLp87Wl0l3uYgKcBlX
BzJHJCHrYVCPZag9ClAtk3iacnxCSKQgDYhJjl3JHFSI7BhIv8I/2vmKQCx7eGn79qlyFMUlnPFh
NbEpIvfSXihY0TVVGlqIwnD/TtUAlQDeJeGEijfUKoJSnxrEjF9F4CpgUQ/RhCM96SjL4DoFO5FZ
KttIfbSBYfqXMO06jgKYgQ07k2WKCZvH4kwncXLEMq69azvtX8RumQpkqhXafCBjC0F4mTWvrJrM
LqZLS1Lt/y1Weu2FG/8WjZqfU9CrayyMny3MRUDIh4twmeBM2jPD0RbxHT6pfFtLGtYc/+3Onuux
2mnKztbEWlwm1P0YN/F1emrkSPSE215r0fIo1HUsmCVKYFwt95aHS5yfZ5bhuOpBZqUDBy1GJ5PV
8m2w7VlykA4eFtgp0aiMd70g3z8lPm8l932wNXk4HsXFc/51/oontOBVAC9saYBfm3g86e2HCpGJ
E846VzzE6fvmPgKS1kc2PONAwWgfXanp4E48HiHF3sv2TvalA0ypmaQs26Cp/VwRYqNBEyWwCIbP
BGDGWTj6Pl0AbyQRTWQNGqwquzemGKHy4969i6zNJTwvOH7jWt9Ia1Pcy7G7eAD8K3ai++ZIlLqg
d6Jgi9DQZ7gdRG1Q51RpLJrY2rBxYFscNcYuXdUwcb+8LQPKbitZJTZrLcppn/D9Kvm11x3wg8NG
TCo7ApI+6ijfKy97QbZLkxcjwj019ZWw1QJxX/79Zs3f7lEnobIWAzUQVHxvfhJNCf++NbMIaZ3m
ABPoM70+OAhcZkG3afmoCrj5i6+APrdYQo/wWjfxejiUgQvqmCSYXMA/IkD544WaXExwEhHWBcrI
WHb4GRAePn8+4nn+Qhpg2CAOhAxSdMWXGzVjauxOaVi02MhbvOVW/xta5+psnWcn3rpkRToKPaw+
jRKpOJzOQboHLUp/ErpdT29CIKz23m9La2Wi6dVkJZyruOa/dMblF6jl1huCvE8Ww6HXthFrOQ2V
+nbdJgx7xRyA0OH0Nw9k+tO960U691KE7bOZrkIs5GpG8iAUiZ9iWghXls6KEW1n2X1BnA1XSO1N
GqM8f1eQt3/x94prM2ivYFalbIfuhPcKEelK2A+JVfH9d35aKrGwPexI17vsHvOMynPP7u/zI+Ba
nfS0WURCbjud5QLYLwnNCbAq0A4SOSVrVhjIDx1bc8p1A60LXreCIjDCXi9F2TSzNNa/Pe9QzJrx
oDjAt6cTKqHMVt3lvYQaulJKrhwxQ2LfBvyQYnEFFSZpSCc//F2quAM8m9/yiYVIDne1396QyX/H
0pMajWIf65znoELcRK/jMxgjXLcNiHQ3KrIluHasv2rLAc/zffqbab5NRTermt8tAeVKtgL4VOQn
8mzMPiP4+kS6uNH7buG5bdsqqteZacje7zbo9ymOSq6ubzDu306fet9WYBofTck/d6KCO9MbKoKD
BVfpnRIeOH2kkQsHpeB+EAOE8PdRPTUBVfyVfPI45OEy33qKUQGp5d4D/xrUqRK2P3E9jr1giNhc
x3QVel6swJo+LlQFQJSWhK4T4Ggf/0jmnjU+uKgTUwa/3KGf7qgc+q3tLFBUMa23PtPQGP6yjlvg
CJJnP6lVnmQ+vUgSMvsGY05fNMCcaCS7T28dpaWoGosCPj92nN7ftty0vOy6HeDoP4p2tYMN9/ac
Hr/DX4QrkkrSFmpfkWixnBLs9aZka2Tst6HruI444gd+auzc20mS4+W8q2nB7KVeVKWowqeH3nxX
fW9ADAIYK/eBaMxbiA0d1hp00UzRHEa0Er76rg8J0J/o4FO4LHa1LmH2KWvf7JBEGvRuBRExF4nD
YKtRFKGx5hL2RAbWW8YXiCdPBRJhin7DlLrw1nSuozMWd/zMAygv7VJP8YWKPersQDny7evTQ0V0
AZ03Ywg0Qz8Q109bhijBt5r02DQaz3ZwCPcKIO112z2tm2rFpZ5ym3Vs7/meKNJkQw0KI1GRVhph
chLQujhp0a77HUqh7AJy1DrEVn1bUJbRvfk9KOs5IN6SZbSPLXAqHDIqXY0Lxrqed47YaXBqOvPG
cPRtRhsD+JWqHJxShZntuc/d539H2t5ml7BJsh+R3CsG2aF805PC/5+QzFnxJdsANjd35H4J2yqQ
QxxnVToxcJKuf+i4ckbK37nRJrqSMLRzvVkws+OuYjDjtFZoaSu8ZEpCVxOTtpo4PwAzAeYABty5
ACpSa3KJamNLrchtUwlwkPCzwX6ixBF7NqJ+/ou1+8B5/KU28lyeAUTAWR0PdBLerR4Z1pDIg0jn
En1MCzAMnIbobADcJEWa14IvkGwR99S0of9BkhLjxvzB8XLZxbWXn9I+gA9/uORWG66uSFTDBRI1
TDEQyf7amF/Ssf+u6+0uZ8mS78inFvV82oBUBzxJ+9cevnst3RLw1zAvQ/OY8mpcj4Mcd9iG2DIF
guU7zsPuzJ8MdLSUYxdPYJBOFvqGYTFZXAggMwzWTNCYb0NJ2s7psfHccS4T4SkknNZ1Vpg7xSaA
6CnwM6p/+8DuOqkedlno0o9NXSG2wy6DKAbk4Z+tSe5Cm0ZpXtGqYkFGF9Zsps+a/muxxHoTx/PA
KQW+8vxX4xUp2AR/HkUcGQ9pe7kpafNxVgI6+46MXaXF51zo8igZ6tjIyOPI3wc2dzzxmLEtWTyB
diRQQe9DbaXPY5Xt+pO5xd10cCAfuNcSBOX1Z6c+OFTrcSGSfphe3Hg2X/FsNWF45LitRI3tYunW
ByMaeD9ezPTj9ukdhc+mSWcla/XCI3iwzQyZokyAog0cqSrBXvIa4TGHSwFq0vWyB5SfQFrwJZ+d
L8e0NPoUVK4caQ92YbEgf4MiZdXeJI/sgOfVRRo53fu2HeILcVKeWaM8W2W6wfEuenxpQWiEO06x
jUJBsVyhRFpyuFBUKAj61L+rzlNX3/KpgqlMwefluVP9EBuYYBPdPNaVdjRYO081rBtyH9/AlRpo
2ywwFKSOp68gLJim8jvv2PiARoK9D5K2XvZKFAwk3aciAEs5qYHzWSqw2HBoZ/TutCHsAE9NwA7x
KKxhNTSQS60JWYwwWkTU2LLc/5vaVMzTZ5YHJH7xrTRzRzRJKyk7y3aL7WqTDGLvl4/1UYYRzslm
Bbb+/3gG8PUK32xUvLOyhDT8PGb5c4Iwi3zo71oIMH88/eJZmLtmHVm9nf/KVOsIabIOhq2bEs9c
2fcOAsFnB5dJoUjzzNKTCC873kEnniKi+BpUlKGR2tYvYrPSTDVae0uuHUOFicce+oyTsPnVlE10
hE15GLEWuWTYQbfaZtRbkc0p38vezTLvjHfiuOlsJpCay8LLjQZVy/VgOyTU17kvZVf4H6ZjYtLK
S/UbtdC/Vc5YPT1P6Vg6McTygcehom6bWo2YXELLZXzS9Ro0iGrlpjtdn20Rrl8kByOffDlf/suM
deLEHJfD+3KLOSSwVAjUsXI7O4e0rxnmcn4EtWQn6Mb3dNc0M8d/8ZGoU1OuFt2EddgwC+Sb64iO
PvWlVEYwcCh8SAUN/I7bK5ITE7d83GLcchOrvRdQjojqN8Omnx8IwgFqCQMZHwx6eCBrbyIIQxG1
DMAlnweDC6c9GRN8/pJ7ki3fwX7KX+V/C86XqKsSbz/GkRK6bhSjSRDlu0gC4NONSqgeQpv4zUtq
1X8bNBKlNXRDSi1n5Q1VnL3XIZwsPFLnrAdb5JgPHr8NaTdKG2Obqteh2A/d3NQ9Og+DvvABCPGm
epsV4xlzRABb9w1OyMmBqX32nrOGKX2V+42nNONixJaAxWsuR0W3aNk0+rDWXWb4Bvi26kU4HLQK
hEgAc9FbHIGP1WTzzAmlDm1i17KkggUt4tsTJ5KnhuI+3nttSdhrCLVKHwG7PKeEnMcaW4pNAciA
O7JCqmVVa7j2hCmxml5/pga+pJToPFG8di7gWSV3qlRBil2NDFhUYzMFmAHRxuGrTYH2u11sDXMe
wVb1JH5tS0+3oc/huySTHgU3zB1oXcn8Sf1ls3Gfcpb9E4SrI9fapy5vqgXOG1q9iGDxfOyfXDWJ
pfPgrxepVPB+QLpQxh7i4a45Ee/0opLeOKiRjsT42yNThaZyNdAWcfQnUlFRkfRS7JOSe7uhRf2R
Z9yXAlK887IS0647FVDURJ1g2AFYxbThHjiP8CoRNsl9BtqhuJ508ASCyFoaVSeqn+U1RXW+WRz7
Q0Xt70ODP5sfjZMl9G9HHd8pcmCw0OdfoO6LZ3faDxEGy1wZuFGdmmzoNBftuzacFliwEytDi3kQ
CshJai2EARfqANztJuPdZBZcVUo+4t2T7w4tNuslilalSm9G58eaDJfRRb5vulM4krBKemwG6Os1
rRw5ZF/t0Pydgs4hW2omtxhkyyCaaZtsX3OmcwtkX9K1ARLLJVi0LS91i8ygcaYsqQxcAHDHx0pu
idOh3onoGTdgU9RbDOewaUyUSE7a66OQQGEPHhnavGa4jYt/idzeWXnth6McHaiklFbwgjRuY32L
GXu/6lSCX7PraBKrHt3dr9IAc7bKSCkkg8WmDKVKi+WPtioSF9hRSN5VyvKs318x1Pzu5Eo/8txz
XTlPVNdKZtpQOrYM4mgHTg5sig880FJhyQPWyuBZK71lj20fP1ehqB7NsM+paUGgRRGbblnfY10X
7tq1MgAE8hEUmgCUgcy142TexecVEmqKGAq4BGCPAzn7y52V+xJ+2AkGSsqF7V8VTNLOnIn3fjvI
u4KsXVATjdyYfRAxFPM5pMYFR6sjLVXbbNbug2YSeOFIHQvVI9lAOq42I8/Xyy5AM4VPTfl7jpOS
uFeLcd7pYSM19iu5xrCYY8k6FSkWDuxcPiERQVMcH8U8080fTcqy5L8QiHFArupll2K9eG/sh5/m
Nj6oOKlDp+t8EK2GtGu6f6mY/uthD3iWn2xW/sQGzSnbLA9Zld7Ak/2Xfib5Tp0yykRmFnfcppwo
dVAobGgPHNFY4Fe9wbAE86K3gYrwJd4Zp7/Ir9UHUNVatVX9kBrCYr7oi7pBeHprnqk0O7nBVLWF
wyirJIOvAMVC3rbUBJ81jp3MUysF3+ypS8FAJfAS5hBRCDY6SANhQWV2K1+XN+FDMsjGv0T68OUC
Zqv8nG1HA0kjOU15LCoCmEwrchALftRdcBl9ZPqT75pcuAI6uLKU1irseWObYRmA+/+wXE/MoiOK
irmXRm2sU7nz60UaSS/iblhtWYHlUZXNNSSo5DKTxHR6vPeJUacbBC2QpuL4nxf+Yb5l6HC84QwI
VuegTdrCHYzsXVFCiDS4MFpYjjvXmQrX+PSHtUzswjgp7K08enKNdqpQ+Zq1s781uZkUQy/1C+tg
pnyqiO2sZaDKZwQ1kDB0gZslOXqubNyf43/plGrVP615p/qk6eqogYB7pCQkbOOL0ZVQYbm4VNXx
eXHjfZVKmHxbC22CMSiylOwhcQ24ZOlSmB2lEbBJJEjJnw5YFlUdcXeiSxgmc0j+F5MnUrUqbX0G
Y2n5Ad8HkAf289x6VyJAT6fsOFAo3hCdK8yvsiKrXC1+2qothcdoe2wEz8e5vZIgsjULBf/ibaMi
BaCxpm89lcCCSkW27xiZq8WiFoIfi6lGNla6DQsd9tnWp6gKIg0YPrJ4J2L5/4HOrZCZaJrK5/mv
Zu3iHD0v82kMH+0UFvJwpHOOV8FCVAjDlWECkVunEjem3S26vm/DoBE9YPz9XV6YZuSL/2nnKjxU
y88WLbtfTPMnjMFxTl87VNPKqWXn+Nuu8XS8MM2i5p/epwNdC/VZA+4lwoeuf9ZqW5WwPoHhi5h1
v5Vr81XL2qoKtAkZC7AcQPDp+yHqm317HXZYhk9xLTL7PLqYffG2ch7xGmUk292CO/rt1VWkLVIs
3oI1u6Wo10jH62uKH/8nXOUAgUIUSo7zlOyPRmItISxGMDRtMG17SDxKEZL9suWdG+qLY7DvFPIG
XaxIJ3dgHGOescxEqKVIGvxJNQr/w+umJe8NIuobfbh4j0bB39f4jOcRgLCYV1zYldB1OZ7hhStU
t4GPU8UJcYxZmqMzhyduSF4W6geC1FKnE/dZhwz3M7FCiLgHdJS4SPGt2IPbuzlbvvbONbwboyY9
ekvFSi+0BkLdfSCnPhZ37fJsV3tqOQcoBC9YAvQfH1C4oS5m4eBfpN4gdnArKC2eFnmlyVIf1nES
tvC22FoSy9xE26AsYXZt0IAXVpksg4YRgLyg9NX936Dy8UugcL4RYAClDlyuGmlMAvn6Z2tiUixm
t6UHcHk6yqDEHmDL9F/CuoF/gX8ysuCqQfrXpmvTwuruh44savMHNDuZHlXbaQj6Ry7ORW+ru78N
E37Sdx9qfYM85S864Cx1/TcDAtg6As8Q6LQHkcSD73ljeBeyWbHVs71EnDMgkt1jpnhnYMOIoYF2
8jI1A0Sg+4Mmcyu5yZfPWJt0Lrui3dAkoS2N1781nZsvGZDVJE5YeRKRmSkpz+Lpls7Q0TAzBNjG
RX1stAE+cv2cWzeqAYh3e4oHCtXQPPo8VYr7btiBD2h2fE4OhzCUANRJ/s5ix5srS2RiHnDfIk0L
it81hMQMglv+K4HquRv5m9mXl/Y59RgVlAJBnTak8l3wW/lolkTtI/BaOsixEWAYOq0Vlywq3+pd
B5ywIlTp+icvAbmtU9zoCI9UcqH53l0RF0ynx2frjWcf1XcvFXbxUFeq3yzY86nvZ19NZ4yAYS/1
78mICm6ebHAztH1dDuW14gAUP701sqJY+Df8ReQpIrlCZmxTDrRhH3ZqgC9Gxka0bl7UcRHwf08V
DGP4TSu+4FPgKQdd4+bxrIPeycwr1j1LE9tHaaOCetPnd08LA4znh4GeBBGuLUZjvj0nlUS9W6cj
HYeZTGolf4yy274Y9eGydLRso+c67oyND9b22lDVy13eomxCjZQ7JSdLvywwqN5QkcOxsuHqD2IU
prMZlbXUR5SG+Dcb+VEDlmdH89M1QCxuD7VUyhAD4WqeMBEryLgHTe82vrmQMC5aNDn7JYpMQREL
/K3n5+nH0uC1HZbVgCc/d68f4mlnJGU7DIIA/4VnWjBt3jHbX35qp3tlIZOMme9062poQkUlP0jX
TpuFTPeLdwLKcb1C99aifpGQF4dVcoSaxWkiwmZix1u6zIrCeboz6PXr7mI6E62v3YSEajYTg7Tr
SoNbpAP2rKTACmFbZ70hmN/Aez1ZtiOwLzBAPE7T2aHdu6QwNNlVVkEwEf6+VDvwMHfR17znagmY
KHCGqcC7+agYI//49yGyzsouwEvD8eu5nythuF4o1gW5l33LIy0QSledsKJYn/SOzr5uhZA5TpsV
Qh14tGJlufImzqlE6PMzqKGZ22SapCdtBPLrbxMuXDTqOBV84UnwMdTJF+smtQuOmq97/RKcTUW0
4dzXYwt6zQpf9Ys3i7s0A2hr5qJsnzbwYAfip2BWO4Ul3oREEh1CD1DtgdIbZtEucLZKwqCJJUeb
ejt1Ru9LODz6BAAVJeMA+ZSdlHOPgP1HyqpaJXv3Uu4WirhMLTzwldOQUtC7nJ9n5ZA6jm26Qxci
rllMaJJudoIlAsMDJW99R07M+4OnoEpeAw/KFf0m9uTRtJ6NdrtNT9BXouQ+O22tX6IfMs3rH8NA
imcUptiW2z3EPOJ11umDoi6Rz0vah7WXofRpaLqKuAP1224QJ3WtuF3121jNT0bG9v3FKUrlzVG9
EQGE1Rn4Xgw1MIqprLldpmZzr3SAqqSgLATnLSxHfVjwWxL6yfGTj81AXYwR60tJJRGYEWZoPzNE
2kXbZ8h/OeEgBNbWMf6wc0Wqs0owc9/sV2E6GsJFLO6zFIclChKFiBHDRf4S74gmaXDk9UL4/sIH
XMtwLZhq7AKVyN+ICK2aXymkV7unwWkSjSqHWowYhXAaXX6og5nDJMJfF0rxxJrCzVoCwyeuBUp5
M0LvRw2/00IaAJ+laEayeqmMr8K0jNCyCwMxskDHyUZya3iy59LF/8ejNzAkWiO2rGUVPfg7+kOW
qPyS1iMmVxRAWQJvXEqMwir75N8EQiOvEASl/Wks/I14Q0PI15p9khSoxsGgVQchAPHn9ZK3NUd/
CdSDOQrJC33EVkQLIXANOs+pweVotaDinAbhZg++2tA0VItFac0vD2VmRIfapvWFx0grK1FF9rku
yqPEOr+vjU66KCnKzGkF7pgmSPtXXLDC2sGvGCymvtyyqB4Fg2L08peeb1qlbDgFxA3IV7QeuLIe
3X1Em4zlghscG32qINVj36EPXECWGA31PnAnURcyDqSIFCevRu9anZCc8T1N2bSKCQFCQDEAQim4
xGNMZ2VJkPJT/v8Hg22UoWiMg0dWI61pIzVPo5zXbo+Q3Dm/AVegEP3ahiygt9IbImU8acEJd94a
QPJ5BlonhZoYZUDF5VFaH7uK4+Cg9gqFqW8vHmDSMBMoysT6KjLTNaWZHXHsIVnAMpTTt2yhW07m
0MNgYCoGDnizSi/kRVN2QQXuVCBaZ68JalGdapdF2u1EIyVTlrjGCle6UUUr5232tLZhJEnzx34e
pex26R5gmjMk/5cbDdieJ8jHvb65gXYIsfZ5+1ukdyQQcTsfrcz9CB0omk+Xg0QYnsU0uU5iPaea
fI4AjDuxnQjQNvHg5RChiWhdwTe7PUPG6wvQ66TitpuNO28YhELhicTLfhoMP5/UczIVwxx2xDl5
5I83EdR6w6+25z0RXEZEXwQ5WPSViJGqy0FPDC7KhrXtaBBNUQb7BBZKM6tolRGQsSiaU3t/bYLx
KWQdDjEY9iMxxRg5BoB8p/i+IS9/GyAbbp7iUZKhFVvENAmiePM0euNUbV4SYHGh+rdyxaHAYhYo
zq9yuSpTnW44JrWH2GfGtvs6SV9qoo5Udi9erg95zUT5FXp4XXelwOYVqEtaLjK/M6OlqYFm2CxI
WDXXZzoM4/wmACV/T3KMPrz6Za4mU8wzE1sBZ+Y2pquUezB4fOXnznyUxCe+5elpCR8FvdLPRe9C
Sc358E8BwYyiL+fZR9CpXxrBF5p9+BAgyp6RZ8gzM1Uttl2qNfQwBWTrJDOSLsHYlT6KeUSGrAv5
QfMElP5RQod31VUpzNqmRTJuXoIF7lNDSew3hpgI0J5vF/c2wZUZ5CuDeCo9dJkr2BgHa0kJ6dJm
J3cy5pIiczH5eQMqp+u5PrAqtPN8amETIweiAWqeL3fJzkaj+dIumLLp7kDcleK9PmPoJ6d7DaKZ
bZkAJG8B76wKPaX7X2rJqrKMY8W4nN7ZkptPuhbnduH06SJGwL7vZp5v///a4+A0LojtDu4/eArL
bdSX/qxFFWXAw0vlWTgTNgwdFm7JNgx/i4GpnymI7Tsxro7FUy5oMfvCyOMUXt/4wmUi+3RQ2Y1c
/9jD6A6gTvEhKKqUCCEsINH68744lYw2eKvy9ONn8J+tyBHiI4gJqQR7VZVXrhuHwrJ1G37dG0AX
s9Jamx+wv2arpVrEZmlSfA20fKU+UOtluq7cAep5mxBxWVuQzpBXsCMbHWxLpNSN6BHr8emCpMg4
9Y8x5zLxtHLHhM/NtVZBHIsfUN0JUhHkOnUFM7SrYPFAfEIO28XlAsP5g28OVlk9nOAwdChbWfSm
u8rohOtapOzv2tCzWWWCrByY8FrAPcNt0x1Q2F/g+RM7yh2EOY3Tozocs7wRDWdcwG307WTeDdre
SfXU40m4+4Wq6NNCcvIfoKdR3IsNR1lbEtcDsOkPieBPC9vXBsdYvSAeengpmBRufgTkHq3Wj2sA
Rg0h9LQysHMCnhqIjCJVA+k373xHkowXTBeLha7WOhPR8RKQjduFH6B68MyLm21DflYb0GVR1gMz
ufkDsP1ehUTN+KD8d96aRTcJzTplXqYv33ZNpo61CdM9zgr3Le3CY5uvW2iwFrQpdVc2iOCoPt7l
0tWycmwA5m5tS+pmtLnwtktE48/kia3FYVaYQ7syc95F5FVFmKEPXlM8u6yOyIG2Q9O75MoaRJ2x
POIXnScz2jRV1fHI+puFZYzmcWw9Jdw61UL5KQucSbtevSx/tC4WW4Lh6NNnfM4WXTG/T9y2eqga
XaidAvLzsgle+59NL+4xbv5r4zLPOwX6N+5+LerxVIWUvXApjYexzrTA/OdaHiXaM1Or7YTAc9vA
pOpUA+dm1SvDPjY/+znVEO979sF/LFcNNZeLQ2GcrUnjfeUxNRx42sclXfoISjT23FbG0phOvZCY
YaynRF2Gyc9mF8u+ZHgSyINTnXr4DeiOp/2tikAqvY3GtLhGQSLyLVPBXu5pr/e6qyKQh3abPVsT
4N5UeJ3MfdixmPtElUFi9EX3hGkWZMQTM2Vx4du+0PfM+munE6CP+Ilp80NNyBg5v8mundaY2GUB
8LdUm+WXrepk3J3XbNEeIXKuXZUKET86IoECzGiMb/Ujnp1C/X/fCZ2/iMJIQmgdDvqL36/O2c+s
/cKPT5RrxPWaUT4XfkL9jtVQiO5M7gecV9yOu31PC2FtWHmhPr3+/LPo8djAyKMZjKg3gO98IbXZ
k7+DROiOVW1GLR9F2PSbTDMMjgnPyNlctl1a0IV7E665wL1228Kq4ktFb03kfu0iOQ6iZ3QXdzS5
/fSSKY2PSBfQijWGBXXQQekgOdDPqUfrM0uX3KxZO1LHK0aa2ovCiAjJIVonhP4PJTn2GAUphjs8
j2+QHnBWOKCFnXNOz2Hr+ZHbkW6bvfGXVHG7SryXzzLtm+DO4e45U6pphND5eanVeQih3aC7y0We
JdaB0A2YGEVd4X/lgKGIRgdPZhsCQY49qO3esMKIq/6Wxf2BNBHdAOFDpc71qoL9YPknQzkmKKDS
bdoCwxDLMNLwohXUTNOyth/AOhiwhTmwx46wwAKoblmkW3dDYrImj46DAZVtYTYniEZ2kloPDAo7
4OubRHsKaK7HoPPGbr5RvZqtjKWlBx/VCebOZMyXG2GzCsxMmiKacxjb4F9qEsKdBJQBGdKG/mZa
L9lXQEZQ7fBREKA9HOSC5PaZrJgtj/JXsa9P9XdhcrbSPx96CJSKVmtZklNcmfOAA3cyAhRfyu9X
ynGzjiFuvhBQ5OUqwXIH/Et5d4KyXNKYZ+Wz9VCp4LvDkLxmPXRhdsbY4QIBYvWO7uJZIqOkqTrh
IrtTr/G3Oib5C57kH5ZKZymNkJ7JLm93fve1zJX2QPt5/wX1rMyDFA2iYFtjGxzYuR0V6/YJpbod
HHOmiFkjTw+ZTvbTedQAq3NQrPFb/rgEg7OuRTo2jUfKyFIKah078+x+IdKyhcG4g5mRj9Oo/BcN
Rgjk5ecnAbal4mXjt+8O6S9CsLMTbTVK/eMHusHK/7J4RRJ96cYAFfnwZJRoBouLuNRxufH1miG3
VEZKKKhwf6Ffft74nUefDXSMlXGk50B5a7j8HgEvk9AEtAOuys9FRacI8fLvUIbnDs2g3VgTOBxM
y4X6QxT7XXZbeeGDDSXelwzaNPKCAEcCbmX4dUqbLQoBdijsYByQ1vZbykicKm5Dwmg1/7X6rlmj
MQ1bJB6dyHOglTD8OLKPt8Yo5vA29rQusTSkpcxZaBRNU5zpk/0feR2t0KkHzlCuxzEdOhIIC1sr
peAXv6IrlOiM3NBZkrOG++2LY+FYuas8PpFoltyQrGBxATuWH/8DUokZWREWrUUbMVrYgTMSCxKF
rKkV1O1xgu83QOg4MYe1KkEKOO+4p62wFY8VPLstWsnTqH+SHL/ztt4ZsZ6y5U3MdplkwPjlEgho
9kkLZ38uqRJfO6+hyridmhaKoRSYTZEz1rsm0MngXDJvx4gLZIxw0rTuQbOV+BhzYeoV+GctZwoL
mfYoV0Zs3gHsGeRmtgdIyJp1Y6jx7ZkijW9/BuRf4AZACuLqAHsSflEQIaYiNVzeZswPdZZp2UxF
r8YLqQK7GqQMjXrx8PEwTpSJo5FBER/b6AABjuelyReIKaef0wHAGWmOraLR11v9N60Y4OhKLDn6
cQtGCc59YCsjR6M5Q08yrXWJTEPbSuBprqHr2BLsmCRKiHaa5GTGItFzgknX4dN8C9Aza2fEdKYR
HLng/Cs3TKPn3ENjn2qUAd8PaMEYqbVTtVI2CojvNt6HcpZn+1Im1iNNF9muMCqGUiIDs2J5PGze
ATAdJgGuCFfIEE/cp2oJsK3VCoFj/SJAmWPduMUmUWqSfvR5fq5W4ar3lJlpZmMT/ADg2LK64p3k
7pw4qTW/he6oVenC8Jg7X1keOmk5KkpeAnHO7HpBQTLx1rAgD3mrBbfFAwmpUKics2/ldbHEqgDN
fV15peQy+cgS/6+CNklWEe0MTR0hdsoAtc5j1+VHZJQok+lpqTKbCYPKJPUe2Cu7dschbfYhb+A5
kWhL+30LjmdfmH9vqzEEs6vxNozpEWtGI5xRvfOJHeqDjcOQBg5oy2tTpjpKRSuflD+EJFLljXYO
jB7D8q1IjsW6/fOwPs8JHFcMk+cuRIdCSviY6W9md6yhf+RjdmxWvAv4yJPk6ED1W+Y6EjX9fpk4
L/Jymg3Ftrhy2KGAc5u9/W7nM8Ud02CD6PMEp1JT/dCcxyesGTMr91jkHL29qthjhqlQ4ZaCky+3
N+mmfR3oLM92/uobblxnO+OUF0F8lD41aLKUArey/t5Wsk7Ird+woNPSSJc3mdGTu8XZKAf7NjZs
9IHNV28pqJgzwpOruPjrgc4HuGjzUnWWaeN8hkhnkXw+xueyo3J6hr/E/eKxjrdHLVyZewfF5VMA
Ibleqyh49lfwbnzJxRGCBN195gJlNlnnyGAjlq4P4fIxFBAubANj3wsCxYyKnyf1mEROWzzOJr9r
sHSWGIPfwIoEbdwufqOLNXZ4aVmBDVcXlaYo+YdJ7hP+gPoAXFmdQ7PFei3Iw1CYELTGc/08fKgQ
OWxAWFFgUrGh7SXAhpJtK17EtJQFDNCR6SO3cvSdifPJrg4KyVu5Ei91eE1XkRzpqslJiAkaCyeL
QB0FFLEqXzCd0TrgO6tW4ZSElxUudUbJU34RbaQ6/6pKaj/LZ2DtWK+Wg0mU+zjVWXgOvBFYaD1F
w6XrJaEcAVFnAP9VF0wL45KVeB7yHcs9tdB3tbrRRJpopTd0k9mNUImOdpq+ZqIal7iGdlV/YAAu
EgI9CxafE3533nqUf/XyYGAW5r8cOO98hLJvvjIfbItgeXGHNy/JcTOO8dU/F6ZV36KE/ZuJK+a0
R3EYpASLuSNxQw75XX4vo934BIErZRMDQ2o/3arC6NVSSr6ASdI9GIiTzROcaP6489NIaRnX5CS7
RcYC8gEbiHnD2/CWwi5KcqiRzRnDV1nnD1kPU9osLTTUhf+TNsI40py/eZ5mCWZ+YVZLzjXSW+a+
u3YHkp3nUUYeZLQJPRGPtpMPuUwjFK1jtiPHvoHPRx4MaCUMEt1oHFRXTJ7dp5MJ+Y52RdoYqNt+
yvAHuzxT75Q1q1bwEZ046guBOv0auE9xVn2Chf1bJ+aKf7G+KBN7rSCrlNNZGFh1UGchkG5F1yC+
otkDYMadvTWnH6jDEEg9fROzx271x6dYE/dAanIt5puMzVVjLnEq0FgITXLJOLZwTJzosteJw6hV
SWD6U71yHdamzpOKQNmIcYEd2WZ/wp3M9n0TavXaH1w2+SPje+TolHpbPa1zs5C/H+BkgAN0JwFn
s4VvaF9bRSl/ECXO4xPYxgxKt+/JzPf4vgSUYkYtp5+vF0kWlZsQ0wZW2md1cusMKTP1XNqMwL9W
AfOC22kvUtE4THtKwv9j2UAYexQIMvHIDW+6RIH8mvL3v9RxPNaYFr5cC1296jwa3clWi+Mi1BiX
xtccq81Jzsy7c8+gU5lclCuHrK+kk1FXGA5JWeta5jYVLCHNpGsx1w8gLYJqPJSTssQ9HbpTzHZm
CDla8B6v7A97QrEIcThTmuHk5zppBG6TNjYxXXmrK3ERYD6HRr5erEu+EcFfWm3ATD+aCNZDOvkL
1PZKeIIIZupvq22FUz5c/f6nwayZSh9zupLk7WPyNQfMmw95cGgoFqKDKMxs6KDnXkp0EIrD3sos
v+V+TChkviYmaSObvn3W6pWjKfSfozd/KLY37gc83vK8TAA8ZGA3dQpmKbz7wS7TnBjnTQQWBe8F
718iw8VFkyVRSmF2FVpe0aES4wEWzSw6PG2HawTGTvyKRMtIzE6qsIE3AnwmsicKZXrnUBovwwEk
6WxamAFSYtounq5BhKAK17lB/Ca9mWlOFOYTQVWGIDsHy1dH8JP0cse1oj9XPfljj6YaviSwtGYI
ZaFj+ndjqXkXons3bW0sIq35+84ATecaxep1xWBfo9ZHrs2Rk7xsNkGzITB9lQzDJP5O/+Jj6mYh
KXw+iumgmXG3hW54QAaLLUlbP81rPbRgLOGpDGjDvMdecUkskwe54J7p7ovvTZYmKfbuBDtKuwNG
EQDsIyZVHswG54H4YnqM1Rp2aN3rK+Pm+/RkMif/kTO46vNXpJs0I0MwxkBcTSnys+RaWrdPxdL8
6VBY0BLDsDYqZulkfc4/x8ANH4sAJsuqaphVM0YxgwRPazoHIbvikqwAt9ooNTbj0u8cnW+z0rcw
0fwS8OhN5zLinBnxlD1ntLdd201mVhazW0nnr/LrDRDbElXaLruJUtXguVZ0/u9YtOHK/9EfPBGY
ed5Qs84ptsPUEB1VbsPOFHm5fmRF1VCINCsPHVEheCx0FV5k+8aQu6rtGf/KtOiLd49P81KuDgMb
5K/WMw+g6ESrP1Ig2lNchiG1kESi81kIa+kLXtkjgRnkqBrvaU8lre+J5hGLhKKbCJQ2jYZDp+FQ
o5cL0dSapcVzLVdGkJD0PDhPbO5I+Myff6krD448q3CEmlGfTPPz/yvE6hUN/n2U45yIWdKW6fxn
jwGHc2MoigY0qKkwlTL7JtKrSYNqe/3CYaFm+3AwBLpjhqQ60vgKPGoHx9OUoP4F34hNbpZnOt17
qGYl26ybm0lcPK5KcPKLCqkvG62YSfIa+4j1nfbGGv+gCPi3HDIvQHpvaVBx1XVgTnOd75nM/x97
XfHe3fW1cA7ykkti1MH7PcwAtEsnPjQqq+YKiPf6qDtXepaQ5dh/5GeHHN9v/dSOBBSVTCMga5JL
3v5TdLVrURYqFj8nU5aEDwgtreljpMBJSK/Xk3MO3QYKgiySBB0QXIJRi8Izr/njV7hlQPurdUu3
l/UqU8SsN8aBvY5yWM8A8ZgpZoTKcA0MfQ9l01TCuWshoB9cBb3NTOu/KAs/GLSbmlam0MI2gE5b
btfTHStXu8WUYagiJ73S4ScRw7qKXE1P9yZJo/1Yf7Rs/HREnIDrF1pzVLe7c97uW9eoyVMr891x
AB4MImKvNM408+SVJslIlqwGeYj2P8L5zBmWF5XnsUxk+GVSHst3YyeXqtMGRUtX7NkRXPPpnOqu
hqnVDOh3SuQV6xmjBU0RO3TvL24F3RmWVpNGpqq+cN0RRUFY8w37O6EqDVHX3obyYH9F8jK3NZpE
xBN0TyDhv7th3FO1HpVubw/aofh6CcGkIxUfnuhWHH7nWTG6llpstRuGXBoEx0Scl3xbLqc82wMa
rqKkdylDzkAkyQnl1fRKdCLfIXCt1hRU24ack0YjTAi/isZ5+rH02B3SuFRjEPp/Q1C7YOKZ2Wg5
Fw3sT1TIdcPHrRICxkcX5Zh8oG5aj/wuAsMcbdTy7sjQqx4MpyF/IMZXP7dFXzKzMPnOyLBOa9at
tFo2fnH0kooNrbfIZDGoEgGpIH/zgih9UJMXXIEKmUyZ0YPAD252Ae1mwFKxxISYqaDswI4AP6+V
dUz/ggOg0kVgceFK+ZceG0xRVwaT59Bd13BkrPtNRWqvaxddL00rO/4JXCuXKHRds+cI2hM2huAq
LsCfBEi3Repjvko1jrcEu0u1TLj78LjYaHOvfGjHDA4Ga3eROlZ49lidLZugMfnYePEFn0C/9WMf
DYPlnEimm+80aNzse5JiNiNp5RMcvEmT227j+6PKptneFcmLnQqf1uii2m8Wu1UpXvc9HVXIVul8
8Q7qP1K0BEgGFtgdM8KJILHRo6VCTBbb8eH8fB137YKKQIOuglIcWP1Um7AST5/AkyxeRElFZHxH
hv4eIVrkHYu1Y2yj3ktF6zlPbfih3DdOi6qlSK9KqPt/DpklM1FTAAbLya51F66CynPcpxC8U5+u
Yrkdrz79lm/03mfbqynffPRpnVA5SW2PnMjaZW9lA7lP6zpt2itHpZDcvUPwKDaEq8R9IkuuHekx
GSDQYYs8iqoyRxzo8DQI6jGBlaE9KHgMpJx79/osaWDiGBDSwFDZ1T5tPlqQ9MUbwRuCBgAmFEL3
I4LGSIsUgBHHtbGULQb9r/+3h+SIAJa5xAkMM67T4pAVf14RcXkQKwDuUq02I2e8O6tzO7sn31ud
9ijXU8SVFuhfwqHeikNw8pW1h4Lo6l2EbE/jJlbegkJ7VW5CUm2O6p1p/Zw2LcXscpXth/YSe/ST
xjzyu+uaGZ2Y5sjxeLTIgw9rAK8xDodnW10ZVVc73MpPfOgXeYdytw4JBBP622aKWuKytu8E9JHn
uk2UAOEqbv33iQE0KQJIkONg+We8A1bLfk4zGKbg1745dUPh8dL+o+21Wm/KrtJBrkmFnW7uge0W
+IDrU8rzSnisTRxtdu82bXnWp76JWIlm0iBzSsoaBWCtteseChR+7JL4/PyAKdtUmhGziwMhvmpJ
fwFWO1SYDG/lnanj5eIa+s9ezluEEw6U4DzkC1DlnkgqA5n5istysyb1ehVv9uxch8RjaLC+D3SV
vRB274hB6hPLKyt9b6iFLZEWnP24+qnwbou9jj1T6agUTakF0iN9VvREDQNx3Xs0oWwDYlCrD5uZ
K/oJXNzYuBJq1qwWOs00XPn9XKYQ2P6bWkkPUXtK+V83pzxJUbz5t7fs7dQbxgttqySRfRML+N6u
xI5iyMjO63mMQ2xxbQr3kVY/cOsu6CneQXxUbwM6N9u+4UMy3KS5wtGGHUJsSMhhiZJAvEJKigC4
68CRtVDkvAvLWeRWc6vOICxhCiMoBbPWaktSZzjyQReKlPA7UVnwUqBsXteEXcXeUex7JCKf+EhT
pvLUFLFmD7/9rdHFoGGK9znOwd7yRtkiZbpmolpPv6pjheUvvdfDmBcCoYO5kFWUFMkLLVKg0CrX
MdGlH9gX4ZiF1VlvkLwvUSj5X/yhDuJ52k4TNlZTq3GnvGQKj+1geSXZYo/LW2t1QRhprv982G4i
QJdRySFbIwlitKIUaQ4jKW/Pz/Y3E65xgr/Ws55RA++zxO27AYX87F0K5agz2yV1COGzQKrGM257
8U0mzNAStOudfOwGYKfQekuIc88xEO9iDyMjL1uEOWGAM5AUQPz6ILxm0is0s0Bhr8CRfworgxC9
cYr3D9N/BrNQrEOdd2529zkJa/yrkYGxR3dBXZ+QmsoHDNx+jCAVcNFSINm6alCob8e2pR5oB9k2
fXQIwICO61uSv/YefssZFR4OJSAsAG0BUd7iCF7KriaY1EQnZKbt7+w/FVguhsf9NxEi9Lt6udxj
KIyifaA7+gsBPpycUN6SzaU502mCNzXYLBMl/YoyOSAH4y0Gj0HsvcSFtj9nutvJ4HtE5R11iba+
HiIh9aD4T1wtzaPHwEQSKWymZu2NHlq2y1jTbp2F4rLPpLTHIOw49eyWH173wrJ4xHXHTJWi9Vpm
Ny4K5sje/929/9yFYvLee5F5qx90HVN1s3k8AcCHd6q7kS0cB587XlNK1zxEwAovzirEur8yh4Im
+Gkkzk1Zc4btRojCHHUVUkqHCxvDKViJR+JvaCgMwTp6gNuQoTlEyXd/2U2+jy8qxstDdHP0tMHx
CLncPvuf/o4nsJ7j1ENpjgJJSAzlwucTcHTNqvNYxryf/+h+LvBAdxXZeordzeUCoOhFrkGRC8fK
qodESwiouiVz1Mo2kiTj1g65H46ol5azhdwCjLEf2xw1iNl5m33TSNrRMZkQNOMPtcub1AX+d0NA
NFZ1kIMBo5Vo3QN6QYNHUXnXvamO2zRMK0yCCykUemm9r1ryWN0pUrogW6kc6fNm6rtK7P/EE9Bb
/Jp8rfb7YtKlJfuEaFUeZXgJPxAdmawWEQuZsDm2QTNW9Tk2e18fRYzW3DZNoeFFDfByQoMrp8aM
iv10DAnSx/wYKjZpaiR5RYCkm6i8LtxTdFXCuam6bLG9vFAT/5Rqe7nEbWIxv/gI2NrWIcmN5akC
7ltb4sb/PNxtC1LZrnVwx5Wftnk4X1MnPmJD1rnW7vFHmdJKTeZaI8ktL57jE8AlZgKFmGZWqde7
fWvu3wMhXvUvUWDkMlD3E/QVK1A2jtY4gQSvW9bqtAytTFZjuTvsBDxPNN9wfHlPga9wKmVqCZ1D
L2k/cad8pz/+E61FWo57FgAfWS2CZYES9gMYColf9hyz3DmR/Ai8Jz1tDqzhQFYC5HAdWvhCOftR
m8IeFz38P3pOfk76/NtoucCb/i2+OZJqAWRbmeMLFtiOYgNLs7LIf3IKD5WfWvfdjQb04OnTa3xk
6nRAULKnVRwA0B4FVYvVy91r7ay3QR9TzfbVsIa4PVUz6tcbnPdExsHA8pWni4bOcba3r61ar4SD
FblhxaX4U7V0zO7KEcU/7NGycJ3VvMQ7p9H0XzeElSYWdGYIFjYIXENLW1HP3lhMXta8kXSTeRxs
fmlhgqYSOkHqPEKjMOWLuYJxJNnwl83bftf1mQI6BeqrTGBhFwA8n2XazZXJvY2WYZCA+SPMoy2F
AZ8oK4zyRK8pK7y/AhdfjvRUJ6qKah0mohs7k/0VAR7wjNzX/66J4/33YY+dH5z5ALUi/4ot/1oB
ALCxshUHNPJmTMUbfd3cCIAdbpOz8Alylo9On90a0D+gl0vDjyvaH1Hrt3fnsVnRfD4q/TWE5liY
WMuFKe9Al8dQUNPdZo4J9Tc+/ezLo8fWqaiqnWpZDxZXfMwOBh8v9lcmwIYLuXPsVV/OEfFK6vsF
/j7pkwGkLo30SlJ0dvWgRm0TJEdFmHeLnvv3V7IX+QRQ+JYaOYEU9NLNWKZUlsE5VU18v/OCKVdV
PwfhDPPGfsCRVlSmA28B8PsLBRydkG/tpYjlbCSE8i05GMdiyw1PtV0u0Ggv4ygQMFRlKG1p1XVq
5H+guRXPpQyU+Kbk5q0g5hAOjKoi/HUuSIdZiEJfQiAz7RMbAI2fDiBPrytqQFdivi8e7A/cyIVq
zkzYMMJSy9L/+jTiOkKVlsBkfnH0YHGTkjP8TH3wCrq953BirsuOmRLLpJcU5L3YvE90k0acX+K5
c6fi9Bs6gj2GG4oGEV7h8uIKWCaw0kVcUjm4NND51Dx/spUQuKX2xEv7o20AFPZnvsUybfh+W7w+
dOwRJHOiPTwYNC0SWhzmy5qkpPv+IrgH1w70PtdNYvK95rFUrPfYYOsSlKnoNWMw6o21gqX0Lp0k
mP1T4HgtBd5lz1hdXpliA/ZZN/aet+K/0nIx02UmJZ8JBgmvX8Pt3HDFvOwGiawgMDbvTfiSyJI1
cd7jJHB1N2529OKYgxJjANVMK+pzo7eLdiQpSuBw30iXzhlxWRql1iLyrDRLaDSCKO9vN9SOjdD+
X1snThLMkFoxsniyRxOULi/TF+t5n2DEWN/5ck/thGJkqzhV0zoXZ6d6JtrMLR4TgU1BvXpiVpnN
1l4T6gdQMm9o0qj7Sc5Y3+V9X5gFP/AbyYH/DrJs3KavK5PDt33mElTWtmiOH4hgx5jl5C2WKAoA
UiDV2/GdYmHTDH+G2og44ahLGbHpg8Az085mhDBkiR11GESW0jbzzNfZ/FzAsCyYj5eeezmDmzW0
yGuN+q4RPBPHW+3aJgUXGLDeuiQZ6jrehuPMy/eFOj3nRvTxRxI5XoQt/prc+TNi7ia8z9G/Jt9p
gjvJDHmpZc1sXhbPE+jSBTcsniuTvOEYG+XfVIii0ahxjqp+UCOVuE3pCpvakTINaZS4EbxhtrZF
RjXkeXHHH+etQTmjWknTwUY69zQqcKiwvNwtBmEAKd4ymsR1Ywczi+fO2+ilyHBfgt/JNl1P35aK
e7ooIn5GPIG8vKTx9A1h/Zx7uAa78ibzln1yptcAjSStPIMELnEVbSf90YTLjwGAF5iIiGF7e4qi
pD5IktVcP4RbYAmSjNnyShqY5Ji+8mQyn5JKhTdKdQ4MR3bC4ISfyCYDANEOyM7ED4TtA1g1wTCR
OBkKTxaAPw36PZtINbturhuZehPC6hn/ztPtBRuA6HDmEwBcDwfd3W4iCdVSbfu7+d27LMAX0TkI
J3223e2kXXqqNmJ4GtF9ZPBxYJYdwpn5woFPwvh+/FiGDuqjK6KU/SdWIMIvOTHjJs1syCBc3Q1F
7ppx27ovQ17/LG7zsEp6fxUy/FuvzGsv+lCfRa2oWuG4oRIuSk4c934cW65ATyaj/JW5EWZKLXl0
lTfi+5DRmN/2nN3XvYNK3jE3ZuPMb2odq9q5BauQ6jINGqSrBoBwqAsEGR6QYgkz2S0m96h3Y4Jb
zbnIfo3HG/7oGwCcB3xoOsH9+lvM90X1ir9Ar6Lw4HLTE8StJ7MlN6Tl4ilZ03Gx4GfuDhDNhGg3
XU1VBZWjye7BoRiwPJM3Eb2aZOSFNLj2nSkRmzqHpwQ6HLTkvKUgGOD19tOFfzzN77LwbHNBEWee
NoceKUNrAJqygp7e2R6ETk2CD0AlNFbfxpwAvnuaE3Kp1AmAtF2PuP6pzVrDXBCxm5OWrhKQY0VT
gyaTEs0gWD678TSSFHO4EBWD0fGhfJhUNqv0AGaUTRaizCv/xgMnzlJchU/M26V2OOjCURBC3PYl
Ii7+Sk1Q5nXLaR/Np4Bm4+owJD0KS9eciWZZVMnAhlsm8SFzl26ECYTk7j0+6y68flBFSta05iuz
TKEfzXo2FOhjj2QoGR9aMgf3AVrmlvtqR1FQ1H1hQc0nxK9RnV2cXidv9V9a7iJCoybXL9Qp25Ty
jftpeKWRyUSP+dS2od7BBcgny1PpDinYDkgT+1ckl4FWfRoQ1fP9agJ92XoJUDbl1QB8aiej9UaC
Hko9OjyBjLBudyOJjo+aZBHwMIyhxrxl/MrQbplw4EVuFgBIrrc9WmwJR/LuUfyIsn60F9wEj4Bu
AupgWX59WXmywlwXbUIyfxCYbfA9H8918+WZIizisW/OW7tlynYlQoqgVL0Ead5lv898n4aVQdqA
/vkD11wDxWC+qVJFJJuLMlazgJni/4fT/X/nxPVpDz5DYvOC8sb6Zvd+oeEtb6eHXQmQxyjldVFp
mM11AoH3izLcJKNZEBnk7m3ZORxIcCdV5B/2ZLselkaib3ONBq710+mLHFcwX8DXMdljLRuoyEb5
UkY53435mz4J2QM1Y4FFZcmc1L/uFBf6FBm6mQzyH+Shj/sNZj/MCrqrSCRyPfgvoe9eU4ylfmMY
atGb8OWX5xwY67I0Y9ZZ49JF2Fy+SAHM+SaZBq+/kDsMlQj9LQWi8unctUJzT0cPCJLScTWchEFQ
2LnZnQPUT3kdZG1QlaPO6MiV+Y8GYXDAvSlpAqYV0sA/aZ5L8VkmqHY9rik+EWtU5DjpvXgHj+2x
oQdJqdCkF9gBnAAfx6ylLsWo0/eH4OE3wYlScAIpV7I0VrW8N+jFkFEM2X1AI9mJHiRtYZvVa7x/
rW0PdA9kaCe7poCHV2t3uUWeQLTRxkbv84Y5NmY6+9sxti4lP+QqRHYNvPGm4EvqkGyDegFKdEwq
s3xwWtEYB2NoxHx5dm9Kt9UXcNLZK7InPBaK4XP8N1t6JEEpNgYBmrSpNEqpIt7aaRqrckMnrpKC
fmECO/9Ju3FKUFmhtG7Au6DE4tOutAVVLd+6kFSlIjrq0b2yBpaJ0sLRqM+NUUVPw/RVNA02hh87
ypJfTpdgdm96M2wFLinToIftl0LVl/8cwqX0SqA+p/MH6m4CnflQuW2Gv7gKEwm1JRIBBko6zdnD
A7cR1h9KG3OLGrNHj1MO6Uk7vf1zfH9O4snnGB3O/icrEWAK0ETbT2k5g9CieG0SnXeYr6Mor8FX
YuxaZc0mmfOF1du12Cn7uyRvkkA24IVpjIpCi4SkDbTk8BDWott+krnhxHUZLG29Cww2sPu1DNuR
lg4tgzkdRYZJ7rvOzrHRJcqHRkrdGF0ktlaifAQ+eKVOqgEUqRC1ETUFwYa4jefcnPKgA7TLbY4T
K8V78T+MwwLfBpY4Q6fl9RDZdzIgf290s8OCv4kabFdwka9EOgmbVY7VSvW0Bw0ePwMn2kee/Owx
TAJDD0cQcULsvQ/VcKBOkpAF8vbQBgp+MUSxfoiKTPT5BkSZDlZpDRfjE7C+li76dZCtJlaGVBDY
oxu/LlwApxe7uzG8k76eBcFMMUlhknqn7BpkU5DArSnsOHqTwQjXRrztvUEerdTxRpE3BQT4vPWz
UQ0/ujH9F1fjO/YHUDFkArYCBvXVrquiuK2is15UWHAgcGIVbPEQ8S9Sjvv9ASmeZRY8acduAufA
KYrXsuPOWwwYf0RYuS+xeiFgIVjTmPHwSzVIxIdekDcQJq2mVd0wDeR4OILFA6jahjMFaONSuiLM
cva6qu5O94szWyt8ZmaTTu0j3nxvIgpEgheZg5H4bMXxal4+fYR6qPUVOp9fDtojsbbdUejGquaQ
r2eXGVH+sF6m2d+CZB0HELLyMuO7Pv5ze/OXaW6GAat9ipx+N5KUkYvWhA6usRY3RiEFpuhktMDw
2h0pLFKGAUz7/0K/md8CfmI6FAL9ZQbQHJysp/u7NMzkH5BmDopZeNaDwi9umF1fC+N8m7+pCFht
GIztWWYtdyqN6Mox73958mcsdVzYxC5xwvWz8cyrMaDQgyV8ZZScI62c7dxoSJ3w7qH5LgTbX1Gk
SHAca1FBzleEEKWq2L6bjnx4Z0ATEfzNSOL+/Y23WPKWO76mCP2xdkZ9Xl1hLgJCmX47CMlxVmXr
2FRC/hqZWN5RxH+bCrEDHGH7hNl+ud+DYnQGRklR5S+pnUANBe4v/r1t25ZlsRdz5WcVsRuKYpdx
7meiCA7kzBewZwLw0Phd6KkYPqHqdnmtWuo4dd7Vud7e5C4qAYg0VW9hMa6ETXNr5DfzkE8q0EFR
PW36dvFsFNoTcYRCU5HK3Jg6CHX9SqSgAU0GUFr1iStSZZN1KepvkO8ITceeSEZ0xRTXfkGokzJY
p9kszs3yptupD4BjtNsBiNA0M7PthuefKmugDuQFRNp4CQkSMagGobBrrDXIqu5o2NDo7wZYCGL0
d6TcAOunPawpMSB5MHbhYNgSANHX+fvCfOxVNDQoSXULqrf/AOVPPsZwtwtgCaaQ0+pS0vEVN2XF
8RpLA7T1r49R3MVkId6OE2niKEm1qdgb2L3t4N+wn8zd9cqzGtie/wIwnCPF1yF7Ke9o51d8Cft6
Uj1F2liIJiPdA9n3FfgZWCDeAHBfyulFSr/aRFETzK0MNeSUG/OX4RKtGybu5JWf8e6srV0awkT3
hx+Efl6nKm+WPu3TDgXRqKEzHO8Pb2RAvfZ0RrAGQS40BmCMpRVuOo49JzaiKg8IT/OiFDgap0IA
mZifOpKggVqmnjiHZ27B7qPxl1070bhuZS+TTGFeNGuLlJHi8KqRHvm1YeU2Wsz0KNBBpIpt1GQH
fAC3LWobO/i1dW7Jyl+4Z17m7GM4NnCWvqVehLVrhn6xOa6DMFkS5KA/C883z8YC8i1WPj1SJMHQ
k1tAbVnIO0HKSh3OPJe5HB23LMXkktgQm5bKFqABnBkCQKwnHGfLLImTPYljAGUbMKJ5Kin4S5Kt
pnq48AcjxKt3B4fWsEaX7dYJ691rMxMnOLIDkSEEBCdPoZ17jC5CSZFqKBEX3MlbduXMiVgPcLfq
yNmafobdw/FJ6Ih2ULjDClrQQaIXVHWUp5yDaPlxA3ONHmKvFcHbx751n3So1jutGUJwEaQAZiTF
RjoHG9aoxOhz07/kT+hiZHsv483mODK7Y8PAu4XeAVPUICfG51NqiMpsTLT1AA+xbiuvzXu4DIz6
40qqLU5EbFlM6NqL1m4SjyDigRvFkvLHMsEnE54s3jWjmUu8BSMm95Yq6ZWF9RYC1d/3mpFKIvVK
ig59uSMWmIJj8CPWP6caZ4MXATLkW9HFZqr3t2+MANy+PzgPEu6+7MkjZMxqFEYhb+WrDL2P9a/d
tnwKE/CCn8qhpzWFDafZhXWpZJMs3O6hyjx5OxRebD5S8j1wTCt88sl7bejoP3l+PCDdiPBOXgYv
AAQqUYeQeYE5/J1aiPx8osWI3ZZLS8hrv8cRajnZqj6ZG5TzCCXm/zie1xj6k9Mhtl3Cr75a83Jy
3sv9t5MTlXLZ12Tgko5tIAVJJ/O8njScXaz6HbkTYCmFGN2S1WaV4HgL6DlJvkm1TuDxqSET/567
+mfHSbKZceaOQAFek9DEI4yZ/Ulv4+LlnPgMAHI5IZhApyxRjIL76NT+p/Lvodfy8sWNap1KhK3g
CHBl/hZucaGhjLk3oLeFrk1UyXjYovmFFs11MUXAP+6qca7JXOHN01MUve7SacOBiqnaDL64/hy9
aIgKeViDYiPe5A4uynlzAzzJrWFr345nPSgQ7Y7kf53UPCaB33VaEzBNX7NBaITHfdHlubAKZKdp
HkOSCEce+v2DrW+NpVyis83DjF5UHb4UaWsyHM2/QMmX618CYXyrEwIBI2QtzIqzq+Oyk3xtGWDD
0kIKrQ72XsMarxtcbGW19MizlUxSm6jppJbumHpKdFFXXXwFrX3uNlevLKMwipsRZUxzfNJMMTyz
u57sq8thwAB2Of5tZH16XB5VwOlGP1I2kWid4PZQ8ylpLdj4aHgtFRzX1jsm0To1s8avwSf+RgOg
w1Suiz82PzD9JkpQrKipYjcBhxWOJaT4LeavPUOOEYUVPVoUfKyUrcs/onmg9HnobPfbeRYqw7t+
h1rHZD7dqECY8704RLbXN//7M8zMpuPKSdCI/ie0bIEPAp9lKODcelSQUZLWZL84Zbrd1JHQlUFB
GMKT6JcX0CWB6wSnat0WsgEZoPtLX4CMA3JrHwYUHSt2AzEPm1u/rmEh+ybgsehZecthQK0WpxRf
jO7N5XjWIKrN7r86k3gKNH+h7QgWotX8lNeC1UgOZfYU+35IBOYHNErit5xqlqUNsQx/ndTrq21I
VN+q0TtwHmXj1DYxa/r9oKbrr4jwXJE6PeuJfy6oGLQyONKKyO4natkhCRvrU43N9AdepSGOquZ/
6Pb2aF7yRyQ4e7K+gremT5440WNcYPUr3GGUdCkoGv3A4NHAK932ZsmvgOOHeax4oRAT7UruR/2w
cmo0S8j1fuZpeshChkbyD03C/DzHOLKeZiZzwLGnbuMU2eHWsVegDWk+2t4rYfM55k+SNhsltZWr
+A+gushNLzObUE6/hBF+ITf14GzthrG9mwcKGiVZ6GVkjzmXukq8h8iVXoSkpByQ7Li3T47U/Xf3
EpsU7JDNKrln6gha0VWkXeIvH7xhvbvUoaOtjqEoO99Kmu8O0/9m1PNpMJDZ1mXFhF7uXk2Unsi9
3Ys78gziH8DMUsnewRVkXo6x50ZfAuMcJOZd+u48ZCXRDgGPG5KKdUsAgwcREjdiq76X+5myNlt7
Ynrvr8ltx9eJ5U7jZtAWmD3/tJIpiBZWX+DQaxAflEOdm2XZwo0KbshVRvks8e+m1Rss0cakO7aV
Hhj1Dn96B3dg0rPdOuSiwt28z1VuE5bqkNLG8moV94O+0aZJ3OXRSVX/gzf3sAPyun1RKL/slO8L
szqUZfL/DEDSuF0ST3nAeqXWOa5SO8Z46YE2ab4LgBdtL4MZ90wcapHillHq3BmgQHh4Qx2IqrWg
YdJUYdEICNPhSuWHvQBpahT3YhhrseCRyZ74KVk8nkUBsfGnH9bvb6umcmR/6PvB6AGVeMhqYNFT
7MMPMNrEWwc16G/dRJvDRtYVUj4+bMU+TRlmUZMqod8gmj7J6NUPxkC1FjC/xeicHuQ3acQYpHL2
akPijDrXtZkzaJkOVjIvEMxP8mow90U+PvIpiGWrUZuCxwI0A2lZs+ncvNcMJG1uYZlBqk9wWfGW
MBSoLliLkWOKlJkrUEjUpvo4TUZfmiZxRx5S+nUt3NcJDXPDbIP6gq6FDD6Yy0cPgRg2Fx5hSjJs
dENYj/IwOHWxAqhVlLXF3WhsPsYIAM0ex1KEESEjxUpu0/Q8V/gfQTDKXqugdQKwaXXdffLczkMW
US68RT1g0aEHfqMpHGvEEfHEw5b2Hz3tUuYz+QIr4zPTfyGxQ/p3lvCjMA2puVqJxriCKli6Llz/
Qej8Kzq5MdkQZwGUP8fOmdfiFGvFGAmTKxTxDuxJcM3W1yRX41cqT8bLxGVxXous1oISnBIwONuN
XLs97pfqk0SVw5zsfadWhRUtoSsWnTcRFcywYTM333RhutcOj3GKGLvMITkO8h7xHB9BMobVSfNo
iFUydgOthOpeVEc/OA1ZxSVpM9gA51QWd1gw1hqoZgCKy0oWNcwLhhGvMbT77PeDThcNHZIVOWUU
TmeRybXyzlrl8JY5hxrUXusXnF57iU50oGu51YQPw+6edi2kPRCzmr21OIjYj4/bS4sgYlec8Q61
HcNDSP9BdhSd8nJs4ZYVTnynKPMFuq5dCo/eFm0SEbJSfF0TZTC4CSXOWJ02XJ425rS6cvUyy+vC
8GkmSS5wUMKLr/rpZuLaqaGadTMQzSTji9EoPbF3ObQavhzpE/PyCb1aTKAoFG3QjCwSn0suxCjA
qU6qRFIcTr7K6hGNZ1kcIow/PXfILmXYmz5VH2uUGGCvqBpxGxjv9NeW0R61niqeeJ1hP8jpl/sX
/J1gQ8GfvlZbz2uxW5+Q5SbgshnK9NB/5GQTOlpCWj8qmGj6E+F9AzIbziKxMPW0znYNgSJ59Md+
kL+2MqFXKeKwbvoA4rmhwb5VrPNmXMRqL5VGjMDrlCpjSRTgJtXQtg4IQPBNmj9EKrfk1T/d3skj
3F/H0IN0BKb2c8AdUccCfwBxOxwsymJOZpQTrnduiGjKeJ3HePVcDmH9Tvm3NiToJx3aOd+wbg3l
cwY6eYXP6kLp/d6joKg5/2u8O97MF4FT0otbtDS7YbKJOUrrL8mgTFX2qhgabXy5H7pR7llyxax0
hUneoQFwsMreMONNVKIQNgMD4/fQLatsnUwjyuOeAHNIXsCv5UT9VIKGfbFa2BpDgTL7Gl9NuU2I
6wPU7lOvmTYj5O8ghVymvRgQXMEn2WD7IhlchVdyl/qiq/U3xAb+qR+dv3x108edYY76eACfUJgK
4UtdFbYEndJw7kJuz9OBA6VgvVP38frCgwpYZBefYss799EPAso7i/wrzBhD23vvYLS7zrDcYKLp
ttA6cyT2ZXVChI0D6/z193+JTSirNMPZ7Wud0sUS5O2NrFvrODm+p7OmuC6xaBMev0Ox04OIUtfz
l4Rvz13EZhMOV1Y3udOi4XlpeoyPLbhBGOxDbLOPj0Xai1gMl4piNX+Hp3NAYNSvGrXAqFK9aend
AdLgGB8sqP1nxMy92/ny9ufui9YYtApcYTjsQI6yP06XfHukrL1dVjZuyX9bzPBo3KppR0nCReCP
oMWN8drQmz74cXkF2Ffyba0J/GNMVG4Uq6zstZhKUD+ly3Wd5FQY88jL81hAjIIvDj7CzEuI45VK
A82o1L5wMWZQ3tnus9G5lDHb1fiiolHYzN1t9lkXO6PWZC4bHHVgvI1QfrBKsgeRSwgPR/bShuyV
j7xPMQ+QXhxGtsu/sg98KFw+vEjYOZY1ab2AoAeGdBYj/FzDZEzXCrXekbgKQvgFsTHZM+80U/j0
uH9GaRuIMZUs0cyiVf2SYh02fi+HPaIveA/OCz/B/+OpF6TAzVqL6sVyfPdKaT4uM61qKXhlTKsY
k8qtdasXDLFyl7Wg5D5c2JBEibfNMJd32PHlroMwun8pdkDAugFhlMQ+r1LX2kS8vJb2jZC14oU1
U5p6ItgH5tuHofXS/Pkt93kGkYUS9BAVuQRl+p9054mNWuA+BPp41GS/JvdM03o6p0y3g/DVFalz
ebgzxyPLLV48hqQ2J+s6+1COkcYTMG+elgWRDdDPezVkyg6tgLlgn4M8WnHdj07gG+WQm8uWjuiG
fGOAJwNYTKh45hTlwFmZDHwVKQk9XbYUfleDevyDQB+dnTXE8m/q+NVJJy/CbP0Dn67CtXi7ij+B
newWphwKEmcwQuhxDfCwk62R/2XNYIQhSlu7TGlr+ZuvrzM6pgA0BHV+/V6to72mGUB5CIPx2FqI
jCSyPJZ/uIgdPOcUGVrHorfmmFzbejjthMh0HhAOOsf3v3EqaVhha6bGol2ljzzsdjMp/FeS9s0g
AmTG67LWuggCYaBbs8FYihMMicQx6RN9fP6+UPYv9yD14Q9kKILeifLt6Zji4t6KxViJiTx/Dc6+
EAeYSspW9VEq+qGwaV1FMnoBrBZBj2anAnX4ObNEcddHEkEzQuT4HYEun0BKAZxV5+QmQsYU0KBQ
Y+sjeBi1mQze+t49a0qdwqjALkWSPo+00bs9EFf79puteTWt3vweyE6xY2Xn+4bwVWTDaqjZBJP5
STMkxQAwt3P+rSpWFXSBh+X9ERrcWen3TNCIVgcQKMzyLDbxK6NTM+spv4dMJQYuae0+GtKQvaiC
3BQgVKNtXIVxLbDOaUttj1BW3/UtKnesEzX5yiSuAIeTBvHv9Qual/NahlDBsncBC4Y9l4Vmp8mP
lmchfsXLpEA56z8ehj6iodkxGq1KPk0V3AMcAmjaf0lXkKYcXt/i6L3MgQt0LOlhe+0IzLB7rYY1
IoiZTYZqLW/mJrWZowJ/zMQl6Il77ZEpjKZ1tcFzrwWsX/zvrCObZwgZg3ifs++C20/A6BkMK16u
0gB2h0fyWxiSFZaZBDU1eeI3zCGRAA50aqL8jlA6NAoXdW8dGJ68vj8zIv7r4KU8XxgImat2hxTb
CRr4at9QXfMxueONmxV5IbtBc/BMR/f9NlGAJi/ETcVsWXaQ/Kh0td4jHmx+zk7RyTFCicgnl8Cq
YF+cDEVP1zvqkR0wQS8mUEiB0OWQdRoyXgOwlPt5+v7mMa20mvRaFr0aMsgyGBAG1ypppkNzeDLi
GsXHEUyL6AhQgSSZTr9CvBSnqJjubFGdNYpoQXhNHjMhK+ipwdwWbo/TYSl5FnpfVypzDdKYzInB
qUa7CMtwBMOdvg1dG49DYI/WUwClaJgQy3P1mw0d2b2cYuxXNwsF6FvaDPPEPrZCmbu22dncGcmC
G/V9sDMtMMgdJBTlI5FF3cntacTYfpXQ5jM4/zMujCc3EUx5gjBPnUmI6zetnw0TY8NRoYfSQ7jw
w4lK1fEvdtrjXKjz71/WRvO6hHa3BOVThA1xRch936bVpxTNJYgY79DCNGl1DujWg/PQM/eHMBRN
G/E6QrI4Hhm9/lkA7U9FVCIOm+i0kcWQU5Zyyy28w+joTzICP5ljNy61B8HCpd5CkoUIKPPqEV55
Aew23VENSEJxIgOMV/e/A+b9XEdNr4yhqTNerv8TI7dSNI0o7pNY5fuS4ocu0e6SQIOODYPJMCk7
JAOKkHOJpCTOuvXSCg5Wx6//eWQXa0QwcWULJca3b7YxrnJHEHuCcVjlWIRmIqj+uDhhPu4/p+/Y
zexsfEdT6Yx1OD7LHaOjkH/B8H57yjWTOrvF7r+CQNqRufgXTyM6d0F5K5dcJGKbQecMeZ8UB/Ck
NmMUuVO773NEVaV3XoRS+FMmcbaz+jPyVO7mutOFKjIJ1lEcs85mPiJhHVqLNVV2j7vhtj3xqIs6
CSFb4J5Ual7Bi+Cf8nUuzSeyID0dXUemAVEbSfOtKsBq4UQiXBQ0qshEl6s33ZzflP7HVG4ipXzl
boEYvh7yPYmXTV9bEEUBn/j92XJb5nuS/pggepLuIxndjXLbEBFsawn31lJUiJUdP4crzVS69dzr
zBx/FE0iHUobM7mXoqiAZcvCvXmMlLUCATfctBqFg7fgeN17UhMg4wMgk3TrYb6JA1xoSn52MJvL
eEfjyTpjMlqsRr3KvMC/29EAiET4TzJqbmt2mZtg7tdY2jBCVPT6ENoQIXbn/WOEfrHccm821jNO
GzJp4B8o2UAYQbNx/hqM+Od5eX3xgrNBIp72/ADRsyzl/bkTXBa7FnCvhzQMQjiwK9nsUZuhU5DT
RLPhEh3per5XoDers1OJxjFTUq5Z31ae2IUDWOhXJX7j5VD0msYhbPJa0xp147HpaaV0G9Yg1KUI
UuGyQ4mDpf2TClkNLEBmV+p+moyBCY0zQzWnvSN540UHvrE5AnUQ7EiOEhlcq1J7YmdzJcfLI7MY
paxQuD7w4aihPvkFHoBIrnHKzirl+77yVyAyXP+qQXQDZRSoGnrsO1mhOKTKGeakeoO736OVGF8O
46NVaOsHH7Z6aKiKoIDCYsah0SpISzwq+TChAw+INsixziu74CD4lGOKIHRUqFNTf3jF/+/isndy
BzMQbuVdRVxmCHk+Mt6sLJzewmRVAM+dXIYzkHb6tQkeCUSsOo/GIDVJO+FZVuUBglw+W+fsOGRP
dV4kLiJ1FaDcv+FRbPpnHLUt3hqtqNmPZ/wVVFFT5am8+6M5bBdXBoIzkztHTvp3GfodK6baLIg2
eQCpPzltuWknVEIpdL37ot3+S5KVGeNG29bc064BpSpVFLuauZJj4Hzb91SaA+qgEOR4u2iEwE92
k+74d6On7cmz3hnbiNZsh+KxeIw+Il1J+Jpx3fioV//ESGEBD0hX2XceNT8uq42TUhwGZnVkh+A5
z9ODerChvj2k9z/Bd6SBIusF/GBpL0jmyrML8yizax0X2aE4VNDtqMnS5nmL31eG+Kzrbt7L4W3m
ZpYBQ9QYIM/d2P0yzAjmT5z+2pG9oChYmVusea5Zc6JdQ2ZPaZGiUsE0G2VSEl2QiuYwCBatAmuR
kdpzRUKeKk82kW15TnzkrZB1pgqM6D712RfuB3NxyHpR64kkqoGR0ESZivnJfC9YXxLHPv373CvA
H6H9KDZp4SdVKBFWRlS4Kt7rxyCRbyzxji5TiWlkPr0HR+qq+diMwe2Y/vfxfJ2GJVOFEF/Hjx2D
eYw+uOlu+Te/3Hv/baJw4KV4f8viC7M/gkQx2yvGh+bd1c46LF3wwvHM4CZB4LRv9YpNguPb4Wr1
CLJ6AyWDqppe1t1w3v5OPD54sBA2vixbJ6qsg0kwwG/wmGJw1CVBf0Q38zKcoR9CrgzvuaFWzxnI
UE6q8uSXfki7sTMMsntTDr5JKoiMTukLSR+Yn3PNpV7IJemVsmoYseo2QbbsStJfhLSu1sh6y316
nHUy7ZsFtzkNEWaKa5PGyAnHp26pod5U4hcw+ijD692eoeaawNocRWTXNhAE/+wdz6DgbMwcHVBZ
MNyHa1lT+9zpTlMwVKjeHTuhGtf6PwtjdVqzQAsktI2L3TFBZpreufSUiUk01QhYMFCPMcdTgtkx
ehiJ2LSbKG+Hf1AGzsu4/vfVQn5Ewq0EprF407fGfpGI1mb6MkPvh+PuwGG8uIXMZtK4gAi5itk0
5UUA3QMi2mg+YYjFozTBrfBrIlXmMwAwqIt9eh81fUVSPKBZoHz8IeSbqmatHe1mcOXiRYJ63o6K
dheCRgGolIIr1Lg2plFgkQBN/KxvMwmZbvEyZ43ROMBKaViB3J4G65FZMOmoVGM2iSkf+fEQ3Yia
dSI+UoFnq25lDzBezHc2AakNKRkc3cV3ew5H7GnKmIO6LCK1J0zVkI1x9NREOz6xv9YpU1e7v9ru
tdxhXOF2FGAFvboi5Ut0kWR/PoGEIXuemz2dqi50mboX4vJsAOw/DMeViszcs7iUhFCYs6ERM3Wr
AmELWPcY77lm3AvsgSe/SOdt/MI2oLQAc2P/iIM9Zd1gjgyArgwYJKNsupDbrSFv+xRU+HvYzW7m
toplJNWJmOhuVxVtQuLaCWuLFhjTStZ0WekuJ5O44WyaeQ3ISh1IoLYNSOlmlfRoKjaWv6OFRG5c
UBVTmz9OF/HYxPu8dOqD8Z5RYT6n8PaaJCtILZDScPFaK527FWxkB/asQ0uUWCDUQRC1ru7pPVCM
Kprtc8U6W3fnsPd0r2fcf7kjcVTMF8nATK1wuYOouU8h9P2VEFCicyh9+6adNNs9fHZDhsNnE6iB
XV7B1tZYFJ68nFRy382W0tFlaCW890AyALvjvFFt+hNuVnjTfnlCKx+monw+XQbkp2ux8l7+NISw
kF59dmmdMTHM904kd0Ma2YxGDnEn2MTYO1kAg+csGq7NVNSnygfEphvceFUzk5h+a6uGdbXB9Atv
zhRGVAtvD2SiJoPiknTQcuKx5T6nLz8kRchc/a+SUAeavfAeOos18FFrVhI5TYC9IUxk5DCFkz+B
EP9oWNnS8YEIfFMm2s5wo4CDpY5GyVmyljwhsMYomi+ZDpvfESoSVBDV4TbRAkoE4vOvOXmXMkrz
W9Trvek3/Vzt+dV2we9dULFHwvN+PUTAUsZZuXD4mJDreHnUIt/ZMzOQrYch9X63eHdV+lCpU/Us
1wxum89GujQj75BtIpXG2vusloh2rVUvDQDaiM1mjoAl/Ah4UIuAwcXK4MkxsZUqyKTTkJoncUrO
dxC0h5LF5OQc0vIbJGAbwLD3cLv7OIsEYWaWGe9CvvYjzUEEemXFuXEX8iDGU5doPom7OSJ58aNm
oWn7rzSLZJeNx0rp8xmKREcdszmsSZ3Z5hh+vvbxNC8Ey6ZmXkoD82QV2XoNTnWHNBDCIQ4mdjjp
xYXGG+4O/X0z/87k3sxWKOsOzGn7YD4YZKjVAE0ZXItatYVcVfmVYjq0lDSX9eHkHxIpwzvgcfyY
WHPc+rtAPz5KnCAcFNe0h/iFcoDgKkgH80H6WMsUaH2dZKou3edfr8VbUyzEog9QvjFRDT5sPeDe
wy9sSrVS1q3kTlUI7efWDQ9GUny+jmphivEvAzaU9Wxgdbndeq4ZBStNnCHrCpPtI8fnT7+Nvu3Z
iy2n3wrgNGB2Trk5Iw6dCveH61O4SD9vmEAoFciWjIYgCepoDNDDt3W64a9CyvE+NzS8IxMkOxOE
zDDAffRB5vt9gPvgXLD2pFud5r9xn8yC+B2TnUA8BOezVuYLJXDI8fViQo0iEsjMDjZvdfOjMvBa
Mcfc2YNiiHNcEEs+F1kzmvfvZR14QzdVugdw/Fvj4dH3jPxnR/Uu5KYg8T/1of3EK6ds63w6qPJO
PxVPYi1/BPSfJL/fg79ENu/UVmun85bPtS+GsNZGFYVe/cBA2i9YhfPhfErOEqhC1MsD08sI6Y7X
h0vS83Z/e+8CBX1y/5igOpbbbZ5vMbqhaFQoK3tk672azNbClcuZSPFJYKjbQB0xeN1pVxRTvTpO
Tc08FWM+q5XTgd0DkJQzR3kNdcvPVdO1FPNjmeZGiG0/14Gx+ekXaXlqfkWu9y+TH5rlmF0tCdrX
wfDj4KInHenSVvAvMrJnD7iHi+oic0nKAABQc2BIX9aayNBrKd2jBTQPzKikIrGJccFhs7qMHzDV
7f6thBr39ArfovZOCFSu5RBA1P76Z+PKUjyk5dZ4aGmF6Fx4fmQJDS1BvW8/cbwzIa5qp7pY8iqy
1wCRnuEEurudXe6OpiTvqzZECIWxSdjZx13nx57Q7uhz2ciVclxyu5oXTKUDafnl8YrcJ78qOINn
2R7rXTC+M1IZCSHO6AqxbmBjpE3CHUHVuL+stg4mx/3K3BM/wjYNGZes08U1bxMES6eMcwW2na5J
Pwk4dwHshm4oJGgGgr4jxA9AED2jzuZq0TNbpH2cYodvCoKn28pexKNWfyHB0Wl8XXrRmAPv9LUH
Z8X0dV85DO9QV1uU7V3FujnMsIOO9SNhF4M8Cz7V6wG+Ix7Sb1BFAc+3tsb0uu/DkfUaSAg2UOxi
CuwYCwx7GP8zHjdPatIQ3bFcPX8uvq/BUukqP3yndPi10Tk9dn2/GRuGsGYNV1xZ/XuXnKD6qgNZ
O89nsGdKDa4lINNVcQ2GfNbdjjVvR0XlodQUovsatxnTS8fDo9/QpEjKgl0ZFBN6YuY7LXmCSNgU
KSypq3wjLXLlVLyB8143eOpU4zaVaaNbe/1UmUVsd7eV4FKlj9kKjI5VsowLyV01rq8Fr0lKJCBm
ECNSGOcgLQFvMimFVmm0S51Lh1YoO/C14H35p/51HQj5frL0QMkC9K9Y2ycRKj8ZHqTGpoo4Uwv2
IklcW2XxIwUQgEQe52MibcgasYNFz9jJCIrdigh88vjSW6gdPrZm8FnMW7RF772eeqXUkiDeovwt
w6kkXv9YAQTBhqRa/7KeADrB46T/zppacNOUUDnmHDZhIDXfBXpGmI2ElMw7Kex882vxVfUv6Bna
9TvLHbWZXxHdu5TsG+tYUGZku5O0lsLWdmk30RLGseHCeaTAsLN98JfgRBDP12ax70bhIVwGRf/W
xfRji33wLo3ZmI5MQyAejmrqGkFGCUsp4x6d3JuPvFfZuuGeeZaR1oMFBpwBLLDZ01MAROarHTk8
zMVfiGMBxMWsH0BkASMY6DXa5ucXXnhEPE+PmCjwqCgYievzcnZFZzr1qgADMfeNQhPDSUdZTycE
Y6HjrM86a4qRLigqMJtWaZNJzccGtRDcxZm4PLJROrJQy6MY4feSVhAJgGSR0NVlNfs3un3UcACN
xKaDr7c8xAS/C4ww8X9dMdlCZM+HFbfXbdFKl89xmLhDuqe5ZJYa3WnmpzebjN0QQM/iNLZc0ZrK
9kI7Ekj5/aYtFQmm3wzelI1WAY3If2FnaoUDzpuJt7KG3D2bORu0X79sqkfsjGerP/8p4voT8xyG
L0l0fB6aZ6v6HLh5EjQGuyLdTR2goYmbOhdwiz1pIrx/AjHZ6JgFGimkHvSfNFUUUbyZC9gKqcJI
pda0vNheoH6cXb8OAIzM/lgJjsV+rBmkDL0jPdya6OvtF8ngNuqQZG4H2enn2XRXnGgMsk7Dow88
lh9QvLJOOA4CSz81r4WnYKd+Stk9NS8jtzOp1ilNYltDIQFRbSL0PzgC9CbH1FHkbymXUFwqWaR9
0CQtljgWAmLiD2gFSGopafW1FDM/pimHlmBUTh5wqSDU6oehp41cy7foxkYmALRsrLIAYSEe9TB/
gz8NybOj8syO4wOzgOc5QNJO0NSTFR2uFTHXJo0HzbhgtIuZErp3s1Rg/5pqTOi20aWXs0NmZMca
8uecyvcb3NOnisrcyXz7VBJk4qWyCm+25icmQ+c7wq+JD03MzI7mr7w//LvmEIw/ell9dopjPLDE
TASwe5LATLll9KtnWgx/t7neOgax8HZM2w4ufJB0w1/sEByevowHyIkJO8Wz43kBCVcjPhFcupT2
E4Ne4AHhDVpbTs3PHCyizx8sLVpdVrPv7o1qM1cZIGxDGyFvLD3GhIcCcRrEUIV8qwVf9fHWZxrU
EvBtBWmkiWNpOBmabASpfNdWoWsiZVJ44sKPP6E46/9irlHr4bHMmIEAAzHlKYPG0U3dGMUPv/dZ
SlVD7R6OWaJ5vExASdzd1DTBJM7siAmSKAaBNxX5iIXc+D8ysLlQAjspn/0UZsseBu2nBBJFd5T9
yLEdjiVHjrWGeavyZKZ8AoBy05Ry0H6aO8QzhJfWhm/d0PvI++nLA289EIxI80rqD1po0eFvFeVV
hmApCFihdZT8ZNlgwQybDJdvtv0PYLJ19VHCGBr2b29Q8izUkW5vmNpkR0YVyDrxY3GySWC6T9G/
XnS+/CkNo8VXLxBLx7FfdGcSHK4NiACCzYUohmOMEvj+GfN65u9tMXsPcN+KoIRbOoe/KYIswyA5
5KYH/U3k6gv4DFY2KvrkCbjS6aii7RypD1yO9pJyio9XNQv0p3Kouo4mSrt0qBNdoHyisBRSJZkR
lAQgcv2V8w/ThXMqcTkqeT1bya8swXJqTxSFAfXRgRRP74eT0CwQ7pX0VzlFb+y/OmiD/nDBQtP8
1fPoLiZ4Tvp1XjqbXmx1OJ41C5R1rzc40wwtYC1VoiyppW48D1a68zsn2ttN/aSqLItn7l0yBBpz
HIwH9yqhGZXDWNGzsfrr2sBnZ2lVPEli9qKXDcB7JnS2zIUWRr7umuNHEZqTILm6GFgT4qgfww36
P1CEW4xmAXR9Tu6FtwDuJe6SNlf7jNX32QMZTseTzggYiM4nr2aiD8h7L44TQuiEbCETizrdFT4R
W6TDabLLJVR54ZxUNZF1jlmozcRaRn58aNqouSI5xP2e11N5cbtJl3Rqsw4+nU6CBlKSa9nCyOK6
BWBJacbkN2uimq8fQvJIYHriusn7ftdxPU+vLuWvfJ5OtRM1vm6y5B/C7X7dM3xstg5YhrwzqiZh
DtPf6+xpDiDF1YZB8QWFNVITVp/UOHn00p04LVhttWuygsC+fbCiPI2Wq0At2A6mjeYAheP1Vc5Y
T7OE4iWzoj1dK3nVXa503sQls/wHZF4qFEKEZGbzWF/LRd1XV//Bk1NRzaU+GmVUygfxcE4tNMRY
iEOYEBG+uawG21EKkMPwp5wDhjGMOWeQXSGjczzC92R1j3KJqwk3Dv/g8oplqdLvnYokicI6NXep
Gz2OtEddkm/uxgu2M4SfNQkkG4kpdwgsOgUU3eVG+fhc1ENhsBnvLfvLKn5SD56XmmC9ozLgERwS
73bx30Ct0OVTVSSoyI9FMNSrQLphMw2z6SuYe8OenOnHf+ioEYGlApYynOy/UUCUQEDlWBGTacGf
D3W8o/yIg9HCoXA7iTkdxdE44UFZ0wicZWgsdwE7F+4E4a8MKuT2FSA2ITyTfeyLrOst+rr6gbXw
F8lEJy72V1+GNhwzACbomPlSjGtOcB3YJNBkkN2CvgKE6pcksdGntjqnurlkvA7L4pVzS+1gmA1n
LVU44LsrXdoirrGXP6Q1GZUKsVvmEuFdd7q229jEKDCXRkfnkDM2TyQyy8r5JBBAnbenz2qvs47e
TqNTvga+OVNepI4u6Ml5sP2ZOQ0tfVYJzjmHX2UfHoQkF4z7/2pat9FphdEmuzxKUCpGI/bk6rCC
4D92gkRLApSiNXa0+ylh8AlGK/kShQqwr0yz8t0NqB2E0MvguAc2n5b8AfmTivtyZR/FDNAnzWUs
te+KEx+vwl3PIq0I1RQUwuAw4s7jI0GlMBH2BUlcXgBj7rFmIXQUoaXN0hSz4dm0Mj4RfYHl0BIG
7VXz0i629XzZuMHmOas1uyl5aREJoo1HgMI511IkhcGUdUOamt3+spgHaA5NCnjIHaoUawBxeZUA
BXsxmRJ9Or/ZyB8AR7xZUcBWUH7rcve+wy3DlClLKYTJyAXItggxoru5aaq7MvE8875vmIw5P0Wv
55r2qy9PYJSLuiIa0JmQELpOQUO6uuFS+RLNrSKMitom2bKcG5FQyCoJUpjG8wle/87XJ5h714/N
yCitaWFKXtywOQ05YGbT7IC+EIAzuszj87Xf+iPjGH+JtP+OVs8VEA10OIvic/x/ZzUyFAJebUTf
iu4sxIAnY7LxghFKgCaDDNf8AyFatYtf+vHi5HXLn1YAzJSyCUjSs2e5PbZUEyA1OJe5tdvzIZe8
1q+cwU3RIDhzvKvGla3fOusxgtDgfWoJ7N17xmmcf7iXJdDmqI/RkSYlKEoKqEtqwtdzhrrke2By
WzxKHzNyB2BnSd2dfQM6LcpPZ53Jv66Fe3PZpSicjI7wZ1YbbAnxCX69uc9d+nOBLzExppGLyKa8
pOsqdK84nTAsFnSItPHvbWldwIxPsFvdmXqTRwSbAH3rnsbZD9ss7TO3ZlaU1x57meik4CKBxZvM
I64TqJUYhwg+DgThaVcJs5Q1cR19fKgVt9HwQJsG2QY17T3jpQT2zm1AhhAMJD0AjH2hAOSnvYVz
cdcKILHSHwrD5yTopX349gRMgtwvrLgNK6F+cqeD+4XxheRtfV+7ENVHxMh7ysiEZpPiqFoKidBD
WJgIIoUP3bIG0xtw4hRMZzv9TIYwKAdzenwDMVB9Qyef1EeDF+myExXxV8crON6vn1XUWz0e6yeS
PLi+reioXZSSeeolubiFQJqET3b8dUQdhTc+xGlyfaKgsKMSS1KMXO1r85UGGBvght7FR/93tWkG
g5fjD0ob+ErnrGPsKbwRz9Cv5biqlv7SNcVctrwE+EiXO56J9TZ6ZkiPB36ybxLm4XQCFXfrsZ4L
JRV+P7GVIn6RYOklZn7LvUIeWkfLlxIlQ7uM2BQPFlB2Y0IUWkX8U8eGCs9taAb5n2EnCUxaHQNm
7RgrfXJ7bsulPkM8fiHef5OCMXB0OHBl4QJeCjj7Za7kjxhfRrRRcO/0w5xf5kzJaRYD5R2mJh15
oonDTuyHD5nmqPRuvKBt50KbiFdLAbhoylgPOT86qNLFShBLx8V9m3z7pfY1oS3g+gAjy0z07aFe
o6BpfUwf1cxmza+3pwo3ecAPF0za1kSayfZzkO/IhvoxMeY8K+CUaMbt/0+VAd7p3r+f8Fi0eEOX
aTa66tm4soWbaXJLqXX0qmlRKwWlmHcsizKqdMvL9mBC7RJEIe0Z3kksckDXp17U8mpIDVnHMsHv
mhqbHBArX8vhOA7w+5CTtIJc37u8MsvCQWHJcmKkxe13Y8tzSp/Ne89y5MbJV40tmKWwXIiiVk9d
YQzb2OYO2ixt467jvG4NMmZ3gWEsrlM7cWxKLbMfl9tmv3xIDH3lnd5ZZWWPaL2UORdHykgpSZD0
sFLCY30UI4d7/V3vckBx8H5XdGuXQs9hia51w0nuh5q38cPcclI5EzYmDqXpBkZpWGFssjYSk0dc
642DIKctwo7sdNPs36F4za4MfmDRVkYAGJCFdQNtvFNLmwt5FqY8C7VFGTTdcCa9VVm47kAOhJ5o
AbAamXokvrPOUgoTz0tfnPWdp3RWymC0X6td9S7qzFWuhg46jyD+YDkP58gTWUY/C8c/vn4Ah4Ne
NU8lhc1oDTsHnEpAJ/+zvvJacwLCSs6rl02ffSSPtDbNwly+Rc4rekZ7CszoFj+mltjutmn3NajE
Fttg41Syt3HTr7dEYwbXYBnVRQXbQDXCp3efy6LprQ2F0XXEFMgXZhDch645sjCQa4bPlJLQg9sU
OJGkvkm38WGiRDVYSL5xbOb0W16UFhLJyqwDnP4PbZpHeDDCr94NnT0hUJWIBVCvQNmiWSBqOoKZ
h7Azq4cJLboBiI6FKa16mN8B6esBA2RVpEN8pRTsvc9UUxOyToov7dux21NOoOT7bGqNJG8iu9Oy
iVVNev3K/9Ku//REC6UqCtKswMemXo4m5ni3AjCddMzZfXlkPTr9zUIj77EIrpQPukFPOkJlpuxj
a5PlaEuEUguFBSfj/6lVuEjgVOwMcJU3ADOaPSUYq3FupoxEuJmwmHXIesgl2vQTc1EztIpRNeLa
CN7xDHCSfGoTYZVuFpzyYit+/3AB7GItGVo4AGkhm5wRaYsxI4b3LRlBkTicPTH2j03wjfm8JPPg
udYV2h+DBFJ6CT9fjor0YdEoIaLgDmDn/d1eezFHwFvbky0myzOn/vsXp6p/YDcnPby1nk60XemH
G1Oax/u+NB4wE8iBw2B7xJsL78aPjkTOJHvDGfyDq+uBZDa3Hfh694VJjRIjr+vNtTsl6PCJTceu
P+l1ZfAuxmGff8cDwGJO+03cAdV75DQACPkNgdKRnHcBnWVrU+12qS7t8l4b+a3O1w0qNPJanKFH
r/I4e0m3iXVxCLq8VBRp/Ll0cQJJYrODeJgaCZ8rN5nDppkwNB5urz0Znxv5DE9kUWvcPAmLnana
RzJX8AeVtPHv9K0+cBQAwYYb3bEMpDtNbb+kA/2ZtneDaumTyf1xdXz5/gNWS77ozR9DvX5xelrx
Ualha80RT5A2GApWOTH64q7ElwgWz287Zwl+/1pgDWjywdOKZJZ0HWiygHztzE+X2XbYhVudFsS9
xW+z/CxFvwTBrWuB6PBWKzVdY1Zf9sGsI/PuavJmfa+Xx48lFwsurq+ts9vVyLy+02zTMVFNPj7B
KFY0iUEMHZtLaDEuXsliVBqMS1xwI0AzMU+QpbBdC5eOg6kagcu5hh9gbyYnpMBKv3efoPcv6Bm5
hk4qChwudhV3v0vhhmTkPZJTLAYNhsw/TMfSWb16RLjTSNpvHG9eUtp+njWWILo9EzGGQllBmZsR
WYIVM2tk0jT/oE4oioxE0LlRHC26CGniuQPYHHXbizU8y4oxWM9eyPKC485F6+vhdBnQAvs/k+6Q
FlUN3cf9il+q6CqlfHJPKOHuj8BDEX1pOtuLQqnS0kuRimgpEw4LHicAAlLwfIuRedf6gM0XUUxy
ZhWAwaPINdSZ7pf6weni7mDPExT+7OxeSFXDnEOcx8g2HsMrLdnMsfuN1Xv9tBCujy2L4iwgO3e4
F5YeP+E2k3Mn9nqrhIpbFbFEExrX1fsmSa+Ou9D017/k7rvFQMRPoPdULjcIkAi0cK1avxUl1rhT
C5cKTi1kdYMtLUjWjgsRwGYiHZaqN7UvI/VNujjTpk4BPCge0u1BVBvZYy3yVmBqkqoMuFX1ctU6
SCTHBRsqGanIL6X6ZOPD2Cx3KmeCAAzr/8v3rg4lcT8J7U9ryTfVYkA2uIj1vzam5VNc/bK7UlKY
TLnG/WUE8PfVhXxHwJbudHNuPfeBdEOEYE8jIu9/Iv+Pkx4xJ+EvI6JTugPIGApXrlEh2z8SjuVs
uYgURR2HXylzduyuP3dMdQJ1fD1anrwn+IJ8aCUbjHPdOS19vYEPvrnmGnxz4Qv+g2AyhqCrsb+Q
1RoB9ORSdNPvM5BE/vOU6GNQ3CCUWwPmxGu1sR2HurpSW1VDEvbJA4pu5Vct85zj+bowl2oa1bcw
kDCmsn40JqBGNw5ckeXhuZGoueQtWJ4VWUBIrUpIxSPhzviiMKeAmzr09KsBGrrxRAzgKzf00po5
R489jFILapkONytVKEddZpaFmvVsiaeMJv3E/BgNcBd3Lr3h4uD+dDi7cok0vNDus0fqi4w1DwOb
+/IB5MdDYQ0LRx1t7sESa5nHCbuW472PVD4wIdTVgnQD+Is4TyCPOOgR409qu96F1EVPFit42fgU
vPWFwLc6Xt3EHT8uYiD2XwT5eXhcOr4wLCTv5CovFkqVS6AfwL66PWVPAjxsgBUj/XKLBDQRvNBH
U35upeej56nlFDLArL5Yqe484gnSJZXzmePdIgXmcA+6r62nZ2pf5KJlnVTDJmx0YEHxomd6B7NX
KQHjAob5icwO2Q0u8yE9XYRvDZgXq7RCnZj4ygr6QwwgUHvV4o12Vng1HZjl5Z3ncwGe9WrUzJBd
NwYXoi6KjdVoayjHpRGGj06aV5fM9pA8wywODcTwrI7XzEGt0bFCsDOo2+Vqvmgkbh3VJzZdXWgh
acLIsgb4Q96eV5TNBmh8A1pbZ+bc9xyFLlVxQy+eKOOK7x8gx9t4YActPS0vrjQVF9sUE6SSYetP
xd9V1BQVRjNDEZQ/F8Y79aJ3cq+7iE1s5XWExZq9J78XPS1LnkIf+hw1nslLbmugPxnFJT2zz6bZ
pO2NunLn5DdLHssqd621eqj/983W9qV1WM8M/s97M0YEobnYunHaOb2+PPLpkE7AIW+8CvJzA0UD
GEB9J7F3JxXIvhGOhY+VqwrY9LOPTkhnwwpoit9ap7pSbk4QejK9EInl1eFrquKqyP//T/a3snjb
0uA0pcPIKXPdW43qbT+MH706HUB4kopiREX0nwL9VfSX8qadHFW1lUujclTDFN5kuJT+Qk8L6jk4
lvp2R+7RcUf1hD96VJN2ll6nltBA+maBTLSVtbpdz/O3cK4DR1AC+f79tuEvlW7TohdsVnpyW3xK
cpnz+M9IvO+1X+8J1gKXbgPuraI2SBXiTLGsNMwrDxLzWpdGzEh+6EKKsUUr76COFV9Zl+Eh34fN
vxa2BD7rIuX1ThsvvAjtqtFaiHMw6SvJljQJPCjAqDkTCX6z/b8kEz02Xbd1e90T0Ddrgf6+/vgV
3rfXo21u4F/WfyM8qaVtky9XwfF205tg3Z2Gf4AgoshKTcZ28180Fs5UV3gUTLO59i5h0fNSz80a
ffYp7AGoCY0GIiyBRHcUCqykU92NCQXGFgdJDFki6JUa04jmldVi7yt8mHZuNLN4of+dFpxpiPjR
xCzCQwyPmcHrU8ttlbWFBp/u6dkEnn1Uo7leHNJrL/PICcD8c1gGx3cCnS7EdlZIioBaK+t8uJ+B
Pd5wwkqux/CNNV66DXOdAmQ0biPDTxa8t510b33OmLuR5Mu0iHQMmGcoPuPS/sG9HAI+uBsBu4P8
tLX6wKuxWWj+JxKx33opaegStOWeGFhaPZ0nP53B5WHGVKcO1Xj58XjEavnRZkIJXHkFa2W1HM66
wzpjBhsxQtrfA8poO3VUqEoTq0IGL0UVHaS0iPgl0aR3TEbYhEvqS6zjyal2m08spGDML+aLhOlh
peLolN5LVGpLDRk5jUE9V0DQQ6FwfbJnuRZVNzCMauQwKmHGxZTbwbKfJ9V4X3/AqxWWC1UVBeAQ
6pqecEK0XyCSS0O9ymPD01N3mh44cC+xO/JBly+2p3/1dpjfUHPjNutymAByABVNWIDugTlpwMwi
KrhnsfXMHHUYxd+jKrCvx89bT8XGQ2gG+ZGTuGwzFUifioC5MNTZRD7NVMZBPVUV9GNklUZILvCv
1T10pL9zDKfVFRA961mVQ1ahZ0LbTz5TFrA1jb6Ssgi+3M8Rs02LuerGmRRbuxhB8sNfstxQQ43Y
9m9MXXqa5eAyNu332bjoAlxAAmJh6MB19QgO2mSY4JjKikpd460gp6Y079SUrmMm0GrIkeqgc19B
5/irXuNc6bSx9hf55urlVcUj5e78blcvr3oFB8SYUOaXDXv/ZRMyw3eIgQJK8/D2uI3gXq+sKVao
MVaecqbHQutYbGPUFBfxROJy0g0iVsRhYeln2fJdeQSC9wa8VpiDzpOgFms07RukzlsX5VHP9ILf
8zSdQeY+lO9wNmNk74YuKThX7Q2JN/T2sMYfZ6mnJgSOytbR+f95A9MQt9wDuv1x8a/YkLrRVkzE
z63n9yFZdfrwaJc7pZoOjx1LWRul4cT0KWad59n97qfjUtyrs9JGVCywOZT4PZevgXMGTix5b2wZ
fgvcti0p7Ms2rjawoLeJ4ptVIKv2WN3gG0Y45z0gLg+kFtZCrHS6g0o9eWAmqrn7eSbahPJlHmdS
N87Oa6ft4HkB05NtJaJh44o/DfafwPE8ai9mnBzEus4v2bM/xyY6tox90HYryJE5BaXi5SRA71v5
0AEgct3TkANmKVFbKKQobcjAy6/gt+oxB+BLp5EraF0zEBgeQH7KpIn5L3XMAEeqqvS4mEA0K2o+
wcDSudO2ttZw5+r5WbZ0Uh+5vaTLuhR4cJYL+rs1zCqPeUFhqD6P7RCSyl8IMWH8UUAn5MTPQZNQ
NjW9zfpVR9oBYvtModCkDtWY+lFL2LNg/cfwihUsiFT6sZXDMSeLWWBbG6f3HWEJ6LmBSpg+AixP
lnbYuuHqxw1jewQ0eQUO3OiQdTNoHQ2gMv6alxWK2WKcVtIjBDTi1ZKQLwxDCTgn6AGlft8z2KLh
xBg8nDG0ws4W5bjJ6wtnSVKwuvW6MzV4pamHJz2MLzHR+XGpP+J1A39KWTMIk+zmFPQeqxePoZF3
ymd+jOL3t3LfC2Niq4ZnW01R5NTygxNyx9f2gMIpGaVbN4mz5KCRAfWcMDvw38TJ8yiqxlp4usZW
ifgTGKmW4O2DLXHMBw+0OZHlL9s0FlM7fQQK87Hz81XcaSoYNpesZEw0MJtz/9xO6NQda3CdZhMR
RhBs3pyYcjHHv14Dg4QVFVXAvuMvUl84rW2Yc9g6oeFOVr6oxwxMKQOGHcwFqEteAVcL63tYpGxw
jkqRjiNuzVwduWK9GSxj+ZM2YprLX//F2f8+2cb83owzqO4XXjQTybZqmjpQqqsWsRG1crfhSfPd
NH+EbXCELt4vq6/nUebRbgrwMylwi4JbsLUV7DkrMMzihn240tTywvGCt62UQmwAtGI61eXi1ayg
cWbuJzv78xImen/nszPrj2fWvey/JZty27ijHUKkJkF0EQls1Y7hm31lhXGqMs5jJlkmpBEOOkRK
L/rb72PwBLqQXXlycPdV9rw0J9fjsdiZMhaccEIo/GakvlfY25c0nU/Xwqh7b5lAf/g+A85gO88I
M7n9P4yilYOfB4zvCenKwpo8TgSWf+oo4ZunfyEEDbg0oI9jUBaiJof+b7yGw0EfFvIKLIyMJ6+B
VUtwl2SgKrdZUtNPGI1/LSp7pCos1QN3lRciwseXxHXegHlU8jhU1wp565HPRRFBj6kIfz/Bt4eb
fAMoKlZPQbhsbsfK7fauAK5V6vnDzc4Qbh2owslpXKXniNLf4Bho8JWSCwkWCIrA8Yri8VCDTudk
hMl3E+uH5Tn49XetXvENT/wi5W78214r6z/HLMQxLgejb7iMkmwHYY+TSgoHnArXXdRZa0SbauF3
yIrrxM2943EEun0G45kMJnsItPBpfKnepCYm8QyrBhOeronwOQfDpxCfBRZfLt3BjD7/+8nuhyR/
Z/gvqqqv7GTcGSvQlvRKyhkl4wM6zrZToMxUCe/Vl9GDmf+YMzrurpRMErsJAFUVT58OQ3m6KWXV
EsYNnzqZBDrsaCX7K8wEqRmUa+UDkcLEbdP7+ox7yfhEjgmYp5aWE1j7xbiCOoPxHg8L9NcHp8dP
3n4EZTCJC/0kWD2eIcHrFpg1ObTqSr2XyGgq9ZFtFLYFYTUx1vMcplcSAoA4Do91YE3CxC/w7gZ/
rq19wj1g5bSufC49uhl+30SY3R9tKvn4eVGLFqDckczvPwV8zu9mNWo/AKEJf72itXffRUlMErue
y9blICJEuwFAnNAvQiuxB5845+Cnga3PuIDJihuejSCdbQwMgpq4WHxR817QsWX8Hs8WtqRLT5/U
Hs5kjtkV9CmoH1xZAxkwCBt3ALIhktx1zpS7I0/9/X2nJnJ3J9ACR0PK4HYR6L5A6BvYDZAA9EYN
PtTeowhY7sqAjjn/2Y2RfSLHRIVlfyVUYF1FUIE54mcEcEP+WueTCeHjInYobsZE+2th0c9cpYgs
9+k7XAmByH/WqJJj22NG4IUJTtksj4EiKqkUZnrcgBFbP7Sh1EJhrdRryaE7erKPXTgepqCmoboZ
CHPwO4VrWpa7JFsAiAILx7Qhg5481Z2JINBPiKLUyon4Q92RJxUcCxfoW5tL7NAJTzLgrtTNyCkL
P4t78x0G4rm15SLX1uv/gPy4D/FLZrG8yyj+FrcF/j9cnxfhn5N4LOXrEOzzNyNR85s9ccgepW1A
p2nura5xB6sfzrT6J864thi43sytR2XcqsjBEv9fQbn6VcMFJYMA8tnXjv70IO7oFXqbGpLzm+qT
eq0xFLS61OKNqP4jKmyZDMEQ/RO+lprExcClIayGa4S55N7sDIn+f6p6NqSRHhyZUqfss+HSH9HN
11eYcqUbTwBJyRl21/hYEJCJCw8nxo5+QTtNruDRXelnPWHqr5hs0LUC0QUVpucf1RjdccdQ+8gm
KkQwuaq6Zt/fvbS9gn3+uEVxBgqFGoAHzi99fWieTbqYOD79l9T44Ka+bnC5n2LJWtC13bIMh9/A
DznqrYkpN4srzSm8TP2VURPUnIa5Z8aHA9YJIT3gNHvNC1yvfOvV9706sn5FkqxEoiwSGmve2q4x
MT9zOlYzcHtL4dROHssCabOkFnxySduFJ/MXPltzWFEaURK4PRrX0fYrrAM7WpkPP7iEIrW3qbAu
stxhoNsu5TXzNhlGPW3rBA/UX53JTGN+xjp2zKk7PCIlY3yee5sp2j9Hua/3jiC4xIPz+/1FH2yc
/vfzC6n05EhHQ+5XYscaxugto7N/zW+PKjuDGR75ailWrs4abnuJg9uNOBUJmXPInvgXBBYKHoI/
qAFcrc8iZmlN7UVplQeH9O9vEoRyA3FCmLYO0G7EK9Oa72JbC5mI51UkAPk/uL13Rry9YanJjocg
SeW1YeHfOFMivJ+GxOw5XdLUjNhzvZKC2voGvJE/s2CMOpUHN4UuTvtWO8GuClKTlk93m8cru9fF
tvh6FxAWKzsIcQGKLm22wEntGKm9v7tBtwYXgmq9cGrnA8aJsk/ueD/b8pNkx761iq44215+0wX9
mjFjK83qvbFm7YjPBPx0PspVN1d9p4DN4XYmYDRYVhmzcXI1avSS9ZztgotMXNNgyYzh0UfBJEwm
5A+32CtTyfzuPTSbhK7hq3c+1EQmlg96xSostm9jkCJcd86BbOFyVwGIXgFN362lZfSFLGmXqoBv
pezMrxsOzn3Vz6UUcV321ao0Kef22gKW0x9QORzk8fUJU4Tq9Bcd47aZTpii0QAwvLmlU6G9Ao5s
tQbXy+vSHm9RfvKA+A3CFcxV0l/1KeBB7d5brzWI3//EAwKqVMJZQN/eFqWodrmnyWuyp5bM/zI/
Vr/IOJ7X6lQ88CBIcVAdCqMxTPlsN/h2zuAGtsATsXK2wgDyFqyzpnGmIdBH1NZQZTWa/ZFx315d
JUvXd3ynq/uNIUGNhBQUjHfZrvx0RDpU19yCwDnX+za9GyT4PzUsdFGY017ZrfnIXRE4YvJc5K4R
HHo0BXioCwrep6iGCC0fKc0OMK+qAGcreHV8PyZtefchzsckI4Q6TulZEWWvwvsO+qkWBz42ZjJU
3aeqDIRsbxX9Gm6KHbjenRS4ARK34JqdobYBPTYITqP56VzDEeg93OjRCm6n4n0Qh3l7SG/Pl5zO
qFW+BI/mP2EzYhqC6fUsxSj1XLs1M9QlqJ86emmXvBFrIjKTD6r+gh64abFlEqp/fWztWAKA50Z8
juAedufJ3T6JJ+XdW9RMSbraUyuiAinGfDPZqN6CAPOBnpKAOQ2z5GLpxaieXpDKogioCh1iWqUq
R0i8pIDhRKHQxC+8zVhogasYM/1tyHJOdN1lN2o3jfrow0lKamU+Y/ViwdPb7wuyyloZbq3b8Grc
iMLSR5r2Wd0/g8FwTnLMCPzUjP4WQpi/t2Dxvxr+cQs5xh/LwDm5IK0Iw8ZS9Ze19bnwILCH2tbj
chkTNnh8BPDvIhuaDxtEahaS3kwXQ3SVv+fh2XMFB48zVg5zfBYM8IjOgMw7UIQq+GzqaEPIaAQE
bqACuwDHcV2uSqUathnZFFuOy2ZQfulYdLqerRVo2swZ+aNlqw4bnu8Ku3wgm01xtInH6xGXLP6+
Xhya1nNwquzezY4MXT/QezNhNS8c1o0TYLDViNQzSfFsKGpxilvLZZXewOFQw3xzu0wdaIQHh88d
msxOdf0+N0GbZ7Lxidgi9Imqs9kEKLIWbuQezja8A7RlVkH736JFg6cBK9j12cnPLZIR5j3+0IMm
VYqi+1Ui+tBUrZGNspEiPKCQuZgrVlVHGAR+MOPYimfwuMGRPioUOjmA9hdrYtC5lYua36arNCQz
wlzLHP5I6BAvhplGtP9nREIJGc8memS20Td2lC2CW5Nit9Ryi3Erli54WzIdwUO4yNJR6rjBqi2e
uTKPZFZAaJjYVCOfUvsdu69o6VRXOnI5Ypm9UeYrVvD1Cz7t2YxOSQqPdvdrj8Bx+4KQxdi+qxOF
3nwgpZF4i2xvYmdGg96wMQoW95LCXVbypPADOz3Nt6fZo6Kapup8powELhW0zb1UBVVXirTCevsu
hubJ0F3WL2QO+5K8Z9YK3O/qlFaecABBxBddiAaBv71Y+hqbqyXJc8kXyIVHwGYE9oF7vUSUXbBd
W8JZ+Z9JoyshZvryVSJi6vmgYDsRQwHuZuGHGfgLvAdJVJDBAIg44nHdDt4z/B2HaTBgOycRyXji
QM+Pki2ZqO2AKy8lqokG6zlC7jtf5ziZ/07utZovQ1YkJYjo+NX2+XBXUO7si4Qcte7fsv/PTOvd
bnKA2AWS0c3Zy6xwHsLzLJKA24JmoVvEqaQysAmi0712oL8gVkhgL5MpWmQcMqkKErH/1g9ZXZO5
m0X4tDufcpOD9v2OkwZ90oZ7IfLzx5hX1ds+VAsERLa/V1u7A2dpgckRVkXh8TWDFLlB0PCOc8KI
Kebx43Xt4mVgh/E/e+7oChLbnZY9eWew9rgduBl+a2+Nuq+qnIR/+VxEhz2gl2Krke1vtWtuxYEz
/B57DkwEbHMvFbmPlTy4vtz9ynQMS0xgrn7FOH0+M36R7Ztbov3XP1boNwiWwN+a58CwLyGP+NxV
s8WYmJSN9ONKvCf1K73h/YxdAe3kYnboD+/E/441LAUqk+4D+TVLZ1BoTalC1JA7MZ40ri1cedDm
dNQEQ5d1wbxskCWPW5/p2QPLgcKAQnUofdPce5KNa16+hFNb574bzLt6vmRX3+Mx72R/VJsZPNWh
GlGRi0h7y9raXkZiGMr+5HACIAGXF4iHN/FoCdDuuOIiQFJUzCfU9iUYde+mZJ5fPyHP8fvh059b
+03I5zqpgcazTg1z62GxlLEqMUmxmnfMheMfQQooKE3eysnoEyRC+Wpu7vX6b3olJKC1SGXCeeas
yEc1Fz9ZPWUUyuebnzJINkoCwf7yat/KoRPcQ8WootNX2zJ6ehjoNdw9U1wf4SjgsWgwxG6Lhiuy
iScxXahcs3dU/MJowrohs/h7IXB19tEct0EvGj+IRUGs7aBwIdUTJ29Es0KHcIjovQTH1QTiIjbN
jtlGrmY/DH9jlQUtaDkuFSPCWBQLmzEy8TNsggAbF7/avoos3nnIkF95drGGeP0deUwd8Bbk3ol4
lbNt0khjUY5yW0ffU48fiOjKqpHca3VTnHyGCwHy5Cq93yz2v9HlqXsOwo0uWihhBGM7xf7y9+8Q
Xt6prNeZV+IYPK+H1Pd77rp6BHAN5wT4jtVVuV2qvY3xEPqAQPa2vYC4IgISNwbejd+bkZtkbn7Z
DBUGV303pjbVdLvPsBsTqbO8Q0+/o2rm+ZvG+UDfoWO6mku4QpkLroYjyB6kMkztufJrN997IroH
avJc2fBbC4s++SJr/Y5rgsHcwk4sM36r5jvU75nw+M6KnBq+IgPw9vHm1S63RYeEXcU+vYRQIdGy
07R3xO3W8xKc31mXstlZ+hsqpHiuapCHxH3+4cro0eKEa7XFIc4Kmwwn2cnl7mp2KReKIJ2JfmPU
9LyIitMvyk31Tsm6mSOma/mwroHFd+x4eB9wnneYw5QG+/tjbbEiD2VsEvtDgyuu0cNQEn7GQ6Fs
G/FnpnVmMdhi+NV5NsBpORabmHtCW/DB3XADkz2l/1cUjRON9cORs5WeOu/STyuelZup/LeVmzuT
xW4N/AqSh49rE0OFQC7LbttIb+rdzFVWpN4krvbvtKPCEjo1WH9UGzrQNKbIgC4Mk5TwXZHY3T60
WEEanle2/xVqzUl+gGMbVtqKocO4wEK7jnIA1DzEOmZceugCYZ9LHoo0ZlRAeFelCdGdknWvugXP
KuRYewoxaXEGyOpUPCMC+igGPX5EudvulznoNFPqJBzAUd2qQJGcTxJuEGI04+4FEhZgzd5BGRBm
ipdjrvhTTI5iOPjtIAPSTlNkuDpdBjMUbzCi0yhQp5b8VdA5DDkTC3hgqpny0JlpCyx9eqKuLxeZ
Fa6FQzScaFoxMR2mDhnQ7Z8Gv0PyplsAkop3GJrF7e8Hk4WN33/SSuDsjjTL7ue5AF2GqeCsFUfZ
Dhwo6PI1lDeZ3U7Zs+MkXRrRKaUQGTIoSPCfFvbZWLSEFu9VkM5WfAcwbxBWxbHZyT3VSzV5/PyY
4xPciLnK6tZReNgvny9Jb3GCYG0XMlUL4xy704hdn9n3Xht2yISaBK0FMjCEGaKa2lj0grl6bwPX
LpxPYZCrUTywt2PimEGUT98L/P7SdM6hyIzmbn2njjXtIQ9ZT3M5arkSjitn1m77l0dlJqTY0U4Z
Ynu1UjnfKJIYupbkvtNabZQFOVya+v/zy9a35lycs+4JWkXrFK5vQ0jFccQ5CjJMhfMK0rWhqHIO
m/kqApUzdSGmrP60sLlHCtxZv69qsAtQhDwE5tGHbWMCdK8l+GBlkXzWI2pwC+6S0HwLeVGp15KA
g6VAPVdmLE5NkC3r7uarWhXRDF6lbxZMsb/NqW14BbameCiWCIRqJXptrZgTnY8dztFcjNk9Tt7B
pvrF65x3vyNw596h9PhounsIHFMQdMcjxEcYssGjOWKtRKPMlIjIrnJSN1hbOxyqTw3TXcvObWrl
xWMckEGOjbQY//I7jAwqi3/70r98m4ehcg085TKMkkzswZGjwh3AiEI3PNY9nMfNW7nUQyfWJGjE
I6d4ZydzD0XX9/DrWmUlCLuiyFalRpib3ZCL9d6YP9GF208hXlrlYkuh1wRTFeWmoSl5phtGklbT
2updOoeCWR3KVwlEgYryAHC46oLQHXLNG5rBlqThz3nyV9xDKHje9tIYULqVLGyCeoU70XqkGfkm
cyUXAeB1EWNwpL1iwWMZVOnBQmQb4BwyRUlDcicK1I+al7dtJYpibp5Q1eCkcHXXtN8MA8x6cLao
tRYlAkBc9zxvzQCzTadBh9TXG5s7vAFUeqghRU5mmJB1eD9Gq3Rsg8iPjfmaN8GQ5ErpVxptWZ4V
mSEsruPSgAimALrP/NSfjvwuw+eSgFbAfiTZbxq0bYrPBcQQ5inPslFR+Z0ltM6X7Oo2PaiSie4i
1J0KN1JqFgl9M3atVVidri3SKP901qeZ6byeihzyW4E+wE5BFpBSV9+i1F7OBh4iZ5ZIQaZjF9Mg
3wmGBmdWvCpG9A9NQieLpVTB28wCyLOihWEDDiZCQOPGs8hU3DXXFOrIOoguEuVNljkTFbvPTkbU
rlatsJAaPq+r2982i0bB6yjGv/Q2R4cnnTk7LCIHXoveDxDuprqSlVF7FQZ9rolA1/WzEB037xwE
aNdKxL3kAVVDqfdCCVoOUe2gcRAauLYlA2tfXsCDV7p5K4mCRyWghK8kNv28yTX4OmkMgX6hZHOa
QM19LoEbEbvBYZcUAohg9+MabxDxox3D9QxaCMBFV3UijUzpZ6z9kewjfPQED/ZVqDTu86Txsnv1
JAztRFB4vVZFtMrY47O9wwkWV6a3cmnffU44iOXl92bKbdPJHUfEfbRG4Vx0i7bodo1K/cmP7T6U
9/GDuZghE907PG/LCMlN10OmLAVjRJw/srN7Pso8r0h3bKVo3vK/BqdZFUQgcAjdlN2EM9DZ3cux
9Z9rH3klNb0E+k0xYawKECvF9HpZ2UhWNugScaZANaoqkcmW8Cg6mtR4cLpLmgjZibh4kHLWZFAM
9QKE8J95QuOVaVgElvZu5dQtG+XWs4T0/bS6614tzuHz9LVLy+InYb0j++bn8Phs/VcZrxTuk3cC
Z3BIY18qelCMzPyuEkPWu8G0fMJhwKNFnlv/j/cuLz9MBF7AQi9LFwguEUR8U41OwxxKjxup6bqi
I9yxPIN3Spc6E/dKEmsCtIE6oHG7jgl8BaWVWac0CTOl6cUYTs81tXAsb4Mp48IS0B8/G91LOw/F
y52k/Gph25ohpepCW9P8lZ0bBgWxHvWztHAolBzbc+6nDORXQouuetCl0Qy8Z4HEjJaBs4cONiUM
TWDlih6FSpM2XyQw7gn4gghsiFExD4sKZor2VCtNLlykrZzQATTfkaIedJ9fYuh7ke3PWMiV1s7E
F/87GrHZtxapSoGckWi01Xp4IYYm8recPOPGCNg6jWKe12U1DbnPI/NHj0naXD2M0rn9S5e2FoPh
1h8hcBsj5R9h30xgWrH57nu+9o44ZB+RwbkzAhmLd/+x6qJcQjM6bwZk1invz8kbq+DTaQRyK3Vs
VDf8MlmEVo2uAFkF6LSK3tkeN6a27+4tR9YYNw2IvkwJZgzVWV2i82EpPo1WyV19eh6D+E0bOZwJ
Iv6+GeCcCMOQX38j/KUozN38s9wrK/+2AdIAZN46ocYY5M8nE0OzkjtC7iIn5nNCFZt0XVmsYbwx
z70Vhl46u1F1NpdhPGGXFPa86GU3frrRvSGFWOZiPIAjeGy/vQaUdyllUJQ80bopxvwlgQLHF3z2
CfkPFsBBrpk9naivhSL15SI52fsGrT/ULqb5xXb68pGfrcM0JegCgXJ7JPOMuraXNzosIjx321R0
2R2IwJG4R4TuoqbYe+6+s8XtM0NYtzly8J6mHnuSUz7ti1iv+qoRIHsGhcCXT3Et2RQZCATtivz3
3BBt4ebk5tdV5toArRPYQXliwb5eXWxNQLkHZa5egCQq57YUG6hsJlwlGJO8eZvLkN/5I+qry2N3
CQHIkeZ0xOJiFrXJrsD3XDqEncv3kp4KqnB3iYAhMuYypyuletDudR0cqxsliXoZt/nINDOj8Abb
juEamsnpEiu/XJmMkIH+3e5W61l/sDOXgJhd4tRmZvuSX4VSOwz/kqxbdHlKIJmrJcM/8hV0L30g
zmPVop2ebG5vrVGlL0XijsSJ7ZFVUEa6xxK9pCHvq60VqOmxcVmQ4Y8kbPHf7FKDDD2nVeHfHfWe
F+KT1pUzD0tdnMySxh83RZWtKnOC+dec+hw9gvpUfHACx+GKdZd3C9gzx4cs1O+n1z8teruB+VTU
4i21d2pkXbElbWzDojC3p4kQHUgnFfnVVFycrAkie0ctVJJE0E0IGrR9bMz+UYiPIarBFcHEXqah
hqSYZ95O1D0YUnA6ETva27OJJtHzZ/DVR2epCn+LbcRn8gIaIgVyXmxMrid5uFTV3mn3qZUnJFc2
ZdWeE/RKqkY6EP7q9KxOsT9gCQoD4TTDe65iQTpNED405hgRe4n07igSs4gShy4mwZpkNIqrIXql
rjG9s4E5hfO56wr0473sukxLmEUd5aWgmJdN1myGsI9zbkKTzrfOiYatYu7MaOjbUcY+g8YVl3fs
wCFUB6HfqpkC13c0kXuI5jFbc9En+xwA83+KpoywQuXu25vNtO/JchjPx3NIvXY5b0RhqD2FYuzP
AYAdEBQBvCMrGGg5Xb9zRvgzlrihd1K9BGTxcjTLGeRIhTyOWQdJNLSGDN0XOoY7syoqzYDqfObm
dVNcxwWxm5yrAKhT1VBU613ZiItPXvYUaJYF8whv+LEn87mjRtACe5bNwTtqVgKKZ4J8YyMKCqyj
pIOAkhNb7EU+12OFLMqxCyNTNbV1NYCVUZlTI7J2MWcEQZrngE1AHEc+t8bVIAH+mE72/BgdBr6a
mXiGowZQnw3l8cGHKhqWT806k63YFUfkQNoJBrQftQElkf6U1RV0UntDaz0mFVrcjmhM3bkBawki
9PX0RVvibLKsgcJ1sG4yxPhtxcXdn+P2ffZf8v1BAdG9mQzTYf2K/kiCsynEvb1cSiMcM7hzM9wU
6NJ87xvjVV6Z9upWbxVHAxU2VmHGqKDhCAly5qj3Ztaoz9gnKmwIvXUGf0+q/8MasbZt6ec+P39B
k1zm2GvBEeOuXu+YtULGoJ5YIWQLaWtq3NssWw040dk5+VZrsypcSUk+4EHUWYi79olBLGZmvTN1
I4YtULBktA7dZv9g2njRV/S4nEVjnZaKo6N/Ejk36J62PPg7mnGRui7AEKTBS+Dc8A0O+4EgTvge
UAfksUls3M4WycUSJlzymonhaZxLemyNoFXLL1K6SbL2UUiViIMDX34GF2Wf4h4NSv0EOVsvw1V2
TtqLzhSHNc8c5K1xtPlU5iXBoRTglgVT+sy493iXgQvMpJXhATIc7r0LZvdZkoAJltV/wdhF9Gl7
d8OPYUFHgArPa+dkvPAaKrcINPaLYYS/6CyB0KtYAxyAaUTQOk8T1JnirM1EKNxV9qG3APEv0cxj
gIclkMwsoxyS5q9/kUYG3fKq+IWpV275HFRGImZAe4d7JFP9iIE/0BKUbgve2scKizYBjMUE59/s
JM2gPINZhQt15FqNeA4uccYqS/ot8m6ky6lRALOweqZGpf1Q2mXrS9F5phR7pGr8kh0ovYIn0giN
QPrnAl6NxrRUmB32KcjzLfkxx9mHh6oNhEWQ3t8THRYU1pUyPsASkVFfnmOejS+pFtksyt4ISQI+
e9J0118yXyQ9bHUlaouNt3XeKwkAYbk+ZQC6TIpTkbBnSznLNayA6PmsFFuj/DKDnUK7aYYTox7y
6ZogR2kKCw2jPcv+Y7SJK7AQLC4vqmE8itXNEmvR9rZp6e69tNGvND55GoU8fiOfcKARcxc1otjB
g75kXnmK1AADnoeqdvXJzjjomXyIRxzzkfeWxnL8HxppO23fuCnmJG2/1IvklhMKOPGr+fTUXQ39
frUpHBb95zn7xKUuHigKU0gAJ1qFLmNT0lm+efD+ZrslPkhHrcnD4Rzom/6R6AOPF/jcR/LeDbFs
xbxdwwzWcHZ/iKGdM79Io9FAM3I+kmn0TJ/ITfLXh3rQXOrZt7fvtg4cwL344QO2L7Ab6DUGcK1N
Suby9F3gQxEueDZ0XNMJr/CbI4K5CzwvL82y10QxJzo1S6qnJQE1S9u4OcDU+G6SF8mKvXmQ65aQ
3St7YHO7vcm7FTR8zQnpfnwb1QI1h60inpSea1pI+NkDGCCZ+aL3tTMwtE0BGz6DYOyFIAOQI2Nr
eqhpQK5rvfm8ixK2NUt6DpCfzoK2k0S2w9GszwDhNuKG5tKggbEMWJhNgL15r+s7x6AP/KFa5HQe
580eF1dP7cMJn7epBkXBZ8rU5GVLuSIm7BCUY+VC3aYAmnhdBr1JCfBYZ82ed5zKaKkRvdcWWyT2
lKMLxCZpX4Pc1DTCYCtijx6sJMy10+R/IKLxOASik4/urtYDOmr+jgtT5XQHyrijoF6Se7c1QGeq
9Bkd8HArJCVCe73nJyC7xcedSTo0+1o0go1DIyqYWW28O0vf4iezEnQlEv7XvK85YfDHB+nUEh1S
uhhXuvq5cnZ/0+Pskt/MeQEtqN2IAwfgWnrO2911+/P0LzGHgHvz5BPLQqwtY4HwhwUmXxG0klg+
VcZ5gbNV+LzoxD3D0zS+UO2NCEs0gyyrywYd8Fcm4vZ94O88KBf7C7uSHzA1SeHmYhjGVidIfgLA
4XhJQD3nRDr711l1JqWhGGSYqD2YME2ZTmfkDnGfZMSrhBxEqAn1kWTyzMwJqfD5uQCGfoSTWFVB
JpFJ9MonwXwjAaYtcCco3RLC/odEu3TpUtxh1TD47MspFyjkpnGb/Dt5QHEtY60mgl2f6Q/cLNyu
EgnJcGqBJH2pVbfPB+fyl6wSvlsSNo0Bz4P4u5c/hEMsEbZWAmiRS3/v6IGXY+fE4MF06WDFATSb
NmgSR0PrQFZ4we+cSTTfeqahABRTkJ9rMQ2UZToLkYze7wrazcNecF9dTKlR0Kr9CzBRwbGBr3J6
EW2jspe9s4lNkWKAmPso55TX1arz23ZWYbiTbwFwgvgqQjDbKz8/nSL9GIR5WYO1qLVTqAXY9sCT
6PvCxeYa0QGekL8kZ/8Wwae7O7oZFgiAhCRgNfX2lazWkitbPKkQf2gBCQ5+qpuEtT7NLuQHzGy4
IyMYaz/YYq+vncBq24URhCYfEY87QdpQ75rafqZsTWJswuwKD6y5vFRkZ+rtPP0j/d/2C+z99cqz
K7B8micxsWBusqsWBJyhyn99HRktV8NyWzGgCP/IVb9IAqqMzTArcRucgqmKOU5Bj/Ft5AsiMhQx
xV4kmXIvUyWpaBq4h4qEwNmDWHyheXp8+Nb8DrPz4kd6orpz9I9LtHyUEizN7y9/rn2X2USq7UsC
vFYsmOERSW0vWMiWJ5yN/Y7y9rYUtsye+TQgzKTe6ElrOLfFALilLtVJ/SLoKcUzH1U32yz7IuzC
Ej1saTIqXpNEGPKuJwXnUIgoVyZDd/4zHU7xkz0XBBQRWbKjlOS3j7rQLEuK9wLMcc41yHIW3NPg
ue2h3MF+1oVgRKRGGxM41+G0/AHMuqzbadCtKd/xHJ4B7N3Sbm/XFWHBmsthSVBy3FiB9U0OxKMF
BGajLVoXNnt+Bxj/0bEzkTFoqnE03xR9O7VX3WtaVE4NWjpFOwJrXvqw3iqD9HaWOpS6oD5CGu0f
K/YYK3pLqKaN3H3lzxxkk8dMWL+WpP416Sb+zg+V2ABNLjnGx6DxmECsBYSXqE6MzRW3gkan1Cyb
grvcG9H4jaT7UH4BYzWrtv5ucMqg9h9x9QcNneSNiMC4ecCUtnCdN3/Kg995QpkpDAblBlNgga01
DxqqKsSsRlhZkv57yRaGJcbKcQUhBPEUSNN6TtpXss4r8/OuzqkivmXHUBB02CAHms2kfuX6p49m
CzM2w6E0AVWSIaV+x6o5m5Wt48t8T46I7s9koljZvUiBMKuZ1hCghsqdgZaNPaSGEPuKtP4MoBNN
MbBr2Sg8Y+IGBAyw+pkI+oaYJoNE3nD88yjetdzw1YoCN0xXLW/OBARMkEbRh8GWaFccUztWr5Sr
wLR/aEg+hpbuWVaifMz5jlQAkeIL3Jao+5gZHFfE+YAL0HLno33wTbdOSx+Es6l7bCapZHksaaoJ
iwHXpxXIiZ6S7gRyBo0+skvWpTGSkiIG9zJgd1PvSrnaB6OujucNkosMvh/wA9vgPEbnpXKhR/r5
vcxQN+15cYB45YttsI7uEvXt9Xdsudm4HCaoecjxdxp94rfby/MnTuNJwgYTEg8QMho/GNIGDoah
DwQylKRlvB9Uab37gOyrpl4/ABgOhe8eZCwA0R+HWNLa3KqTr7endyKVd+sr8DYrmgr6/LFbrCG/
ZJvZQlmWAKk0UDGxg8oldEjy0txUyoeuXF2NG7WypTVlf+cV0hyOEiCUZ0vlDpaWRtAYLqCAtmtz
aoYd5FE8DjOuGHH+QMysANbv9HphLBe8a/9c91jW05jtK17eoGdJiTYSruFsks4BWorcgpXiu15p
lC8ZAr5Otm5A5gJU498yMU/ciJwcm/27YgORTzWeXj28obtSk8MidLggQBTJxm5vwe8dCeeNMmte
9DJgXr6GeQ2McRdIXrI+QrpO3dlB/POHrOTuhQOtgDuLqpDrjdpJabBjq8rSuKNxA/Nk9zL5ya21
L+8Dcd0vJdUwqvznTsFfK3Djs8yG5HnF8RmdOaGF1Q0iXdb6ul9Iyi9pR3DQqwemIihRGmjkt4lQ
mNST6hIVzM9V5OSpGhYwssiZWXgtRWZCp7vOjIyXVRfWpmqGzT+39hyeXBbXrXHb6ACHt5qqkTVR
gzlQ4ZSt5Lh+UN3q+WxVjXiS/IbEok4GchMO3MYqFi2eUHgfgOV/IyqQMehn4DTWDazpzCp2GCJP
bPelKfCBj710JVVSGz+FiPbtEAVAfz2DaQxUiCVeiXKpYcGqUXvR+YEt1fo66AsGdmg/dh6Qxpvz
mgLyZBBIGr39xZPCE1KFbXQB+B5SBquElOLkWcMcK/l6CSbhvhuIBQMR3xRRy9kuqne7IzFSOa2/
XnSrD028b5TC8kmEOlfAZhUFeurCi0m2Ip5BkiVqdKXOP6EFwgPlt4GtZGJvluhBzqVD34K2nLkB
BZUk6uFL/8+vbFY0LV45M1bW3LxCEvaOzJE6gbpXHyxSrK2eavwMc4ZmTzUbdEjZKcrJsQr1cEV1
Sx45Tbx7nXpG3KYGDr7jY39qDHYjmWSwpYVx74xVIYG7po1UF5UAbOLfK0l2zyd4CbMkH2+5LIwv
Na9xYlNIvQnWvN5Hi/aKdekfsaOuZYhYvqrGTUqqE1msqbE9LlDTnuF2K8HZMQRlUWUwsSCd9F6j
GHONiiDkGPC65n/mT0wqKI40mxHJcJ7crNcD2M8RC/4DUJOgLxt5mnBjwBk5q6T18e1SQHnXTuqM
u5ozW5SQHUkZE4O0G0d+36RA7h2uMJDOk+gEzc8KiKZzqLMIb+3hgb7j8Sf0Iyrby6NqzWAwWNca
mJjkTlvxgfCqBpJyPREeHg+WeJPwozoAIAyhorZY953nSS4j5O1NybcRCVRe9uD/GKl7QaDBpVv0
nKhdw+NMSfOKa9xmh5NNTXgpxQQ4NgxOEcMRErA6I1VqSOZdCZKgw97HAwvtFHAEmYkUAX+sY8uC
sslPciBC8rqGTPWr3XwUU5z57pUoUfUxaY3oQLKvTnAafNEtj6yFqbMK95o79395Rp7ySj+H5mLL
fjoBN/gXvZnYrrzOkDDRfwzEz4sK5PPylQ0a/0NQrslXz0Nokiewzwf1FcsppCJG9LbQvC0gf1PD
V+OrepZo49dN6PLZ22+W6UXBTnIrV2P5GlMSdzwMTa2JX3vouvjeiRwQS69XktFCPp4KZvVDy+L4
9xpD7XsSY8AQkiV++O83g6FScgeqHJqbS5pZIDi/w12xU++U+ryu2q1kObJPmRcaDG/u7q+QjXM5
lpmgdZzJ8VelHJgDcnm/uHMIQNHFHEsHgv1Q6aG2LI4YUxmTJmvjdvv9u/a0wDHvspyCig+Wbu8a
xZO6Y3l4ra6zQ9/5Q74jCn7w0+0M3S4zJ/yJwmX8yLNWl35OwPFP75CqMD4unOhlqADLM1yvUWL6
dg2TqutCY9rLkxLKqGTZhKuNRmIj+LBvfqAqaqUPzGABcEOFVY1J/c30287XptNfI79kPajBnxKS
l5u6fNlO9uPxejqy4lIFKEt/6/ne8+LQup0T3uFcNxbi83VCjzQXSRbFallryDOo6LX4yVNt4t+e
u72GGZadgnGelMtct2FUux/m0ZcDHQ7obNhNCSuNMpyqNTMTZKDKKOhr0eFL6c3SVf5RAS/1rVho
PUVTwG4NXebmlmde+QUliszUToX33WIYbZTd5HI2BVRXjkJFORjehfRLk85cueOmP1WpF7iXpnGg
5RF0zZi49dpUJYHFbIt5jUnb7b6LKBKj3ScckFkUWIFB6N68Lu3TKEikiWzThPPffUc1oIAr9m9M
sQ+kzZODdYJX7Xdzsx8ydayp/4zLdshvPsN95W7akZFHUabpJR8yfRMmjVqlZ9qSm9lEH/enOZ/k
hBPqhuZlw26gNeWyIxOyqTzOPt3U/zZfpW1Osne9DiFAua4tFcdJQa5eQeqeRZKzK16r2F+umd64
Xvca/crhjiBXuFRXmI91koWnqS4Co1xVMXrF9DFf88HvgrJZwpZkz8GZwBJLJgtPQky7zSSrQAEV
Sf7jQcYpm/+yJCxt8LMvUr7TAkUsVSlB1UN+PWGiCMPuw+MKNEEg8uZwFLzS67SQAOZU/QRSAyrd
0jIOQ97k503IHf8henvLLMTZWYYPywNFf8pqt6MS4ddhlwkn3qdDwmZjRhv4tezfa6Spa49EaZ4a
A9sZI7H/xD7QIAjbemS42s86m05sVv7WPmCf97+iWgwBEnLJU0Y71YtXSvcVLWEbardXvXStmNp7
axWFJSljoanS5K5I+cmO2Ewx11+niETKZ2RSfKHE84KzjJGm0CKuseF1ZUo2mf6cCbhdhNV/wZ3V
HG9c5LGgJ3/ZgpohRIclK+V5d5xFQjsl9d7YEE5hr7g16pmi8DZ3YO8Dcn00QNvWKULQhg1aKWQR
rTmSZdL6fbRBsQhpsKj0CAcUCxTBiRHyafH6YH213crp6ojg2CKtgTPwk83t5LG66O2U0EyoyPtY
IymaUwO4qhi3zQHRd87OUa3svtQLiNBz3UuTYM6SZ4h7Ts5SncaawpT8HyU/O/nsOa++C3s6d5GY
KDqzcTjPDTphZJybeceP67s2cOe1UQloxJiU2VgSDgafj7cpQnpxsDiVU8OObutpHaz8EKiwn78z
T3XX3UvLtK3zOyHJcQ4cIquFz1EnBfRd3U+9SGDWKxRCu4cZgW+WR2xId9EOA80OljL0CQy6atVV
QcaaCewQuO/b9uR6+5Rj0WdSIAH///YndtKeuQaM1DAakH7B8gi/PXzGIrZnV62uqwCNKXl7RHvV
RK6cNPBa4ccgikFGzbbJot72LOVton7yd4JT2DSAcDJWXMJ6aKu73QLN4PoIB6K7gHDCnEirKUAe
K8RAFYYq4V1C8v3hwsZFG5iTmIwUm0ITbq2yY6/Zre10zOujeJ3cqJg9Ha1/7zXl69ufVL1pfxZB
YYz/X+Zll9ClzpN34dZBEyNa/xfGrs5G/cGVZDIGRrjGaYyVI4OopBBG8l39QQ+vXfwx7J1x28Sa
O+16EAMZ/6ElLFXL3qnyvDYPkjcbMgOX65Nlk6HsAixvR5BfVJxFwR+0GAi5hax1+KApFuxatgSF
+guL8QgNpeKorR4OkZcRDH9ucR/6lusNjkeywKXp55Jv+DCs49k3duNEb+4Ahap4/28k8l7g5dEo
mXxYBpZ/dBQ0pE4czVJbGtf9LzU6pXzDWcQzAQVYLW1g0qGHIR3uqFuctf41xlQ7cjOJY8PvjTiR
PWhukm806apsdWzUFYmcWgkvl8Ub6FUP8j5sRPdhj88OB3YYDc3C7SeVYRK8uhQWTVMeyjCCFwcf
rY5OT2n6k2FwLvYk65+Py/Zzbo9S7xQRV3Xgvdlf7OOn/IzOXSDfE+wa/dD+KpGYRmC1CbjVMO9y
uyXIrZIJvLy4+xBlOdPInfCQYQmWuWWieZ4+g9FLigoxwNDplCeMOlreYrj0V1dIaM9z42k8XQy0
wAn59fG7zWKXAaF4o9wVCKaFGCQDYK/qCxXawBhGTeXFYo9+wXucTZjaKfwnX8F2uQY1ilQZwQA0
trV5kGQse7JUN0Hc0qYftqzi3TNkiO3BtLDhUMBhArnFJHblDqEY9Gi77Hzh6ORSKglBSwRZ8mN/
htJe442h9oSEmDjfcosa3SRLtDv9C2Az7lLSA8+45NjJgWvbHB/H5dAxLg9A36Qng3Zwn0Y9IDRx
V0bh0K87c/ocNb7QJEYInBVtb8CNX+J/KNGTLQWeaZuFAOQ9stQYkVUk1xdIuYAKxSAB0cAZhOQv
7v6aXf/KMU4NUc7vp9c0Db5AayBq6AqhpnwVk4PX8UKy7xa5GGh9qdPAcluqeimNj0st+7/VmmT3
QMfW7hI2/OnpgcjrGL5TYnI/7cwmmZ8wDj/22Zj3rULrdHP/xCN3dlwNf5Nno/DFRt1rEG4+Nb8l
yq1wGPq36FiZE2gGUZuFrOtdF4Ke2xxyQbBI8EPraWjo+HLVGGtMAPEAIdm+P598/fRiAoam7Xw7
udHvClvQHVM+qaKCy6K/o1qjpEy5XTJKydeZU0rHCwt9TZ8HxKvykx8A2uMRuHF7Ii6DjFmiskpo
ecSpWMMJcKjiPFVOv//99PK1yaH9nDOcUyYjVUAGq5oECDdZwz2IjUeJsir/WY4QpCw5f+rCmV83
Fu9V4+BE5en9OrbbEvcVlabEgEtuv4Cir3jpSfx/c5SBm+DtdKJICrwisN952zvhKC+heJmx4CE0
ovGjBZoCAsx8G1YSHwjCN08G+Nkc4dKnrVM5Ng7qyq0nMxqFXipAdilKK9HD4LEEM+x0H8FGrMrL
bZ5s9Y2B/FGoYMJyeEh2mdJfU3j3tsaHVycQTFi32ukUqKINnKz2I6FPbK5KUiomdlrvoWTNEZP/
tal/yMnCknxLkcwg+HQyLFkSNmIuXoxhWKEKRbk/mNZxLOBH84QvnD6JAhibKkayAjb9D2wVgC40
yOVYM7oQ00oNGJszrOaKFXZvaTiXVsayByXk6Vo8a1cZn/1VyW71+g1GeityNrsSMCpfA9qpCjMp
oCF/pfJHk/C8vSOzFIGuSywa34dtcLprxeOYNg+YW/SId4lyWnRn5R0sRP6bv8rJygm+vKHoq7sm
mA0eBgdlru4GiKRNJW+qDJjW/uOCAQA/6166xkq252jzJY6th7E9e5S/wc+wMvzXya2v/uGty1Oc
W2ALzk2yCvigyrg0CNzng+tns9gQ5POLywZSkV054c1pJHGyih/M6gm2uOiMO9uCaR5uG5/O7qTZ
MRPE73wVgdoNz7Hyqp4RfDA4ydMKbSQXHHMCQttprAUPeTxIIXEdFYBiv34ZDLZK2WZZRmes0ATi
5Y+zS3yxMiwqSrf9onSnBqc8k3DKisXP5QXBiQinWKa+uqMTKFlpxKCSLu8Khfhi2ssj7L+tr2HV
TM/yb1fKlxemd0BTUKGRQiWj298ml+AR3hOYQMH/uH6wMew0ZZmQfGGJ/ZvxAdGqWmYYxH1JLXMW
/Fq6ba7mtztKEYKVNRWOgw9QKJXDFhCl3W1PNqAGQ9JxCWhtZU0IBu7zD6ijuYn90SeRSn8Mghv6
T/F6i0sHi7WS4w1pNIKcxHwZ7Gq6lsH1aLaTs/votLEKbUPHA0o+iqk3QSNdaQOOwoLqcjkqV7+O
MuYlo8oCqku8Ak4i9udV9imT+o6BpDBGYWduHCSRvfJFM9Gj/RynCREl0RyEWKtt0Ov7Kea9PNJl
ewLpDmqI5LZI9Z5wuYgz8h4/UR8SJpaMNWAywjGuXAfKGfEr/m2lrqDpDKvpx/D/whm+5Yyeh7J4
M3Up2627ZixpjeUTd+1h2HpS341LjWklgCYV8mmbbfMkjq2Dlq3H0GL8BQBMvEtBEQlzhSlE+Yv5
3Aywqdm868fA9Rt7E2YTKxJ6SDNOChPlE9q2znJnTSN+xsWvP5i2bXXh3qCAYAx9+riq1liB9iIT
0hIaqOXioUdEzWZsCtxRspSd2k6XiKhn49nzjdkAQ+3f2mFG0XcnD+4356qgOXBDm2u4h0AQxbbJ
HpAl/c07pcMD6Td5UrI9oXiBJJ8k3BTiBiw9GIGcPEwCFlBAuF9d/Z9aQohUTptYDNOSvnuZWFYo
YYQTcZzc2VKytvQZxplex3h9Dhf8D5ewxn7dkr6K56882jczSXq4rFTRsBO2M9phMdS2GDc8174H
jWU9HbbMDbEbPpxZUJiJOIrhXUDBDfycMxv1t6bHivKi4/2xWSaHs9osZ9Ts3aS+8kqZRsI5JR4G
/eHAD5eJcBc3f2yHSAt3CV6UlL9MkYa3Q+gcZd78NxMF5qiqaOHgIjcvI2/zvGgQwmBfbFCq+mpx
oWG3tW9eydcZ35yhgn+s+iejLXgcalAYMTvt4DTaLJ7V4Vke25VnF0kp1km4ACvP/MA2M+AbrbQt
kMJwdP1E4tOQSFwbD8bgA7Mj0LEgvyX3wSC+RT3rcB18cdZH6BWcf5I55xyqNw2Y6Hy4C8DmIGhm
2P+rGiK5+MhCgDQYeJiCIFWAJhlYHYyrfAodcUzfW0wr1ym1jIb+OXOoyRO3RWR/EHnhu6VE1qHr
J82z6T0NdORC6IIabylfLgKM5M78NHCEye0UKwJbS9hGxrCDY5zYLV57GtTZ0twrRIqtLp//ZKt+
+NwVbg805jXW/NzJ34oOLALafqv9Lq0xNU3uC8MdiRhOz/lgnADRQIzTloyduNq0P3F5g4mUOQhr
xDFmeIGZTOILndCWNWICDwZ2KTKMe59i7mfSVnrXbc8avowYpoipAhpR7dP74jU1Zc+9kYecsThT
/MxhTmsawbzqrayssEEMWf1PEfhI6BlT+hcTof0ucXkTYjy72iYRlzFcvk41XNpUUY8HGWUCRZ+C
el7GJ2S7paLY+GY+WSbDCBFz1/GSSEBmlgk4EW6DDhX6ewBPQIjt2sUz1aMCW88O2v9vy2moyLZq
xjcfmO1TLNtg19ZDMpMca3hhISKXZzJg3/cBbQotqHYmIgKACf5XTJooKbDTo46fija7n0OgHrCe
jFWoUs5cygPnyAKTRjpRl3P/zWFY5g4dYIGfuo5A4sPbG9TtYfPLmwcxC/IjV7APsnilF1zWkb49
lUcbQUcmFrcP5/vBYZgO9G1NLOvTX28zdiWtt8En4uUw5RlvR0Pjd6QIGT2F+lX6LA2PrOdxNkIw
GRIe9BgSl5iRgot17mLTh1xVi+EHy6TbfAzYCVWv5eZdSXeDKvu5kmgZcDniYvtPelVi3rSz2UcZ
kYtsIOl0WSf8IKcz0+ze6IYSqqCdDgVqao3A4xEG8UQE8VsBFgaHVr2mY/3iHeZjE2sfiYLUyWFU
mVojOK0CS47H7wqgztxImMsTtG0xbfKkXn/IRrWtnjccTQ0gLs+jsX3Cf+N3mcebS8vnXk7cPML8
vfu+NyocGZ/9ud17KwDyvi2VxWa3WD0PNjRkA6+S5hUJn/YH8OlpJq4LEEsHhrgFoEsiS2Wk05IQ
Tlu/OnSPerX+8RttKuH9tSs2kUchBUZkRFoMY3Mby12G+zYULLvrQxRp5Kl1aDxwXvu2GCTW3qBv
JBHpcrgB1jy32AVJEOJzGWgh92s8IX43/wMOZIIWtLjfcTCG7DItIQJxUf33mBUXHcLS/fygMeAZ
scDiF83d5kMJXWNHAKisLUPOjeIXAZdKHDfq0XGtfFmThmkI+4eHPu3yipW7kv6vqg3LHTr/WQLX
rrXuC3I2V5Vx6gMgOFQfR+d1KmID3p6EsUHoRZory6hac/aSPiBLkLSt8VNRGO2lHPL9LcDvPtmL
kXcNAToCGbsB2pPZB0beJU8KLzhNclPB8utTus/VfYiW7FTaEwEiGAar7kWIQNyjJdd/oNLHfelV
ZU4I3jJxpKDsfOLC2WGJMoYpL+bQdmsQ+Mlh2m6/hwOqTpqH6rsN/T71GaS3zWDKW6ih9M775ef0
fc7Fnwu2SWkEYU7bzB9x5c19nLDPenvyjbdK+U+1+Se0rPEzkWMtl/N8FVGHf6x9xsZyn0TOdqX3
Hbzupr3KEjqqQCIr4vvQabCT0htTNdrHeRnwNpz7eUTBoxaiqirK/fHgUi7q5Low0aWO6+KgF2+8
Prve3vFzl9vM4eTHjTEL4RrWE0/DH0FR/ctbrFdgSr3lavHWVh6NJ7CVNNvKNvIsw7ic5gRYEy/i
lqHYmbRBLPbjABZnxAJD1JEswsjmZkUOIAcwOiLKMxfFEQgpp6HO1Nb/YyI7Bb/rINIXpN4AtVVj
8GIn2vC0QgQNAq65+ksIhdf5vP2Nl+opaAzIFSCJlwYlPHS7vQ1OT8VARtmTtnXBZplA/76FjvR3
E6rd18ETlvCIunrFRsPwkxT8BUzoHcfu3emvOUJ3zrHPCw/EkaKqPXe2ZaWPGvKIkqXFMwmnUS4R
S5n02Ptndt66/sAa5c7EiiNyAwI+pl/jqCfWQPkJhef+JMAsqREXzbzb1SzCZGbD819UtYLmGAFE
FxydoxZXtMGPCUmt8pr23LvJB2BEv663oFwhu2Kr8Rf2MnT+HaFQ036wF7khHLEzxS/PD1fQshiM
5a9VvYSn52xx+IUD5NZAjaSdu2+k4EtkDu9LTpBU4++hf7l9alPAj7npTjnKgSZR+nQZazfVVIZ9
3/LX0a8PtskctJuhEfS7Dp5p6wpa7YGmpF/HxyA+xQEZWeXSn8/MzOGUpzfTW1Z2hAZKBtKZU7D0
c2hwdlSsDg2n1L9qrZiqBXBw+SicdHA3OO0T8nLJibUHuwMSeiK0nIJPB1kSHFr9ZGRztrV5HHFT
oG+AUCSrWwuVvC0WSowicZgcxUPJC1x/qxiqNmR2kQ6xlMoTW8+Jo1FLmVZagPrRtdPmIBLRlZJS
xz5U8DrB1KWuhBR3eOWF9ylZQWOP5BDAoua7eGyjRZ+fzZMJmewq4zL4ngFW+DOvOzs2tKy8FC11
d3xvXTsZ+UJ5Tb8G+wosrHjk9/S4s0NUDufNJzU0a3hd/YpCCHjMfUq3v5B2xL4iLJbmm+4MRm9j
JA5o8lwVBXagjCpFbWjoE6bYSsw09pd4f2C7IKgGvbmHytVSuCxOBs+gD3vqZi+IwELPh/cSQiXi
qsHUcznFXrnCEFxu1iivv1mAQqTbSHTEMAmlg1McrqQj+aaF5Wpz9JSu4KG3aEWSBdcuB5z5yyvO
Do/R1zgy6J1RH0Q1uY+1mEnJGw9wsG3AtPRGKPr6/yn/Xzhvsy+3ntTbRTWD3pQ9r13zn9hZz+ih
RfQzR8zvtDyZ4m+TXM77aTRmZtkSMWnPvV0RQyz8UiQJYJBLCgslfQO02VcFUj+b1OxsjgkFiZ26
lJyFIR3e+EAd1+wQ4sdozKaZdqT6mZKPPVVeXpWcRHg22vmUWrCaSRgUQ4QuPV430X+9pjA0wDa0
AnC/Wm/rnG2nItJ8JRTtSMhqUOZ8EB9hMwR03p5H7ieXlD+Nv9JNvVHUk+aC6DeeqTQIl+g81FcD
blMh5/ztxmCxcxa/7nHj0a8opFt70g7IcEY396H06gvG7PvYK0L1CVtFHAXKtpOG+QgoW75yrBHI
VIWH7PQQ8Ng16ACT1qfM8zvmoFfU35qGbAfSiKJfGB/ksaq8JKxsA8yj93/yfRpiSyLFAS5+5SVp
nO3hfstYUbHyIYSvzWhVDxQa5yZOiqEBRnX99nO/9EmxeUSGxDlUiW1RmPqPQpqejxldkjAUuW9A
s5sBKB8QxlbVydEVimYIcj1h2BwMR3RlY5/l099QQG6HK40ysxwwL2CHfo7y+NPkKnfzRFOU18ds
BPbez/asUwt22N9YnxYZhruZZzSKzc7PbSB4i2zn6XHEir50w896ID3DgCyUTjucrJxvKyeHb5fx
uG35hVFUOwDzl3Olj7TL9pbx7J+q3Rtj07a06zFhWcAKPIQoNtU6Oy1Oaxuko/KFxhJ59ZbfN7r9
QzuzQ1M+erEP/gI8Z9AVTI/BpMvrOiZKFn6Jp9JtYXPJNCx0oPuyN5fET0NCFd4x9go5XGAy+eAr
9dPsXpLRGYQP4A1bsC3/oRgq1iKeUsiN9OotGGshbQOOxgdHy8r4zkkVtma5iHDEJSGEkWPHBbK+
3V4woI9NehRZ37H9+KIop2pHpzpAfP7yOlAl42BCeQtYHwtfxWBTSPwZQXDPj/14Y5jepxA4jOE8
RahlU4G6rWH02GwhVs1uDGHMHzzjAwk9G06sKSmW6DAIGgo36+4UL3tL84Ong6eWlEQbX+HLJeNm
7X1rQ3SL97n4oQNfqcnBCWbKrSmhroVsISkN13WEnaYtz6IpstU1sokuU6Sjy7ZAqwnFp67cAA3Q
0H6DORPyMwQs/DArfvI2faSkVwWQ/u28RkzKgMoclwWFopN0uhBK8fofb+0XnX7a+pk2MQmn3MKw
rTviDLcVLQLOOs1jLoZDJSCAw13ij2Tv0Mila8Gq+KiN6gUyoq/a/yFvF6uKoz2/G8mQxa7Jf8xV
r9Zkbv3y0D6M5jvoYx4fDW7Xj19c9rpPDimB7ugVAH1MZu94s9rFLZJ6Aazkdwk8BlkdWZ11Idha
J9DKi+yOsL26FYqWRxGq+lDzt6Kdcb4IccTWdWeWokP0+bINiPjHvDR0eVPZVK/3wOjB/PpMFU0G
XrNObRc2Ix741WIOKTpU1wyZeKAsktk6YcUHYu1v5yj6rm4bJJV9npSdO6tjbv1UHSR8u8or8Hem
492ASUSxyUDfKHsGsayG1FSiJu7wsA70KP5Rivp7WapgkHrFabWO3VyCNkjNZDZKcMOfRbgN575N
Q/Y3RctQb/nH2ZD31KWTlJ4OMrYGqPwK+4nRgH0tKv2xmU6ZN0VEKw0Pu6WMOTTTqbfiF58c7cM8
A50+VJodSCV6zr4BB4nlYSw68ZCCUqmHvzX6XvV8fheLX8Lkw0Zu19u6OefYPcPPDn79jSXDwfUn
/d6X8u0fqZbsdeDh/eqHJUeglA3bxzuqW5imxGfmm9/b+IJ+0nVfTzc6uGuEhGwaQ8vo+fodiStF
rjvuysg+HgspK4EpzkcH08rxL+R+1zVGGiMgQhTh8PvHKUCJ0jBPIjERto47P/IYMVnyDqUlLrS/
47XmIGM/xbPCXFKlSa4hF3HxvuKAK0D2bUniaAFgEoCgdQlJAudCss8/y4rxwPaOvOV8cSoX4eHl
rIQ5CjS/z2pJB45npeny5ID2Kr6unoR+wZ3HZk2uKV1tyoa8lWzL91Lxah2PxA+BpazLHGU0hydA
R/2E86XM4bN2ilNGvKSCtqQImlGBXpdZQbgTwk/u9vNqZVhsbKolFixKjW0roy0kOMiQA7g4KCEO
F+DKC15HOq/N5ZOydmzz/Xo2NjNOj7Em19VsC6RxBi6mjRTtu12A/3dYbxwBltTyd4cIO3IC4RwZ
ZUBjh4k+6zDlZ51XmhEBHqq0j76vSpLXb++Txs/+dyKm9w/Obx7U2Z9nxdM668laGB4WN459KUk+
TP1bBRFTJ3rSX3WHAnrSuWhFRWqiOvzvXL0S4vr/jGZTZurfV6Q7cvAuzkelqZhMTqipdk8NDRjB
uffkcV+Yii1uc8ke8w43KtowQojyJB88im9ZN/TKreUM3T+CvyNuhZn94or2MLCe0UFtGoevhDHc
WLNZmUIi0lRrgG46xWKPRZgp4V5mB1eEWY6NUj5oR37aK1i+hjB4rgml58ZNHQnp0f25DjOdEyDB
mPtcyQdL7g7arOLozvTULSXhckOidp4aWGnmAK3e0enyIpjCEUUlrG0itZpkQoc4S8AjjQTfy/bH
V+5AFirnnANE9t0/Mm32nDXctDKJIo+vMuf4H0HHcfFFQdU5hjU4TI+sUOUCg1fHrEmuDVpAGdBI
QqyHPpRS++mrs6P9c361jG79k7hWiKfEE29VEnExCCQd/rVtRcyQHPetLP8O/hh7qRTK5DiswBT7
UpXiIrYhfFjr06hPVJ1XXn9f4kWaLmMXDIx315wMYrgajtfsBVaH7x+z4TwLrwxeuDA1vvbVW9yY
bITKwOJHqKJJcS+fe/lkDy07cb/92/ajyRdeVLrlGMA7NF6xw38+6GyjVNdfNrgksXUFhDHKM6En
GX69FTvVc6zU0bMmkLVcDRXVMNUTWUROvaQ6T5AoW3t1AhCiVVNepBD7D8mai7RnkKiP2H0qx67m
wCDcWmysve1cOlOrvYwBNatDWbWQ9vR4Yw1KAL4M9ws4YGSCCZhpo3j+M7M9ITfnNBOPuZsOPZ7m
8pW6007ZMjCBLlgmx/7fbBirkEb3Mbnbw4dToszbyCcjFW3fK3z3UhOwMPxd3abq05z8aViZhJ12
mkuo3gDGPfsBXKW5iDlePKMXxPRgvsX2QMpx4sz9+0ayH+Mp0Ogz24Yk1/fR14CcmCT8GCHCtDWJ
2s8mO26QXzIoB5rEwAFCwFeD3gCMq55e+rjROviEdvBDsTyTijo++hWSAbm+zo0f2RNra/CmSnA5
snCT/GqN/RxCkZ9o2ZZgH//tEpZbsjswlk2v0sgE2G2W66H/UDyjsu9wMlzkZVnC4EmufEEy5ra7
CSTCJ5nFzJ+KEnBwVWnOU2ZwXX7a4vXSaqpFHAfZ4kWYlEElp8Gs6khXpn4urNNEk/b6+suPmE3f
j8n6+Pwr08sX20ko//Z5wCPi5R5WW/TwOPiSEyiX90R7lFWBx/N0nhM48uGmT319NQqVYOAv4XHZ
n4OY+gEfk8YK4HDOslEQUqH6CVdfozV7jcVBM3Vhq2E9stPkVWgcssQV28steIOVIoh3sCOSLMj7
Taj8HBZOphKB4Z5p7UlIzmmDRJm4DfhEy1HEN1nWVlXwTJRJsZDs1VFoGpIzMSWXafc86zovxCfc
y8uw1YnwJs5hY8slUhHK4I7KhM0j4+5RVIFFV9s8RGkHg0rwQJRdg/pH7sujdTMxz3QUEelHh3km
Bisf6sSxkcTH5d6CwslSHX+aibQMhk+KWF87v+572Zlq0og6WKXgRM5GfVLv+EJWsQ82HO0Knn8Y
VqGnITVFGbFo0Sj6r87lQauwwZwWGlPqLVMLajuKW6JT6vrsDSFMgueeVMkbEi067ThP2X8uBHKf
cF3lr4Xsmi4ZrM/Wr30iHrjfXPsJQ18xgN2+LkziUFO9VItDsikrhYKuEfumlcH+EZ1i9YNNoe39
RxNBdukuubzq+yRbskZvNm8ECFAAWKlCsGEK22e4ZBAs66BfcYAleNauEUCFK92R8dWtG7iFLiAp
0J+iyDq3SB3Lid7njy7t52AvfOWdFNqmXXc01yzQUaQIoC5X/jKP8m9g/xm3K+zIUS7HLl8yvdlf
NgNzA8t9bAFnAcnc1VjlrPUrJRId25QiMqHtMF0QKzcNXr4kcaZs7KcpZjg30088LpSb3v4A4Klu
9J6+g4s9peMyxMpWri+PMjF4xpFlw5xFwgOnJQiMOGY/o4CM1NVH/xnxjay5tp5ZqrzBYm84CL1C
F9JRP7/Qd/oyObeIhmrsUdMpgheBVpDHzuVdzHK2fUS/eV8eSzPfB+NBg7OdVb2DzXVcRSfrPrny
7Z5RLesb8QEIk4pNNFdCvzkDn2xdvWZC7Z45et0Me630zV90JeI4k1Ssb5qifRdTuwrVQo7tggiZ
kYYlrTPLAaeJ/if2lvqSMehPPG4x4flDQmG3VwxhGkZw5v5IImJq6i8cho3sZJAnu1QifZMmGHBq
HLbmQpGz4T3KyccEnLAbqkAA2HHeRayHLgDKLy09jI5SzqyMPcmyA8qfVwgk3dtE/CszH57pACJp
H3vXpYiakTAY0H+YTqas8BsSdFd+mTyRAPbanvPbI0evsRFE/f2My5kgrug6Mtgj60yuj0ClnyzO
ca7E9vf93z6UhcZRVqxpfzimrT9DAHO87e9hZ28TRDay3kREGW4lD16SnwfBHkdkpbOsTtouDDbZ
b3jYvjDx6HnjrLJ2vAoFIGzqDYS1ccr+RMVvwSb2Qa4xaR7QX33Z5+ebHw1zpjwWpDx3UyA0rxso
F9YCsQj1Y11tCBObEUTLkf/YKWLLqktVco/0S4B6T3W80LpHkMIFsjJ3T8RaXRe8qavOui6imSuD
FZlfhze2K8S741Tl/Sk6LyYxcxjq3h7HlxR++ZtEbRAvY+a7RDNVXkM/5DF4lDB8rkPNWtFpWkWM
ZuLiXax/qqsCfruWD9udZ1JSL9uRfXHEjx0RZVVpU5DNjLxWuqhTzCm7KbZba7w2Ff3MADnDIIeA
cSW29yBRWS8TUS9vv0MtIrOi4dh/lQkNTCz9JGS8/obGvZ1FxydoBjQQlaKsWY+UKBeG3DfF/9f+
R61OY5HsX1LtySn4bkzNeXm+kjNNUTyFvPHb7Q+W57lIhE/AfmjQHbxa/r/MwQL6Uxsf5eK+5r+6
HX4kykayT+COUnRWCH2qAMS9ZAX2Wjmh8Yg9hIuatAdk/WoBv2jOL68kKSvK6dkGNHG60NmNPASa
GCBkY72Bn9OUEZauWW8m0Je01BvPS0DHwd3tLwtO2GFTmgzqukyoqA7uTTa2qOLBj+pLm6o8lZXX
HWlO131ys/xmzatqUZbtQsYNyNu8Mr/75XrMKz2ALMxrIUvOrLjUimUyihrCayoJI5Rmt1sxwLYR
yMLVVBh1F5XNq692Equ725sVi4V5/smZr+hP+AbpvFO9UpyLGPtqo6O95zZSODuq0r1UIflfER/j
0g218GcL5NFlpvwplb6ELOBCghKsYRMRew19i4qAmSgsErX7D3PElP4XkHHdasBSAe4FSyA8yfDi
eRqM6bMzkoKWLpfiZ3NVdH5qSdL3oEYJRuTavHgBktwOzrPe55lQ6Sz31yStvClAcKZzAlBvhfsP
us6ssqx1oIOLybYi5W7MIAlpNRTRdemBjTEVhV3I1VuWlsW7nQav8bCnDRl5m9Cc2Xh+fsruSIVa
cvWoE+/SvGzSbD/ApqbcM5qPSNOMA7Pf9c8Hmc1C6ZWWGg+b0pSZJr0cnonm65aYFeIT5KLMI+u7
gmCFkVCHlmCebDwXWBgeAQdctHHoke9VlalIBAL5jqi4dYC07+CTE/235H3SofOwtd9wXsmADjO3
jVRRCXQhNvJiGjLurOzQ1btRLYVRqwqGwVBLzUFJeDJ/c/F4fkXxxIJKIywuaob0MmLerwwfZXk9
BszZLU7mqkV6oupJBMriOYSv7FmmEyqDMh/CHOfCD0p/EGtj1Dv9xrjR4MvqZsYCa1n6tvcK++B3
+I/B1PB187tzLUr1pp8pHuDdWcCUEK7fneh5SBKglgkUxj0UJ6n0vez4VH5FKF9NFgcf4fiDu3br
j/fsKG/Rz3gbKSvr5ukt/XvixH4LSgbfUVmiYaloM88gjCKr9FY6uDkZfDBsVebpxtT+Dk62vTvS
pQvt8SsYush+v0tp0Rav6TJrZSZ+GZG4tBzD+1q4FGQvODE+DzrQPxG/sWkNqoTucQA/N77kMm63
/Lk4dd0wa+696cJzxZCPkMtooJ4a8K4GRaWI6dCObrj42eZfZue4ylNtHpIY0PSGFL88oBPIlWvq
Z6515Vhc/Zf+w8yMS/+615RPNRBgFccJFu9GbraOyVP4XRIF69Zt192b1M8xFgOf0RK3Q+4XDWR/
GQ5qHrko7+8sqjCQ/kESIM+j+mcjHNifPCkqQusb2PXy0Hmje7MPcLsnxfsMLRELVhAaSxH1tNrn
1MaIRO70RPIC84CbEJDyk7kLoXlQVBMr2/kREguhUAdPzQj3XrBBiTYVdLHzYfjZkc2tzdr1EeX7
hD+D2PSdIZznL+KxZFAm/v33KQD88VwMY5TL28yjSWkuf8qRPpbmU+d2j9gjSergU8HoU6WY2SOz
vmy5Ja7nVb4wTff4zYxtyecEidB+BwQEjkSahFNhRffxhFXBQgOV2AZ1jgoK+9WfchenoDHHjS2l
mjm84Bp8lmpfHOrHtjS3xLkdCYVyffAjCE6FagGZkcBn+mSVq+h9vmCSgxkkTHXgc3b8WlY8/kEH
aoWnvPTMfou6oXMOuje0K8W6fwK08WFIi/TTo18HMyls2thbfucSHnD74lUlOPG1k/khqvamVwHk
UoVd7mqBRByR60AaanWGGsUJ3+CJDcfuu7Be5JTrqXwrg2+uMQ3lBnfVMV25+mIYtmEjn7fjR+Ee
UAHih3Sqo+u9qsrdM7dOkmuq+UkW7FW9yA/kEiNDGFfWHyEHQnnhnA2OBEEKcJJ7RWmGliiyOCxr
XI7G0fupzYkNkqVs9PHK6Eg0ZcXp7GiyxjcDcukKmSeDuEypOHjzM+txvTANnwtz6GkpZWYJlomM
DubBF6qhI9zAuWMURPLzl8jYifshMXITJ6ev68eQhIVxE5MpQVx2AXR+bbpOak7Et8kfVYqiAJdj
PzxhTA8XU+eBoS8hnd1CIhiLjwj8vvpRs6DsApQ0xnAB42BOIoqFCnPRDhZJx4b3kLK00rfjDZsv
1WehmEpaskMRlZjEaFi/4IlKHPjjU5yDnawSZ0WqWD6yvEBxnG+QlzZ+c/gL/9UvDa2zBgczrH3c
y8S+EDgJd2sYNsx4hOnI1Tm/BG9i04nS1Qv1z3uSolnodCe18D8lnkvrdrS73UF9OicNrB2e5Slp
hNsWRRRvtQbCoIO7fhQ+GvjPQggjE9ePog9YdsCWT+1R+ZMFbtfTk/sJBED+lQovg6WMHlUcro+q
+AP94ZwG7p5y+YhpbBo6yjCKU4MfFY50tDnGueV04Pf1bMu2g6uEpthayTbF2yEnNSt2m9xAFrdP
/CaFGH0CLUU+jGy8u7SRuVWXHOLj/fJOYj5kWQL4gBlT/8pTORF+ElnvTgX7FBcjvFw7JFZZ9z/5
ad+BEaky3x1B2Yps4k4vyeWY+eqEcoj/DLsA/9u9Pl0BK1PxdY4ssJHoSyyiMEdxg5DI+uVKETX6
qqGIInCJYNUV2UvZ1mnp9QI8wMlMhH1SyK8gAugIQ7mh2X1mDSmqZ18q9bp3krWp174DnyNO8OvV
MSdnmNcYk9vKjpG3Q3fPVgBvT6QESt6Pw/Y1gHoR4boMhrobfvXANjdeP3sDhgvGLnUxZnC7ztqX
vKkNfGoKVxdbe4Ivyxe25+hjb7elZ5UUwDVYu37eBhctdmcv1PI2Myfju6raqFZhPlRTsHEP7h4n
RCxawAckkae10p12YXROvzK9p9BTlBScsOMvt1bNOlhWsh8gV69FFgO1VFR8ZYbP/AOiOWBKTx3f
uGeKQ9gOsWE7FWoY8gK836T6ThSU7sQQXq3JkuIemeBv99AYy69YYGqVIT54ZtZ/LDxtxCvwzhvJ
TOAm3qVDfgt7UEeL0EP3E4vT3J6BYDsPu9pjecAts2g2Dxgo1alQkaC+dHCrC6RTzCSFTdF20Plg
H0qlHZIoNPM2ztKHB7iBcF+V+2pi9Da7qpcjH75kgGzAzWLEQ9iL6hfllT1uf2GXQtVlX7N4eLH9
gDBicIdqTkAZHad98PzU6UQabbxenPJm1GqsTyUyZDRVlDkhJaUEwHbyTYQLiJh8z64eRs8atQEb
iLDmpsCh/aWw6J9gRBk+3Sg+Cjf/2CtFAwZGP7j+Cw20kwPKFs7BcUtcp6/NyxG1zaDW219mUYya
hVnCqaVr05lnBvG4coceZIhFEJXVzro5v0gD+26/NpDJmBVTeTKW/aputiCDJRqVYTtI6VHxJZmM
iTm20QkJYZx4iNox7h1HR6knj/7tlaWOu23FPXt47IlzQ6rJeCuh0eGUowSwB966os1Fy2tPyYDB
lXXQ/l6BtvlXagzR3SNs0A81BqPYiLi6VpLRqxNuK2/dAMZbN3iL+RuJtyMI+HZWHUUBmgtYkTvo
EL5ZH5LrRqML2GKzPGAJNMNUk0hwQpC17eeH85WdkJZVxuN1Kenevy1g22gzXr9grEhTawNdywrT
biw7kH8IYxQq3CCiVb7Ig+q68O42w8M4KDUb3vK+96/t29a/k3+KEGjO6MI3G4MoiRqd81b369pV
tzWXGMz+vH9pZGAEul6YahZ6w5SEmkmX89ET908NOlZngZ6u9oHbzqUrdW09k2RoJcGohF0W2NeS
BBtAB5A39QzBU7IyyR8S6zB5T15Sz8p2L7/kjP6DWR9Y6AdBVn4xzaIZMzmsV2F8deY9Ut1WCqgt
VpA6pkmLw98asbYFv+0kdkuci9VDjvgAjjXQiInxyd4XAbwiOphPnpKnlQeozlv5GvYK1vsLseAt
7x3Ae8fSqKl+BEUsZYrsub0+DwEcdXiBpbo95rphAyHL3HwGP2Lh1iAOcx98zCd+d5FVHks+yFkQ
mTi6WnQQ3562iZuNYFoFWg/3NWwzxmIPgFlt7U0JNKjpx3Mu965dxcVHg1+P1O9LY/+kmjHIuBP3
b17fnRli3Ahrzt2E274feolsN+EY4a4bFG1MUxBUHjIYwHfbMFMqYc3zhJXEzvOr+gZjwWdjRyfL
S+uJTrnlfyaIYz+vKUw6WwkCmJUYl+cNF4ScUeKAJ6x2LPpupnkwbHTQp8FX9mTwDePGGAWtvJ/4
9uZfI3YT8s1LVrO8hgY9LuM5g/iiZTPrLZEGLtqZ37MBbIcTNmYFNZR5FOZmxE0j7yNh8dUz96Fa
XSCUQPx+Knv5kMmaRjLgG27OJcF78Idux1TUT8ez4FOOO8RMSz/CZk3SSd8hB7bWZIZGAli2ctz+
bz8MqCEdheu6uGiHMC7ZplncUS6lflBHqj6MmSNP8STtF/EYBVrM8x8/B9fCOAT4cMKKXmk5JdU1
NRKsAWFi9RCP612hrcf8QcPpaWpInTLP98H465D7PTdbylPF3vesHbV5ekxPd7kNVavcKLbnXuds
LVD9ULppILoBrgeGHdXDTFXF14f9XFP5W+IpO6S8U1Mx2Bk/1FYSZQXrdWH093c8m7Pfsi+1JIaC
OAfOG8c+iTL5dmTeTKARhCCz+mRWQzjjOA4ePU5Ckf4MGE1KUkYvR+JsQ3rNOk5z6HiyKZK+A8+J
6zngSHlyubpT2xIekBAKmCSw79HTbyfJyg7rYDpcavgRqwlpZH6glqTsWLKZsA5xN+JwmbMJ6o6P
g/WqoXogFRMCL3OwVVmXyOK5f5xnYncYXlZpy+8sDV2emW4rWDo8ENePGsNMwdfOSmagJX8pxXfE
7PF63BAsdg9arh++YDvH0HNtOOtlspqBllg20T17JSFbsiONFRHSjJB2Z8/IG8Y5HBbPsnsN6pDq
fp4f2ii1V51WNLRswIUIocHPYcatqbAE1qhQo7/z+Kkm12BF+V7xtZgQaY1q8p0+AW/86KJTSJBa
3h1sPgIg65hy51LoYsv3pwRJ890HUDa7SGZB1Du2tJWlg/07q15Udi45k3By9jEnUsob9GEH8YdV
g3a3Jg9FXymTvwxrzaKG5OxCi/QE+dh0qc+UUKWkEIBYPnuwcEFGTljhUxk31uZGC7i5Nez/fvrZ
uq6uu4d1o1etgtXvzAp+VXgi3CNPO0+v8g/rPZLBNc93gLRyKZwr2l4rZ5eEr6x/5gxxZPVFCnGb
O3iHhtUxvl9Vj8fWSUertJH3OAQpsybD8lKRYvhDCcDGKTyh/Txt7bEwoGXS5FqHf6IvCvYjMUXn
SfBHqFHLoMnpDf6SV4DLfmIxvIas9aTdKFlOR0BeWikwHy8GC9VCeuUcp5t/WF1ijkHAnCJQpcmf
n0kQaoerKwOPV/3mNDcPAqH5MoV/SV+1Tx8G38j7QmMPIv80Sl5EAfzEG9L95/INDjjgIgTfWyMX
x92242443/4W+ADDqkjiWnRpzXaaxUwT0BuaWj9huDtAPyropEL1tY3CgZ6RVXMkqqc7gMl9iQJk
luxps8cC9IrPIxU+QNay7nyRnifFFRGI9f6WA41n+h5aQXtRIzmA46dHbj2aXCc9U0LvD2m1uSQQ
zEM8eKYqFUvuq8Y74eieg+NPCjFxGHfDQNTlMlnSe9aX33MvOIqHcK31rplUBO9Vn7LBR7EFm4VQ
loDr07cWi+yrTWyORfc9P8fgq+3SRnxUukeezOREUAY84NXoAE7WpzrXVLKUGtlRX6FBI0Adzbkj
c235M82wuzYijCAuhnauFlIJA/bita3G4948aE2XmPl/XsS/P2rVa+7LwgzgcaDUiHzmnyUnaaZd
ntYzMi87pKCOtClNtlt/bxpYSv4gzoP+x4bzXgCA5dwVBIdRJAX7QWS99jKfWeOWOzi/GFrZhs44
E9FvBaNveIla8GbMHQqD8a+kl0S1Moz8CyYe9gHPzR8nSO4PLsjhuOJ9ZOYqv9hw7tOzfco0Be4e
XSzimtn/SLHNKAQVYPcOKKj1mVWUcL3GPtkZD3bYD2v65FCbyHTHaihrXvPBUX1HfM1/hJANzKDk
kgEYZ3mNuM36PPgVSCq++3gJYqlXfVndhHswgI2bDAeWibY4Dv8xF80S/H1JS1iULcj0xGc4Krur
wZACCa3BOpiEgZrbYhtq7OOrcE52aENp5OZc93SvBrupm1McpHFQ+XXDt7eluKzzizAOtXUbToyN
Vr8oFrV3p8DzZYtIxxYaJcmcNhf4LREoZehwi55Ipjs2yrvfvQcXbL1JcZb6yjdcm85IEX/mbTwV
1JMbnW3Fu9rODxs5CBkuE0LmdJZHlAR0S2uIFYR6WMr2qccrwowwg2tEuNzFEKHLUotPoeV8qS68
rBdXuueVuGBHttjRwI0eGIh88jTEk3dYWX61mogtpLDzh0av7iDT4/FePksPDHJ3wWkLYYLQ0WHc
uXdMScrwTZIIWbKu9jZD3sNTZYtp3nB7if//fBRU6yotmxuoTKMaYN1FwZY8IHcYraBkdYXhLnth
PW1SEh9itGGOuPzMSLZHgagah5Adb3TDtSi7U7oWp1zeycKkVRtFAq3BX0k1ezk5RkqdilbjQv+n
3S6UxOv+Ud7dsZL9pz6gJSvU2S7vx+FHMWYRPP6VhQYlOVAntH452RrRDNwDBJXEqOYGavcmK80v
Iwu3IDkUKzcr91DOOigl2WW7r+EEUgXIegoY0kJK6s7Le3mlUpLi56vYW4YTmvGONoRe+OPmIkA3
jH4eiwrizOHTaEQ2LQM7TozGXG0RsVdUCtaN0+C/fQrdBvoqKPx3SwFdyd5ZmcFmcsaoRuZ47nb6
9SrAZpA1YdTAso0e4BMJY+IEyUm/fBPKVK5dTIbheN6LPGu3efJeL5m5j6S5ixlsVKwXiOiVI+dz
T/bfmG27dHXowL8szG7p3ziQPoKYUxF1cBjR0oosPe1xpsnHh3b5MhHvFJVoBzkrukzqdrGEXvPc
aW8T+6Ms7Ogy8GKVNhrFkMdIFkaFjKdECHVG2RtxHu4gW4OaMjQjjSzVRT3WeChmuVT12NqrE7LZ
u7mdkTio5IsS92hj/Zn394+OJ1hKXKkoryri84jtfgKu6HePzYI8kaqIKsbKY9aNDXk3r/kizp0Q
h9udd1e/4kAQScC4/xqkXPZOCSGOWB5vn16Kg4pqQxyYGXjIEQG7KKgAXdGed914WbTsi5ynrQYN
W09gAL0Lh+yDJoq01+BQBV7GNSooAEsi5edNFaF2kPG27wLoM+MKxd67kHnzBJsuWUwXaAHDVxQy
/jZNK44rZmJ7FXtQ1utTwbmOa7iWF6jmTTbNuBpnPKon7FI4WE0z+kYEbzdy/pzs3b4XdVIHNkWb
PWEB6Yer8CYWl2hTlJ4sG1G3EtJMLTuvs32oNkbt9ICuqczP2cIhMKrvSqOykg2+1MRliLdKtOmi
YLMZdjNKo90RRkIs/mYUlfYzpgD0KQLjAVgQ9hizKaJF1iER592jw+B2y4GjVFFqQABQ+G43Z2pl
r9j7x9BVYokNB/55/FL7V/L1e1YZJfQ4JBaw1utJyKFv6npOTAPF3cYMU0pfeyEZ+0YiyIXwo02C
+lZhjZUEMh86iKYyRv47opGUGdFP+QzsSshGGVFyK/+y0RmZivtLI2b+dD9VXC8GL3mW0D0L52TA
JqgB5zVxvtuZUqJ1Fo8CjFiuhub0L/1KT+ARA3xMA5ZhhztFoTU/LQQUdgi4e+WCiDwEtv6ZYBgg
kiwVrYZX0SSRipL6WJItsyDAcxFZe0gRuTSQscg/AMSkIQpiqJLMk9MiZHOL3LD8gtTqlqMjbRnl
h4U0+I/I14RGI5OsEM1gQ20cpMkedye2y2mZd+39d3UZ6ZqnLVsJeV+LJ+JZ363d5wN+6hrTWfxh
ByTVn+/Nc1mGq00TTElb1WWeutggglYY+ZguAK2Q8CQwY9m20FI9qYTAKWnMRE9G7Pw9aZhQz5HL
vJ9aRLmRTaxOqu0Nf3UHEGYDXLkCHkah0Hs3YL28bycWazvGcjLrLqQOYK+uPIwAkq7t8vNy8TLr
9IPd9yXQDD2Dftao7tRw4OwPN63dUHjMgmiRvgvBp3gavJGAWc16KNgKoTvg24cGy5H+i/A3wlAk
1JscvGlFkTUfm07F5TD33A++tnF1yzSEL7Y6cQrpMBZgRIx1e4Nl4YzaCVE6oc7bIYr5K4OlDeKa
sWDYqmrgeGVXC/fxvCRcKCzGSbkQN1+V0G56EMNTjyTIsUmaRiya0omHu5c7cY6Ar/gFqVmbzdtR
8aV+vQ9sO5BLlDD0Hd2i6gA3Flg9ubqMa8JucotdpeLXQEb5kbYlhPi3ebHx6b5+sng6ZMtzW7Tf
k4qeWVhzUbwOO3blkBJGdb4NIfKrnJuL4GMTubXlUV1ukBkBI2t/4PGUFPUTh6637XGhH2QWK+e5
9aD0dcWG9h69P3XHgQYh0IjI7YtT4hAb4ceXr28lena6WqzLg6G7fjnDt1thv/S9aehX05v87xlK
ZT6wONJvmz8xdn/xI862b5oxTAbiagJi9Akz7hcyXF0kVK840U3DvwJJRGzTw2JY9z33M3TDYTOS
EVoZA0agYitYUNwE6VjRnJPyYuUboLWKwp4E5N6vjSJ8RM1fHZk35vkjxjmSZISOtPOCzz6PpaIt
TpOt6hwKFsIb2fwj+CAVGtSSwJr4wsBFQSXN3WYTN/UnoVgO+IMCYVdno7SjdnstvwzYkjf/aC9t
JvtRDctNKYQtVGAvQjeSfxsdJv3RcJiWV7VODjLMpR8J318RJXfXJRjLwnb4hoIqFtbp+bSc/T7j
LPpB098/zaVOBlXf+nqmA0zE7q/TDHcaERxxSO6ZwZdtFPahsQr7SAaA2XlARAQkJ+agIM76OVPY
Hb3hXbx1NQyz6eAP6Dob5EDipMHXTQiyyUk6ymGS2Saea4kl+c8vV4o65cmJyTBytsbou9tYUh4Z
N4Lz61tDGIxIIjt5ULIjLnKmCLFpjIoeomMF3gSps3dk5nj475OzWj6vBbRiqDe1vJ6zMPsRJh4x
nP3qpkkZ37OUG17noY6NDYT/+IRkJbCg+dSk2Q677ZeY7Y+Cl/EQnwHgWpv8ZWlj/XIs9ZGbPSPT
G+OsyFMunwZVqHehqQiaYQtK9q7TxScZpXbTYIaNoDqRcgYOesunb6x7kRwiVqCajD9WP+b6KV5m
EbylqzMzWCyWzeRIpIJxuYrj9MNZNQwGDINb2yAGtApc8BwgNFf98colcysYS4tGimQIw14pnNRG
ofspVhmwfHAwSLVVjyuFNAAjV0xOH85x0WWlcl8OAGDi1C7UC0Ax4hoprd5y9mBU0Uib2PmZOB+r
i+STubYlwLY1sK6lt3zhOewmSBfLqJouyseOxFpeQPFJyw/sfHyGf/KR155s0vZ6v0kw8rw9nH3e
VUL3eMkGyQor3b3Or8G/FTuptqvFTpSF5ta5DxZyFsHh8vGHzfgZE3XMGsa7H0jeaVjXcHtTm1QW
wn8Y7I15VA2nDT7UShEFkO6UvItwlxLxM257ItddbgPyRV32iFSE95uEjZ3dilXdC+bBIMcrxbQ1
NVgz3s88Lga+cLXwidXbblGOgGQLHPot91tn6JrRFVGSTOemwdwVHnDhzmtxkv9X94Q/B99AbnqW
/ochP8Dc2gK6t7nqvwQZ7MZFgfo5e6Cf5ZN7oQFuhNHV8oe1t8+cB5NJsLtou8yIRMxjTQSuTxUy
vHuWy1fpuVJMr7P2dyirS980ZrQYbqmUAznixrnpBH8gDi++gwX9lU5ujkjkWNy7/HNngIGlf/k9
C2Gm3jKmxeA4vrtapWXIAyyczWHPDOE9KK66oDEBiIxi1Pxj/mKTfrUHvsPBXATJqJOpMcmIIGPq
98ub6MuL6zq8yxQMhMPVShsMRakrT8UXLz9WimcCjP/E6P1tBGG+XFY6r1+Or9x/fApXOWgBrftU
OIDvGgldfmI6TPys+WPJIzRfVJG8vxoR67RsdhCZzt8WidSmgPu+iiESCxAqIvEoZIyf4e9dKFCC
mPZWmO6S1V1ze0CMhXXycZ+7kjueiIbQQHK9IU56yO57lY2iXQN5OSXASg3jsswBGBpN4F0ppS+v
07Pzt0Db2OJSXLBB+VZhRRPLLvNDtnf8Tb6CPDrHPya6fuMnM8/4pcILXd9tgZ3uCv3xp1g47Jxw
nF8tJr3whxGYkfrfeT4RJM0zAMIMhf/dVndWaT4ywLeJjiH7A528TpnDg9Y+wSRzgr7AuvIdvjPF
M80+rXNIjcKf2envevLtLlGs9Ko48luAA4qjldaigmS5+CMcOhlrhNZmD3u2bOa4x2xDUPHa9RK/
FtCmeyVyWyvdXMwmweT4+qHhcc0lNaCuuj3U2SPXTZsMRQ9g6lQ2j/xxi1yABFnkAAf16pKhdp6c
XjAcUThZXKqCGb50SliS+Hwj/z1xO/h36tyTRR+IuCWQqRaKVSEvv6TMXvXLMVe2eO5lhdcrzeN3
SDRI/9V0XrJpqPM4rENf69X0hCEsTKV1NQfH/3B70/y1cKUWPNdSz6kuwLRMjDzTlvfAd6NDktPt
hl0Rj7LEOufNvRxVHrtcoz3YFftdqwd11wslIRaph9t8hUxAeiJdviqDP3pq1fMCwgqCzujcXI71
HoikJrAyaxi75aUtoQvOEVmDe0Fit5DKg/VWNi4eNa/W/FByLAK9969z61CxraTIpt/lyDaqT8yj
ckTjDhNDHGYVDTcyIJUYULqszUtYUeWldHvbDFJ43xDT98nKp/TPG5cbK8ag5fjbNybFp+4KyNA4
hi4N7ZjUzvCiqSDq4IDZFNrIvL82OguIiRY1EErk0ZSMy0tyHYBMAS6JNraS9q1XWRDfVLtGmQ/N
vQj5+4jico3NuAyaHq+oiB0Ggqyor7+SHpy5unq+2gFl4vMqcWcX1D7IPumxqegeGHI99w+mGMoh
VCL8WHYLmgwK1TlU/4qnjFMmcmI3Z2tIitIYVzFeiq53/vZe6pXFXyRplyez+CbVwthMx8VJUCiA
JeIKVVSQQ/H+u7KTrxUpGyODEaq+GGZheUzizgFzIOR/RcW1rx3QrIFALo747Fs5vhV7rzEySO2X
j50aTZBP02gU9dFQeQF/vj7Mw2qHWuy8xHhr7JYgy4FVm3R057tbFhQjG61aEjIkhVV6ZssN8hm/
iH4WHKJNlhy9563pMfBH8InYxEY7r0jp9p6ZqlH/8LbFNJOf1hzpyGV4nbXGYCB9I7Vto1BiypaR
98XqyhZq5HmlkUChCKrpTB+V0QHwp1PlyjjWeq6EWJW5ENAHM9oH9FVk7MU0Sg9j4ikSbX/uIGhf
8Wa9BGsRaU9oVUk1nMyJ8dSPR/WDYCfxIylCcY9XIhvUkqs2W8WjEYejKHbPUD0kxOIBat+8AAa0
M6VTUCBPGZBMQKbd6O31IQVaLvOWJsm1Akh6uV6gNvbU+jB2S6P5SsxGkrLa7dt2TuU/r/ks1Nyy
Yg9HyNyiCrdoN0LHkah1bEatn3V7fFfQY0605gVZg0bzWiTlvpPXyuX2EfMjVqQaMf5W8eYAVZQ1
IBSjqH1orUlaTxtE18BUQrPKTGJHLJNfJHSaoklBr0XxzcXSBtWZwE9pv64d/zBW9FRHthxYc7Yv
V1ZWkbrkH+GY0SvK1Wdbv+3G9EbxFCPLfDN5N67l0G1dGg7Hcy438ZVmI0wMSCZ43drpqq0L5VQb
K69JiEXaq0JHStBF+8Ry/8we/5bgZbC4Vg/tj8metXEwfE9PeCuAU+7SuveAHfb9shQ6jfPzu4G6
Bhk8FiszDHihIr3Zfr0Ig3bGKRGlTRBI8HKQQrmxSrrbZB9JWj8WlkiDf21C5JYRxbGremaNfNLN
1/u3rmQl7P1PMqVQ8hKyv/JkqXU4ZfMqnqEdFXtZJCXCy4GIFnluxdcGviysdYaSgUS125nKfc3k
N/qdeTjZbmoOKC+roG5qaViOqlNZJ0rHGv1s9nQL7PNawe/pOTfjS9JafdBzw+bz0U6QozmKjEzR
GqluflWBnn53Akz2UVq8rhPw/qul4SBlJuLxQfYBlJHGRE4CIoygM7mrY6gkmfe580TLCKs5GaIV
UTM9MaemulqpdL266cTARk3Q3iTkbTs8NO+eMvI/cYGnwfGk/29iTZWDzLUwkO4mWW4A4NskCPfJ
3vw2djvCvHzjPB/TKk5dK/7nWSvlPI43NzbwlhbtwfIDSGOGCxdHgPqMe1C3FPBZwUmJMZbUhhmN
KrZairsYE+lM08+R9poANr3Sx8SiQyNcfe0Mj0ultJBMgkUFOkeAR8gd24kFOQBY0IDZXuMoT5bL
017KuC1+cIe6B8Hzb+WR4TZWAhKTKKvdtTO3O2a3lL32Gw2bS4QJ+Lq84rbrZY8Vd1Fd5d719wIM
QUU6VIg6PUvlp5u3p9qK7VMDry3hh+RPNrwoUmlG7bh3ogC6/VvcyvKSfKopVT79LkuwnoopStbV
15Ck2QBh/39LbY+9z1i0FdIQmL0fWD5ooydmOVNbDrxXm8YdInywNUoKSe/S8FeeloB4ve+zbsdx
laqTRUlwLyS/XXzLwCfpFcAGB6cujtQ37dq/i1GeETWwcj43PdB2dX6xZUjbiWlOq7PsWr6MGUPM
l163KTf1rgGDx8ePpq5bWCkFeyTOYuLV3qDdF5fCcS+7mUsGhhIyEhfjj+57pNHSdl1EmMWjfwjZ
JmZim6IRlaTSWPTezOBrvMYdLM6jAy0eE6jN5MZ7tkr6P+PoyxdpE3pErBOMFuW9BnMwNKRUEqeV
7p6mF+tNUQYqLdQOy5hm/OXRI0I7xOHlXySld5be2WbUgwxvQgHfniGjvhI/Lia5qXhXSQX+IFJf
pctaISUzBbCVf2gQP4dnTyyBXJxnY6G+jp6UR+fJ82HgyMFHoFntUHLFzKAADyE3fE/LRyvAiPFR
dla11q9LU2SK+oLghnFEAthSg7N6KcMK3oxfrHjBLztOPeJFD5ZIbe+SHEe1CRbhDphPPjG0KGla
LNmx1p6MKobPw4B2ENW2fYiXM2vGLCZ4oHZ4+sXHUVd6jh02MSGnGQnhgvZYXdbyREShdjVQjMgc
udo3gxfafgDNaE74nQRSFaaB15hLyZitG/mg2yIog0g2+FWGD4DigTJxvibbcURoX33P0yJ1IeIW
Mk+6vIQ3P/tTMdOhGTtFcznjeBPoPsM14TyA7wn7mXVuef7nxf0ytRjnNWXz0WjGb5NMPA381HRJ
cIlzO24ja9SdJ15DuL+UR5ce5rzMGDgxweVNNH0gLSr/t4pkA0ScFpIJVcB/OMym/yDIZLzVQqqP
zEM3DVD5fCAnqTG3B/mMXwWFUz5TQ8dHAEV02G+AElZt8DVLMidyOcOZ71ycsb/h3HOLrsajkh1z
FvZr7MgSdOH8lNCzu0I43bLpmeE84Sckvfg9XlW91OVGZ71sOQ+pK3TIpM8tmjwedAchzxZMFpUf
vgLKKUQoN+o52zY8I6XTMLSCW0np9ng/ZpaKUkp6KouMM6uFfz9j8kCuljakIK30kwXbaL8QWCnj
yty9XTzl8tgIJF6XdXr1hZcryBYWe7V9zYHjNB0IixEeVwYPrvWKlAvTwR3AH9GT3xBamUAbI5xv
t4XmVfvgrso6HVOVgqawWsfF5K6TeYD+GhFpahr+ivQWkuI+3IQg56/vaqyMiC+YpcZVQlX9FdLm
Rbmtlkx8d+Fr0B1n5Wfj/QfwWXmSyYPRsQNHTLSaJM80nzuYAlBYLEaF60puFtDDWmFWlFCW4yce
NPHzKiAXoBWr2UOd1Xnq5bOfKBNGIvngQcIBHzBlPDR3M0jjcdVtqzTA4Bt4x+YQEYYNW+giQ1Px
LK/zJ1UOBnZ6IyZsewNkRULvWcW7wzEyYvHY1TIXpDemeIICEseNaD9RO/1C4hXElQTKzSJbWFfb
VRDAlYWe3hXHdTUK+Z/qDM0wzECSL97YijU5RQDLQo/YYMiBKXIDWDgeL29aJE1LQcHXSMBnJ7tf
hOeEPlB7g7oEKR1yGapv5xOnzxZfYUllzs8+6dnJHUX08NmkVdxeUe7G2ZyCuNGLZmxbetqiYXMx
wpsTq22vGbKpjUDHl64/+B4e6nuW7JsZhfVJkGD844meiAGOP5hp27c9McjHi2Vt4UD36Y9fZnlX
ZQOtcWGZC2rrX+3l8JUHEZ8rgh3ZH+1EsvuXJ6j5HgIMKBPZhYmJIS90OOPNGlSsguTD96dO4HOw
MzxSJciwitxRCn0rx173MVzBZMFeFssPacane25T6uofQJiGT4RwheDiM4ClWGzGCBRnrgQUQWay
vzHh2A2BtTKc8fepB9LWwomt6eXnqRyi8gDhHc86cEuR4XaVbcNBVf51RzqENFjgYKGqYI2Cl24d
Rfq3lIM/d3/UFpOJLyEfQ6JVbHoAyWrdiinag7x6g8X/irIeidBlWyg6/VWKKm4C+3SPHA7ID5r3
sfBDiiQqa5zOiwxtC6paxdqsa8pfvSvw0ldG6xTTO2KK+snCRLyCkSPJsRlSbWchjJ6KUo0NNBvp
JLtyCG0CSZS7qzpAfsHL2UXWQ4TpnmU7Sf3tQ5AdNSNZsBLCzr6loDtYhaxp61Zyo7lw0S7RkS5f
JEhUsScIZC8rXcjsqFtZm1Skk8YvhG3NOEiKt7gB2t1O+vHmuPN2qAUUR7CW9YB5EmpG9OifTW10
E0hp0X2pbtDV+CP8VcE9YpjiFTJ+jXFQqSzc0Rf/+9H4dNHAUmf1Z6gkNBWxcO+AlvarEs3Zb2H2
e36m72hWneu4JzNqbX/AO6KniY1Svn/4VrzYLyA+HU90FDVxnQZHYcAfs+2sLv+bAJNPTk+qslA+
LigoVjQFumHGasozIKLKBC6JQKVppjoD754WXlE2CbEoozd2V9GBiD0xEVFRCi5W9FKptc9NiJCZ
mByonyGw7lOO4hEID7gxS04rOP2x43HX7x9Hyw+WdHmilUvOSzHamQS5ex3MfOXskUuzYQEINFRf
PQMetznM4zBrq+IfZ79yq56et7yw4GqOQ7ZGWdpWllVqcAnw8Cmhb9wyYxbQFGWxSQfYKtGhsdsJ
5222G+tMmgVIfgsLCMuFebGT5Ozzqr/RvlErCvL2lbhu6T2HHWspQd+b54VAx3pKu0AGabQrgI7p
Tojnfxm4vNY/ZUzM1gk7yRCC+c3Yhrxfo4Ow+XZy6HoSe2IBbkuMC3ArfN2gfvltb5awv81YpJ2p
Q9Ta464DrlPl/NUnbpLq6CyEkgJ4nFeGlrE+4b6a1AGRZ92hOws4d44lKxZP54NQve1sB1X73bdm
rWDmqU27geMtSslGERg2Pb6Q7jdTxRRKeNTsgH0UI1NQNQdrHteKS3/RPRxLIUjfqjSD1VlNnS11
Tlu4603rhZjBeijqzJ1kwsyvS6eZtMy4mWgmBI+2XAQdbzff+vjpsilte38L5zTv1bbBoMjM6Dg7
r1nenzQsPnx4lxqhpx5zRdtBBsz005lesM32k5ifBvBsQSx3pSUpV7Ai+pZr/829XLX6Y3M570aS
49dwzK/ro9Gt67fD03qe5n79/awEs3VIacnDv3nC38pqzBuvCDV9czM+bI97Y0rOUplH8TH3rnQa
PJsehpNwa9sDTcBcDmoxQB+q80XtjTrUxuC8x9R6y6bMIsMYodqdR1zuFyeGo5rZ+HQId0t4wEkB
TE/4Mr+vw2mbVi1T1w+ySL0sKwMnvMp7ckHw8OgsUIlkUA9Ye/XiSl/qSio6YsQvzOXq6Y1BUV+5
yo7YQvMuRJB7oplVQfEK4hmbHDQaZU+X8slhIVupSh2d6gDQK/4H4h0hhWi7mpIn7uZPOxjAM5RT
CMV5RjyB+V/9z+XQOpDV3EP115a6AaRVqUs8SIiO/H0Hup/xan2kQYF33nqlFy82UgUM3SgIXVSP
+k30aEZNT/CGTsGsrSZ1FhDpH9MMH9VXX+7IOGhO5XB+4DI7J5zgs4VJaOiINuYTFjIoafgqq1G3
BiQfHqLYqoa7iJd5WTdR/Fy2IY/rHOyqB4O7HHvqGsmB2NOqUAwyFp0SbJMfq/vCseWMo5qJ8fjv
5fw4EsSLi8CyE6Ye0MEgOIr/lbnyzU3q5uvHDvayNq+5sicBTU8RI/2Mgq+iw/w/5ENEhGuSI83n
Dz0mgwPzEOfhbGRG2xugSAjHYD+WGE7o4nqIf9e9qcF+1oGP0qhWXA2YDdsXzoFQPsvoACduXoUo
IfaQyOdri/3DhZCV3ynLVPTcT35tE8Koblvi/GcAvj6JIaS+70zq/Y00XU2aGPwZcViHZQ3WKX8p
FnER2rqukEQoYd5Nh1DZRLRcqqWfrRh+pUY52Ru1TQvioImYdNqnP5vftmZ19L5QDbLfZ2RSzycc
cFykWZx5NlAXcvCJFSTcnESRz0tQBtfoVVSRqjWiGVOflOuiUza1Qr0nkEo76P9c0i/mveyVz9fw
xocBAoLaIxr6vQxGwMu3kuCZEnyXLfetP8S18EARIhWS5hQ6AU/3u1ggFYORb2J/ifrWFTwm/Nmk
9wRwWcNXMgSJ+vZkS2+0xsgCRlkJwFgBwVxLcB5vQp/Fc/7kIkLGY7djfEW7YPUuciZIemImrcE4
czDNPKoMW/BpAeR8Dv5ApFo0kygC8S72OfqMxFPICiJOZutPyPwyat4Q9SvwsSOCLwYZTxJVv02z
43nxLQvLKs5pieiGDH9U9NVK3mcGdeExbjNjVYkeBf5OBYh3vn+jYCMbzrna7HO78CIUHleCrquT
5tt9Ybf3r+xa/r13mz/3hGspPkSkzOcOR1y+KTkpNIjZQxytYxOBr6D+OMagktoWiq8FwLamoGJ1
GLBpo3raikX79S4Xby0gKEk5Upi4utRMztzpFFJPIRDQFmDb0aukjRYvWalecuJx2PL0Bxf6z1xP
yifZz9SOUoM4XB0+fPKXXlqOEcrW8yZSpGdGsz7c3doPJmYkzAkBYsHDblNuqB9zgW0QM0O+ubHS
rogJPkgeC2incb6IRQYOFkPJz7rUj0Al8+JOKW6hEYN5nAn2NvKp0qpm9xnky0IIaziCIa/VIb/2
RlBATBfFrCKwC+TnSLZYjGn1UWMN0WreQ9VXizidyRknLro2EOtwvxeXaBicXCCXZWet0Iv4wDNp
9e8hPF3HevD8jbWtcXitK78ttjwXKpPqgsNc1SOxsbgFxc3UIR/AaZPCsUzFOG3fP7oDp/zIj6wa
fS0PQFSz6jI0oFPriM8uaAxeWl1cpxTtmPRUnTEjjbRdG8hECqxEoavBpBZ7xUaod8KcxdsFPk05
q+DSitXkNoahZv1feeUZkcVONlsdmb7RFRTEhwBxrePBieiQQTMhKVggtgWHFup8O0RFsXouTEiF
prZ6x3j1zdui9HKHPmSJJ1ZUO+8k0/mgTsO/pBDepJVh2das35Lw635dvM/X29p8JoNxC2C+n4X5
5Fne5/86ZcYmdBRrVuteDHBHVS+IHAmEoW7TiABLN/CABUTdI4ZHxB/J81JPJWncldIIAAAL8Yo1
Q89DaNA1y6PgkHA2sRKuwAyNDbZimWwXu1A1TKrictmplUz/76N/fNM2RDJqsXEFaZcSh+fcI5cC
JuCWfaxAD/fikHkVrbRksd6TAeKmRyCk8vLO8MN2Q8aHxWDEDv4DMJ7GgehBgY8OdbNbFJkxyXEq
/L/Gv4tMwpC8N1DAYq+a8QTtlqZlfvJf4XtwrC+tASb/ZqcvcmY3+PBRe/B5zayaqxp2s0Kf+flk
OJrD8wODL5lv3PvzivZ+x39P6phPoz71oIPLFoFwtQt4ZXpS2ctGxjq8wIpJw4fbdz3KAzyNbSvi
a0OJ01eHpdYjK3bgKl4iUwbD8ZUGCgpwtrnvdNHGs+PJGaEBVkfkrzZNeMcL46TQX++IEv+IEk/Q
7B9CuHwThycHJISy8HuCBVK7NcQ4L98nH2tQwMmRqTqnaxgftZz2XxRSG/OFRDMoSiZdt2sk8bXd
K2NYiW9hbYuR8J8NiBA65UcafwPyWZL+9XXvIJv3elR+QJAB49ivG9Jh8mJDTqy3GfIY4cgSDARr
k19nq4RxB+J5N2p9+4XSfx7abqaDgFvg8TkUzVJEawbD7pGvt2zIHSCdEyriDJOBdDHcMKIyTJ/R
tYgGs+2RZbV5y9A+pHAOdgmPpF5Aq4ywzxiTFkzARKz66FmDrB8r+H7azeI4tiSgrq0wOXuAa7rx
W3b+BtW18XgGoigyBJnDrfGqaWtjixGWPrFTmjHFIC7hNPe360bHNAX6o17QTFYwn1q2jm0ydXNo
1UsqfkSH44HRoKAdsXVrVuXGpNxs+SaPxbFs7PzTXc1S+uPxI051EkMKp9cPRrkCHSqGuP3N+VxZ
jXs2MERLOcs2VfKRv8O1f/IqPj7ycqEZdkdfDjQN//Yxh0d9RBQlSm+pjiK1xWIMKOFd00Q2Bx8t
O4x0Ve//nRwcp4OIbq2n8et0eXb0vDnvO+AAjU7LaNsbs4iIUoh8OupROjuhAffzzqcbovmald1h
VpUIa5BqapCGrADtV4hC40gPePMQx1Dou18MfCKe4LEIJILOcdXPufswa51cx0neEuk1QlYJ/olp
p61/wvY72mHk0+flHiJ7x3U58SpRDrOeRKj7QWsaws0RndwH51Ee+R06Ey3lt683qmyKT1YBx4Me
zDcRJBDWL4rI52zDDUFkMMuRHB+v0+NS6dNzoeVcYfayJdCnEvxOn8eUmy4QJIa0rhj4w101mbzw
Xhpeta/VtVeypzNaw4WlGQ5FknFpvZ9s89Ude6fvF8+ESJ64/KK6PjvNzkl0PrGlfczWJeDpVUKu
g+acNzIRClqNlecVcG4CxvMniovzYH3R/HYpTKqWNQkYK0js7K0dGfMZW8B+tOkOsgMDrvl6klBK
eU8H8Z0hZ+4VafLloyTJ1m8DmRfHyJaTXIaiAt1uHFdJk+/eeZtPgnq9r1v7vaYWxy4mh9U36svU
hegoP5CcIkyuyR0item+kp5NHj6iOztx4r9okG/C/e+Jvm1nsUnpXcC3kvdAJqBg3ai4OQ1LhDpu
tsD2D3kD4mBrGrHY6HygF9mNDvemEmu9e+Z30jj5CR6Ih+u4DikyLMVmlqj+fY40TMmdwG9Z5nuu
uPUB4HlelRO0vBTDjZvMv30m1P7UHBnaaavSVXp92GN56zOMD1Vf7j3gcP79gFNn5LZq/f1V9U8e
Ho8wG5oq//tMr++pOo6XOejIvXKyBaE+GUbwiES+pnHL0YOjikjWTKTQ6VbIiCAT16ndUWwQeCnF
bU2yOV39LDVLpvVvvnLg4DmVUHM3CC2JddwL1H5kOtxKWG3/AsEybjXwbdcE6Clp1SIYpx3lETu8
GLp4mHAwdxmU9dsIEZpGRY4FlL1TJApWdt3nI5ZAHkg9rGeSY+E+YQvyd+H2iFD6ZUGwmn/7aLR0
XdL49qAYpL73AS3Kn3NUU/nX32vxFR0qN1dKMS8kO/xCN6Dl7FD5d2/3x9hsgH5xrY+TbHaxvNZ6
McfHyr6d66Y0dUOuR/8WImSpMGNp3KMgekx60TkT137xuv9e8uGRYLFvfWMPkRYKmkW49IKSLFXo
W+uwksym5YZhmomOh15VfM7KXQ+csodYVkoaFauwraFL8a6iQl4bsWzpIDwM5iHF8IhVzjvLHcto
CzkcGG95DvKdWJlPV0l70RYvDt4bA/hFG6zpJIQPnj2FjmOUyP2DBUj3F06hBNSGhovUwPp2jbaP
bCL6o2Q5CqP6Dgia4utMvwT/rqxDlVCuMkz0tS79CoUFEmwj3GwZzKpAx0RnQBVSird2Tbct8DSb
hBOwfzmLOtz5p60/GV9P5rNaMBIGixJLwUeVvXJqd2Lbu+nXh+oU2TOK3YOxr372/ahGRAeBoX5v
h850dBhEiLioTDQfZLGSNrKCfTJ2Hlvo3elKg+ibHgetNRKPyFHKpuqtvWi2PCwH8igujuhngYnE
D+jZiKzAmXyS4cCN/z/z2y+Mw4fmG8Ge9G3KL8i0PNbYWAhduQtbaOvVhzqG3ItktHURIW9nxWGD
BMICZ9jVZi2k3/7+Arg1sNy2RXv4G1AqWXQo54qLFtYu8P/S+W99odPNYPSW3Af6sz3p0R+r8U9m
gzEu0l2QEUPk444S218PMvy2AWks3qv/fC0+C+2hmQhU/iJ/8L9pRUla6t9k4RmSXA8U/cbeAwik
iqpiEwRTp0uuQn7jo9F7IfoO9vt+9ziGNew8oOY7Xag3pes8ix7M9RrXGyR9mGLqm4EGbt8/winn
mcUggvHIyScmZAXJfYJhL3xVVObrXm+MlXSd5n2VShw9spDx6zUBddLFix8K/HMoI+qc2PDevYMi
tk8SviGX0GebMD50+Pl/K+7FyDtjGD2jSm3p3yplGi8OYybmfGvGhT96Tt+/iK7IKMVJDw9zwJqF
+mLGWQY7fZ5oedrdLlk/8NylKR9vVjfe4B5MRoR4dha9zuE/Q+gdMK+KdmDEKGW6nf4yPW4nwTl1
PIi4rzG5rKyhg8nkTpc/VWG1sK/cJI8rEIKNLE0FEPKaRFfvoIMP4QsL0jnv5L8LVym6cXRt19sJ
eqXHWJs+e9v6K04pT9k7bbeiDvGf5HRsP6ixW2WcRUxqIuaTZnbNU8M02qvaSXY5xAznBG5hv/NE
lpUKj4/8zMjmiLJToN1u87GyOSFKJcu3bbgLMOCu0Z1ZAW0Ktf/PMZNRLqGM0hGt+PhfaYlLjrTv
pq7f1pWHcLaEot95kEJx3p3yR5vptbimKnE9EMV9Sp/LzAif+xkKZ1XpL/fy0p4ydTehRRFJ2Con
Sl76XPLJvJDSts2yZVxZUZCXd6E3YkbDHtRqjiRfUx8fG+hz7caoVKxHfUy4PnxJAr05v3B7PlNn
F5JSf6qrEJTaTM4eQhvfDOcVcfh2mKJoRE65FQThS6GUiLd3oz0SCCZe97codSo1OHt7jrzU3hq/
5Yjm9mdiSCxHI8darGEH+MI+dlQdw9zUNpgFEmwFSlz20HAdlPBgIivED8Zqkvm1GXm92W583Qxd
nrrFTGvxkFT51au6obQRQqw82GAR6dM/uYIbii/ea1IaYC/plFbI2jmk7ru5fPKx6ZeC4ZufT/WO
b4VndTVOBPxeMj9Msvth5O9cEI8GuSQwxes/ZP4VxgeLS1l3OXetbwHV5wWjBirBHzCQHBebGcRt
ADLdNvBS86CiUfJU67u9pUron3gH7JeYH8/5P1jVE/ikACnCpR5FW9BsGSwqQV8jxxhfFBSu8HIj
GG/zVff+n74oJkR2BMzJq6P0H34wvQFwrIqwaV3jrNYujrFLkTFDiHGG4Jp67qJ/QAL8n6WhZ7uT
7sOM6H8yO6630PrpOW0HDDjVE3wptpnXRY9pzF2Y+XV851JjRuek4MJnTE4aJe4fT5X+JF/4xD4+
wm+Y1NU2BS6iPiIU9byuCIEGDrjVJLKcgSxzAcZJvfdUO+iUalC3adVNHgx0hFk5PBQKSK057nYH
ws/udGP2XS4QcCeImrIeG2fD/0QNLruO9xVg3TaafCSkLEck1oPi+Y+OO4tWXgUf6pvT3+dKYcIr
KjurCuc+TXjnXQfDXwI/zdReYSiWqX7rFNR20cA5GFcf8CSa1kbjEt8nxwee2RK9l3cVYfNtYk8x
pp6jzb4RwjCPe3+nxpBS9UsfdzkX4Pp+T7yGb8Z7n4lSNiBtsn4t8fb9ExYqJ1KpUhkL3RxQq7Ev
fw75GR283VryEklY1IrRpho1SPe/hPpX1rxEk+WGkPehNm8KPGVm54FFnY7bYdp0cOttaXsBzFBZ
KyLy2+zZBr5KDjay92yglWc1zlokjcqQ09JvYNFR5N5fwbm7mET3uxeDyNwJjm60HWPZ1P6ripll
YMYNHWNkvy4/jKIJykjekbXhR2n/czGAqpRIxHZj+4aWF8tRi07M7A/uC2TQ1njbAZSb29WZ9mmq
tlX7WrMSe5NTn9UBSo9OoEOgsRpFO5jhG9kqtKTkm3adQWvoXUybGEmgD/zfl/CpU/kqEkKia9+3
oTJvl/krAT8sV4NSm8qyiflYbsVTA9d1A9l5GxYny3Sb+LF+2lFiGE9WTD+ZGPYkxV9RWZXwYvy1
f1mK9i2BHooA9cIcrKPf1XY93ieG9kVsUnfkDFyotheTJlEdXyMR7J+h0JvE3UaMlj4DXfiu8yN8
s1BSY/oA1pNvEuYY3VzjqdFKwGBePHD0LUvp9qjalfAMdnpMvaDwKMW67KAZ8x6RKMm5toCTXXu0
VFrehtH9ER9hpq6YlaPq4+rGvHvbCyofJVFrp7WVucRmpEcCSrOXXpQTzZkOGF5OdaX6HP0UGsWK
KyFP6278YF2/E359Y0SE7GP0a08lT00fHqma7KY6b1T/Q2snF8jlNYvpSwkG8y1P2M0izZU5rvup
dayADGMhwMKUORTMx/R+gOyDRHDTERrSl1N/upJ4IVl1Sqfyt8Ogq3l0iTdX5OEfJPAwUMfGuX8W
XfkOQXwCcBvkin48EJOjg7bp+86yrxyU0d4htXGQOIsJnGNo1W/InvUs1WfiV0EluY5Lv/l+JolD
MC9jBwDUXaxRleRbn5uY9Enr1isvMPOw0Orp5/XBnDYE7jFb9Wza9M7EgvB4WNDow63yjvFEfXQa
g7zerlCiUGiBboLTX3H0meHYfUkvQ5jqRW/fy6EJSwwOJgViF0b7ACdRiT2qaru0yaZtqzUEzIHm
jTFeui6B6L1JXjzMKWYREBCeFtRZ8q+EPJuohXvSrcj/9gsfNnzDCvukZhTpqeKyiLuHhLtxEadb
bYwyyrA0PuNeS30mTIbEn9xVAlrvyJDogy33C7IZaUTkM6280BarXBwCYLUamJMko2752rGSw6Vx
z8QcSo97UOdNDYZ5yQHECOTq2xC2vwYZcUn5hXNB9fXjcEgQaHIO7EsUYlUKhox4efceoNIdlnJ0
ToZLnp1SGVlfXmc1ih2svjCUAwWrJJ25B/qC2eRLezLhQGhj617BIAZfgwEmFo7TPsz2RugshWEQ
l3aUKypN7OnvfZvhXwhuAnw4/Ip5C9KzD5pxMOfGZVHceqkx11696C8JLoxLkihYWsudOboesy+d
9YdJkPs3Jb89WOGSujL0yUkqINMOttX1NhWwIqmHZMDgpmodQJcALDlI4fFPBmG5nKZYCmc4Nnz2
R2A6uyATwB79WDXYQvYzyTYD7CEb7NoxXAC9+BIsKlBJFd6sEIEEoPEhPYqlmyd1W2/n0AXWVeGs
YPaWgJMt4hqejOs2X02OY2ynAuF54qLvjg2vxRZ3AvEyaEaNi2jwSl2C9Jlv4Un9gIrm1bmrgsm2
iXtkMq3Jdf22M1QvX2h/NvfDsKnp9Q8Q299WEDj9HK0ieBF+OZSQkL7sIezcpTxzaVFbVT6VOdhZ
4xV5KMx3hQrF8Kfa465Rz7X+nrtYV2PRjJFcpY3skjNkhJC/1THov4EeNfpJ9folXjN+spV3ky0t
WZqRcIu5HYnWi800hwPSSecaH3sG1//0LQoK8/WRVUUyFkr/dnk1To4DuRlvTOxXTdiludWEBhYR
3a/rYVcFiYrVdXbln5cZOwDbUvrx81iTNJwdKZs+r6TKB2hDJsvz73tlX6NLa3ee40TaI76Ser2C
uUF50Uk6/9NmJuBi5tCDvqtNHQQbu080FhtgF+E5g+95dglI/4ygBbsDE1z5iUB2f2TZLgagNnch
JJGTTqktUQ/PSViYKjz5zEaGVK6gWcP96R8UvrS6ynlRcOSlUy37vByqflxlxNRhBRGsrOMwXYZl
e3ShnTmvApCpl672drH1lGEbK6x+z06XorAd4vp51jJz6A0TU82KZR7OWzwo78dmT1YgWW9xHHE7
D4cYKLWx4wDepsDygN2M7vrO0flLIwK7fRNtBmV99gbcqflLfnV6dggtmaEt71RgYhMQDUYfpHw1
M1yCgmLY1Vs372yyLwP9VIy5rG7goGpUfgE6aI9jkuUm6Rs+awEMiW3k7CDXZiHU8AvpqSnknWU6
e7EkaThyHqUlVEWIwIkYeCq3kCA2AtARcGxcU9pXl9VglNlN7JT4cyNEDMW8AAvRWky2Lcc9F7NV
z4k7yLNf/4cwmHhsSLBRhJ+rk5wysurFvVxYdHQiKPl5ESL2LqVLTEiPeRLFbO8J6n7D0IZpVeRY
jZmeYODVbfBo5oEE/SxoXLQXniV9ELWgbjQgZHYfqBda/i/XvPrmnkihH/7XsJcS/Or6QMHtzIbH
Ks5h9m5Ko1o+s8f48MGerf/66rH9yxOy4bvG4rLxkIb+UCbRQbVj83f3wS7aWQVqRPFZOKmMzsYO
qqRIdCYQOkx0Lsfn6UY3O+vrx8vo8pbkiEAuiZxRU9mupla1JmVhvQH6MoXpsCQnEcMi+8x5znCc
4K6/t0v5NOkCmlIL7p2REfL3xxws3HUkU61d6/2noh/DqYHH+yQiNhDnpo4jvHWbsiKtvdvpRA7x
UfS3fNluckuDXcVwh4AxVJSanoC76yCM9jr+XG7CenP5JcYpjD24ypmR0zV16jY9XDF3H0SXfMJx
13n8zXdR/kmv688cmXj2hUhUhqAjaHI7gYm15E6C+41gow5X06HbQ1lPcQrfR1SarjzUc6zqw36g
yFf/XRK6epFO+zI+eHGJU/9kQgsHFCm7AtsWGn9lFLIRcfXwAbqHrnweKcVOKPiqrs5qdFCUeC9p
lmCEXR+S+HUZ95lykB9ju6EzVGlFJ4S/xesyW1t3YioC1i0SLDJ05diTC+aHGg2OVUfMCQ9XirHy
YPMlBF0i6zXCiupqoa/mjQ9TNvyjWE+4judgnotV662Uf98Lk/0HNMb+Nufjnxp+9w2EuHb0ZGS7
z1NYkF1r7zdMBiyi2xZCKZB0xXBz2uySfPO3/DicPB0WIUIChyMy5G6YeqcWy17SEqAcnVjc8cJ9
ITghT5G3sIe5fzKcMuL6Y0gEYOlCmrd2PeWVMTf8CnuUZfZLKL1i2mhkpOYQ9tmeeCfchaV43GRi
LRo2CAI4nL8ysFvwjXyQ1PONFXDDUQIOu1H74Fl6CJeYfMroDHxUZtz3L9leMzITB1cs58NtkfJN
8cxO0PG/i13Nu4Qosv/SssU8hC6UcwGRXqq6r5/Y/rgUeZZD0CqN1/acUVoK2lGauALJgTu9/IvF
sXa/pPmY6sLolr3Qy/nyP42esNMGYlmhbYiDoOZfzHNzbkxp++aS68FTKaBTlmXi8ZWDxA1t6+pT
+C3+eTcvmPnENx/9pvpVhADoz5y2wkgMeUXWZ4MC8tCrXfevKimMV/+exHxti8fk84WYOxY/TB2w
2gvsKBmAwL4UhmNnp4xRP5smIUmB3TVx3LKT//UWMeRYhKfVvyXilAZCUnDecOI+P4Nkx4ZNWmOS
vRJSxvLST+Per/WgwH+zwj5IuqDncUq5dxlovslzb3/R0wK1lSjAXQSEcH682tkd8ZdEpx4vu1Zf
TpNgfNOPrqMoxP/wORBAq+LkcwOY1twchUcF/YMUheeRr0zwJyV7AW2PmtZjY9e6mlM/ep0dvlkN
Pma1/QNOj/JcR4niYfWLC8cigWXOz1aThLGALLlRXyFSO/vydZGJ36qnYJJ1INiLLaR85jdNkjRO
qy8JGs70QTb+/RhACsMu1D19AZOmADRWy7+8fIwOORUl+fUkINuWrlyQsGCZfKDb764i/q159rnJ
0UQG0W9olET44AymgyRUmOLTwrmxQvUdFF+DE+ZgLD9czkacOsIElH1JudsR4aupGC5UFPZ1uyxX
JxLMpLxseZdgc6Ate3w3lHaD36w3rN9vBiHCGluNKncCWuUvPvvDi7zFZuWK2e9RoKigJIojw5KT
wBB7oMcf+vlrpbQiAsOni2YYuRSdgaLbDvqdBgq/oc18u3LHRd/m21rg/0hxtHiw4Gom3Dzhd6se
tPTE7f7SHZe6uLaVYRSiAKS8WZRGemD8JEdFQLfxlc/KUA/DtjM49f6FydHdIVnZAkHYx/Yp32eq
/cigmnKWTSvGWFsR1kpf3V3Nxafy/gTYt+JLFq6jXLjurJu4f+/L9X1r4sQ3+gWN0zIq7LqayMdd
J1qgfDvrFvzC46OYUEnuCM2p/oq6rVrfaFABSYRKI0haGuNNiDXTH+Xi2d6a1sTkR4uWhjpSmeNs
3WNYlXmri8Xz6HJlO6l+zFvmEuD8zjTMWFqOVz6+JkEXBQw6CcOtqc02Y50j55RerdrLMLGcn70v
0I/wKYQALCSeyeMQ8oFJ2EnjZ4s9KXGJtNt/vswnGFr0PCwccso5ypDYWAizzH+0JTbtDIRa5Xs1
allVwYqAa2DvvmVlEB7Yc1xuR4ECn0Jn6LT9XB79mOHfWWuNLFtK09NXKTKBTChiNSVl0jX+4jng
MELMdlQQ0xbhYL3KDlGfQMdwiSJeu39KnpNHJIRAORHPoHqQbTD73L9Z5e6T5VOOiaGA1n0LCl6Z
vHBf+ccfa3yzgIo/D6pw9Qu90MKMR4sjey1oqT8X/9evHvuczsmNiAQzMdMaaErBpJWPhNJzd9Eq
sHARfzAdMBhXP7UG3Ahy/PcD86TcH9cJnEPOlEHZ/VSLhuVHghZrHpRMbDHXeH1ey6eSBYUWDVZR
e8Apex816g4QdQzVtjwpN5N7v59oFTXcBTeWNu10zSrWEaMJb7APEs7Lqf56gNB1J+nV0ttFnafA
ggwOH5KmLQjV8kGyzyBw5L1NVsv9EFLl+/1ew79o7EEg1jY5DmETIBDLu8S+N7e5ghvLJOUkUzbq
SiM9dPO6ZGb+HchBsf2011vc9moEgkUV8hpN/Q+bbxjPykvarFoLPZyyq+h6osrWuYrhXkLgm2IY
9PQ9b+LcoDqqAaw1coainMLCkH8/FHpcvpNsIsK+PjlIqWio44IvuY4Se/ZAmwXuR1rHMoHQJZvg
Tjk9j27x6LvvjVsKWWzeEbZhGM6p9Nk+CkBL+8jTbVUlsquHh99UIrZkeCD4uaCesEZhSyev8kzg
E9O8yrkxO+Hoai6jjgVRcDauZEcEPAQ4YMblu62QWZdVxGcVTZmSDLHHNLSzD/yFIviGQtB2OkES
EtLwbPzuGrZE5/vgUqrt6AWd5Wbsn8DAVHyNdKRMumkdRNU/hFjMLph7UgP5Rf1233TJMXjdehUU
YNyHEMyDZTtTMamADObihwDkHmAAIN+NSwRzpFLZoZGRpfTMDMoaSMEyuFLUTrx03Zr4KM+D8FF7
ko/TWlVpkI1Vt81gUbd0H/OGEhjcZH3JkmjKQTSV7eudKxjS+ua8nu/rui44Tty24FeO69JvA2kg
7LfcLPvx2Tpv4z0mfi5ud0rywEzNw4yJkrm3fMSSZjV4yz4uxS+IqZr/J9qrXKkJm6wbEIOkwwfq
+hunuUdVtOuJqHYxdbVXEgTCc7V7Wygd6k5ENV3cEdWeFUMQibrXI+HpscRKeVS0iKIVFqcTXJQG
7ZjWtABznzjpTCPTCHRdDofQDvpxxCXdTNUUadp+kKF1GmqXtG55WdBmuzkQHA+1NjADt99QXv/8
Bfxe+DDsKa8G/wE6uxKQmy10B03CEgjWIV10uw2IO88tebnmO4hk6SnpZs/3D1ZTVHXr5BXoXVz5
j9jSqYBr56Gh5HmjxyRDJ/nlHpEb4CwU2artqEor2r1NpdfWAg6GWnqXohTO/VnOPEDIbeoOBNVx
IyGe/MSK1lP7erXd4N1ZILJjbFQsZJJtR5D9kImok8G2BD3NSolI2C+ZFd02rtcQ0V3YCeojilGK
8j1qKy8l+SHza4CJys7OPC1Sd8821AtJFWT4ayeCkQ8Zz2Vj9DufMOj2ViEKdBP1mpTxhMDhhUnq
qvu6gQBlMTv5jFBdrmbHK21Ck3gYLgoJNVEsyBAeRxPgwk29LuKL97f8v7d0VkkYd25f2Auo5JLr
KZ5YpvM40eKsgoBGhS54YWzK0Py/v+I1dd3SFH/Dm3fEe528Moi3yEI5E2rdHXyPI7iB5cHwKy16
aluAXDfCebvUWPCfSH0DanLiLeUKGz/PFbaVIQcavLkakRQyP5Cj9OcYbHi6j+PVnkHOtAaZ3glC
2kjr/CIeomwIa6Q3Lyjuh9ugf2xEmDPQrPD7xQCP7tztHVNse+wuIpcz8sYWo6PufuKpq6OZVsUC
JYm2P1RmW7YzEAv6nz0v25Tl4OPL3qwJYJMURGaaNKGDxFmAKJfrVaPITEhT6/ByRQ1WhhVPMsfX
TjGxkp3pcgq5x4KDKB9vYZ4pS3EnqbGk/zXNbcZUqBIBAHI0WRi68ejeyT/QvzAFRlt+9OIZep9k
PcV3nldEFRU+vpr8mBw+y/runsNdIaGzTB5pBvHVQLuSb2O6yiIJD9HlQSNV3Qv55O+tqYJz6VJZ
2vK+1x+i3u7/mqgiR2XuCTR7wZEPAqJS7P+lsL50xYf7BTPHHxCiS0bCOdSw22O92jmrGpzVtxbF
MSzpQpMC4vHY68ld6DUekfM4fRtALEHDEmS6S6axw7fEa2dBsPPhXE5lvraBaJIwfxYqAh2x9rPv
NOQKOlz0a+VQKxNwNkqznVGlyvOp4O2dQdPOAnbmE9+rsDFJI24SrNkFrMRmnndIb9TiKXQhiyRr
6UHrhcJMPxHwXSajyAEjT8tPRiIQjF7dSSgKfTqu0qGxCveI7uK0UetwvHl4FgowCvoHyOhQVzBQ
jeNga01Pw5nIhMfsSBhspzV6vjlJX9bNEGtjaQAmrMpAw4biYSF5h2YKbOmOs1f3Cn+OuP4ZUX68
W/LC72Qs459RSCNz0/Yy8GryMg13pu1+54vnMbBo2y6QJ6g5ctn/PXMS25xhhkkyS3H6hzUbQUfn
LrzOoGqlE5Nx0oX3q3fVVpAxgfVS/Fena8YM30EaI0pRh0o/O2XhpflzkjTbtTOmHaMI6fA8ai8g
irTVXrhHz0yEoeu5ZYnUG/P9ugJyjecwpOd2nPmW76Q3x7B1c+hWOe3Hw+ZZFEepOcKrArNINp2d
oEGekBRdR25y9H5Z8LoopvdwIka6oU8nwzizvBQMzyWdC7fDqf66dbMs5u4/jQ5VIXLswdoxT1O1
6YRjPEVlP3goe7XwAyk/hDbcLKiNvRHAO7bz1jJ6nRNqrmY1jh5CeSLVFusWQUArarWRBrO/0wzU
ESh9ia0SqpmvyR7MARQ5ipqO3qtW+VV6maiSrqCplJTAIL/LJZOhvsHhmez5mXz16IHAWFU2Wg2h
djFtK3gO5FcH8bCD6h8ECcB/MICb1SwjLgtw73fpBmA9X5m+Ck9KNDuuLjjTt3P52+icPZM+j8s5
xUJ/R/5iZ0lEo6/ayIOYHypjCsIE/51/9tTrPY6DwP3Wgzfl4t2KgtusEp3+FCiggfxy3th/zpz6
K0GczLmbaaBZUF8ikjPoJsk5WJz9qnUspEZR2579zQmZj0CSS+IEiGF60zBPss5+c1QTn3PrKB0X
G/sK3AcTzV/q4OkHGbfyJ9USmERHRsby1Y0zrjeVDdGykxELzo9UEN+jsqfbxHgbz4pRlaiMVnWB
fDdtTu23JoBgWRWWxOHMk0iJxHxk1v68kfrgchQ+V31idHRBooutGyE40e4oWfBAkJRKnAQ7ANf9
zP9Jjz8VhIGL88ZDp70rpkgpUKBUj9uJEDpjFtxJHNiVh0slHEm2faPBEL3tIotWSYI+xDRD4Zw5
CbTa+rYDxaQVaziaymrO6gEa3YD+v3gTojOcu/1bN3Gt9RCEvisF4SSzGDtmtyDXjw7g7T8ZVyEL
e7pj5YHWBwoDRLbVK0d4ZpxxEpQNIKmanKWJimxaCXP+/fYCe31YAVZCqGYIQrlYt0UoT4eDoYQe
I6Ecp6StNybyO74Dz7gJUICx9oAhdh9qwv3wbYxCkZjW5AwPk+oJjsleHBTy+gI9NTz5VSp64PTC
Q1mC4579aEkBSB5I+3GHhyEN5rXlBUoRbmcx8/meazjomMwKGgJL28W25IC9/gomXIscRpVHFJXE
a+eXiXTQWcBXDrl5TBWg/1DUYn6TBP6Ee8pErROCHvqmVz+xmqa1oS/32dAdtcK5ayfpB4De6LP0
74nLZgOs10UvU6nUT8jfYS7ZlBM7V2PzWdBS4Et5HEOIkV2b9PKT0PicLM80jm0cEvQtRRHhw59O
gv9tTphPK0CJkNkIedSwU8UoBrTHNfeVw/Um6dd/ZSpWy0XEKAMyFbhIxHcJPUYzdzxDck5iYTEK
HwMzvOAhuyIQSxsIKZT7JGGzceVATUnzJ+hbdY0YWPzARtkq6riZ1QaGzsIG9tvjxOWh4K1UV8Au
yLNeDlepEH+KoKma2PqyYVNanGDNSPeiqDjHoWqZe011zdjiT+3OKWKYDCKc1BftZww9PmunSs7/
pl9JreKQ0ScgUAH2mxjcTmo/Zsh2VX8icuHo47+3uRtckw2jzZeftwYpb+XB3/aKGenl8O0rNqLE
82j9Q9MuJGONN07dm3bL+HNZc1oDgQ4qpSU+OziWf4zXu8F+BUixkNt1y/nWCPV9tWl36riedcdv
MnAxc3Eiqqxuw8LXdIbO5WfBoSkdGsnLuwn1Gr1+U6+afAfaphgsmGKX37Zmjy7XSLvQkgYR4hoz
uRlg61ruK+u1kQWRcs0RrDxBvsC/zr8sAnPzcSpa4KKA0RFBj+1mKtvr8lrX1cQK94zRICE1DDmW
u7R14rSOPD9lnX76yJQOa57Aq5LGQQUtcoD09+iFe0TZ3SXxbWg7JGR1aOHS9jNG8tylSctrz9sv
HuWyA1dsx3FEGmBGWB0WVZS5yUN/2+3f2Il75pi2noXjvHYiMhS+wML5xJ1ghAK2I8fYZmqt6SHY
e7UoO8EK4UWMWdoF6kxDzyBXlJZ3qNxApMvHrc/KVhIsLZVv7P8XrIvU3UuIYnzliRzu0fuLvzg0
jSNdRxsx2hdaNnUrFyRwktkZpsJfxKL0SRn4EDJFtdZ6FWsB0RSEuX36GO3h0fQz2lDQ2839Fi8P
9qtPQK9EhQpt3LV2amRO9HfL0AFcr8fUe396StEmY64/P4AZJUKmKqHlFo+hTEuCLoHLtDI6sCpD
L3B9uJS5xRvFryEnT+sLfNb6wyqyeb/apHBMeB5hJDItT6eaLyrqgDZVhBFqCwhs+Q5+XJf99NHW
uR1uUYWgrA8Sd/T9lQMkAoi+5hRqSDF6hINLvU/wufU+EldxJ8BWp5NWyo4Az4s1h98R4qGhaK1+
9EVsK/zbVL+LAhfD+0RKUFkD+aBvVsvLq7f1NuvlgzPu0lqm3w4m6lJKGhkdYWa6ouJy/en/CzJF
RuEWDtPhgTEEAnnGYXp9IYcYDAWbZYyQZwOv1UYjOO1FdCpE8Yo3jw0l9gizSQ6CWpJEhqfjTQUg
ht/GuNO8664JNsvhmHTNgA5ijCqtziZEjwridMo9M0Vp9JfkOdwckE/31Ivlu3QxpDnR9VK4jsAy
lezm9n/zRjCeR4clQo5twfBC4sk/vUJS0YC5VHqY2nUMFUdW36T+0UG72Y6UMUO/g7z0D2nGf4Iq
jmdyp4VtXAXGmPMFkRbIzeMeA/M9aD2ryedH/PnFAITiSjYgyl9eYwNtPyumfoyNGGlpTZ2aCjGY
htGsuxrHkHZZQnzdNgvjNTciDftdLOK6H10JJL8pI62eZnZHRzv3mRNbntbSc7rvilFxefzoQlfx
QkaIw4fl3J6U/BeRxnQCFPCoMJcYgdMg+MXkhKl583yh/VL8k8rZnZcjsC7ZfXIoDO/Gy6Pmz+py
CEOtLHha/MPfAWSk7glZ9BWl+DDux0ZEKW8N/jzqomMPeJ5ln0f0b5sKdr3HFDZo74RNCGY1MCwI
ILHtqjlBs6J129Y3Vjj3gF/wzopDPDCSzbTx6mehxc5Lwccpp4QUAisdzk36lOoR5L/8tSN03eL+
DoV8AXMvlHjdVzhFUgbf8S2wwoeVoaJaAxff8+nFTPluzmFbTNdKofkCHZ8NioxSMTBSJKxHxn11
FpuK7w8G2XIF/Xunwck6+1Q/udkDYAVPTN6iRLsLNC/loEc6UY+tdYzKlzIaBKYS9t237ZU7ggDF
Qlxy/CWaA7RRw/qtTp4jj4mLoYLuyXTgys6DiH4X/8rrSv+IC843fsL+bz/mMjPXBewWVNckYayf
YTD6kVhyFPHwaA+/TLeKrydUi/O5sjgWnENc42Zuvy9fD+ImFnwi4dIQzfySiE4XYeA711ilbl/7
hgebu8ui5s26d0uJpuvwTeUl4BshKeGI/7SxqGeeXrxg9eSlWz00zpKqeJ0R/R9AogH8SvIuNgWv
JwQgWlJY+1Aez0p3yjb5cfWDftSVBIkOW9lDHuUcN2oS96EGLjt+ScvBWpQNSgN2+D6fjqK16Hjj
2vzktHWduqDDE3yqzLYhG+jGCVCeEAHkMKwS3BpZbirVLPseNF9SDuPgmdT5OV6xjeMzcjgsMUDn
GVYoz53O6xg0XDuKyK6BLKNESFn+CcmZiT0uwi1bZePMcUnWNEl6kzwAPqYcrM0hMHfhnqCxYUul
0ocODDpER1tDkV8kGIZtIz09BTNSO3Z3PRX3kFeeO8VndVMh6vhMKb6efFIi/9X29yY/2wWhr+nd
NbA8dAGOEN3CgUblIdUZPSothfAD0jQHviRN2L6y2OeMNNiAnQEquE/KbX0ClItKi/AxJ+Y98EyT
KkfE9HLMbNfK7ZMPu3Z4o/zz9ptpqtaNCS9thOz4dxMf8FkGGCMYBWQI+5+fyEhMpuQzcJLFEL8T
SARHTs4BKVVYf9+j61DYqCe8V56GpmGj/CKgQzKCSrjSpem3uEmtYPyQzZRmPlFkJcfC3pEr0D8p
iS3DUMtieFSt2PzwRWW0rlzNAOuithTzQ0s8JMmzKnrnlmVQMtpZLXJf2cH9X8o2uax/bJEfyIhm
6gnz2hvD/sBQmRHEEGcbjn9mwM26kZ8A3M/AetZa4zCyU8qiPJS1mlC44+f0l+lQvhZMBp/CzSSa
JQqQHHYxDTYEPxRxTH9xjIeLPC7cchR3CXU67FPTbG85q3bsTvSx7UPV+gOWdgvQr87RrFhXh2ny
M4Pc89bBJgL05V/rYHlvtFS7T77p6o4YFbKFwto3vUKETaWul5zPR1r6ACn0ppG91x6flq8HNVyY
SlFZkST4SUtl8Pf7fU1WPJs+K9ZI8KEioUZbXjurLCOyREZ9TjPd9O/OyxBAc0rNjeh6+JJOQW3i
Dnd01qekuKRqVj0EzGMub6f6yckeAzxmnbz9MNAuIlgKAaY1aIOwj2WIznjGNThkhrlV8wzkhRcq
X6CuepR216xfbrtTFkMDTo3HO2KG+zliMvK3nF/olC27d4cW+A7XKpTkissv+IeHF+VVLC1LAoAT
3YG/J3/U25NipMoqbyXe49M/yYfIlPkHfxJVIHJEIkd3eIb2TXAbh7CVdBPsfKbvECvSgogofjor
C7RsET9RErk5Of/HHTrqeqwABXXM09OLcRbvLLVq+p61fQybNNG6V8nZZ7gOIfXcMh/eYNxTU+UI
/fqOtb479/i1DFSW3lSlbN14JhR1F21zI35Dg0gi54FLJrLCzqMKahlzjUlh/PSVKdKdQekfVf6l
spd5aTftvu7P/WQ/59JlwB/4bqbHCxmWuH5kyEAlb3ubyDve4WDeJoDqYfcYSy2OJe4mhBp31ERV
D7MuXYB08BM3ON/ntyWsPUsLupMqPiflB76NPiKYaRx4vCyTFEUEKEQ6cQEfk80ajmSl2MBPmsro
YSsISrhbA4/kwkAS5A9IoI9qM9zB/bw5226zLnforBXV9aM/r9egCKrxDGqmsH2FPOCCA/l+BQWp
yrBDri1OxwMZxDD9PqwFMazjPtXzXyNVY/aEwYJevff5uZMzDzOO8ld5YpmgzjzkmVcCzCoUzZ8F
nGoFgQKPz645eVG/nsqHpXizoJcIju7kjDyBaJ2XibH/dfK76msJ0xy/ZrKKVUOO627oLcKsQuL9
FXkybYXn6EoPJLpLPHrrCZzMwVpOe6CDi9xoQCOtsc+hEWK1F/foo3SkbQH2Me5pMTuZJlIF0xXB
gFscphzZ4KecDCXSJZZl0KmI1J1xGOwoglTV8SOKvEs9N33Wbq0kyLPiKWscvOCoJRdBs0x38gzs
WGB+Vm4AqOSmNfu36aGLzBlmEJnw/wCD6HH/E1iACALLRPY8bpmJaHZ4gTtbsPqmt9UrVAw47RY5
XFQ2bx9RUeStytNhhwEsPTC7dnBYKvuclOSml8PapnVcugXz+sV/5Ty3xmTU9851x+VdAx/UwLlq
P7BMh7R3O51VH1PciCP+z8vPd8psV6N9C8FC6NcpGsbA5rFmEJk4pwUE0t6oojD7K4X9PTTjAaXO
0JodplwEplEsGQEtsdLnTXfN1wAKRRvZDOfCYTxWtU4gpYIL292/2qjQD0gyukjKlT5Nmz6UX2KZ
sWJkk+O/iApX9TJ0hU7S3C4hq7oVfrB8jGyBEy7JnYXtD0M4j/NyqREYETfOjgs3gfiIgM0KDVR+
xlbD9X07l4RD7oQq5f+Zas0KvAP/wIgdWXYkprtvz61mffARdvrpST2j+ngAMi3OPrnRYwhr09RG
rXH5pdJxHGoHWGbFsbC+bnknYDmYyrWe5MhONXtHfPX7HTPuwjZLoHB9JA9HClVNACc7cw9zLV4X
vs9AI94stEXPFkEZOQHg5j88c/D1507x7A0BCJEoHmZs0QiCIURAqIaAbUVFM8Rxhy4IayYe5MY9
ChqrCVlRmRqg9n4HHlGDnTLANkUEARVn0oNKM/iK2TvqXWz9yPbJ5AauyKhAq1I2M3OvxC2hbHcc
jR3FlbC09k5KFGyfATuBpki8QvNPmVwtw7e4kqRzgPYTGU40yL22MJ2GGM7KTn9e2uVHEWSiYWdu
2gUTU685u4supKQDpqVU+V3Wv5ezsF20jYZt8Q4vIiZ6+N8Q5GFvEPLOgB8UMeKUWWIqrc8pWmqM
ByyyGQ3MXXYTTjPzmo29W5wnJ25Ti3Kyr0hCbxoQWocdo5ry/ukidlRAo8QEKF0ipBasTloLz/1f
v+2hK2X+fyfJcfR8cQzFLf58Sp7TMno5Uvsx7q6ECeOFHhhCOTP7w828Y/0CkqgmGtBC9B86ghW0
Lk4ZHiXMep1OYvzwJOtOerX2+04teQUdnAkOT1m2/gSjEU2miOGky/8rpgvO6920GJmuIP6qk0sb
qB80zwNNWNxaWARhvLbyHWrAVJvT9Zrm77y+03l2rbBttJhM45Pz/nKwi3rRn67l9EaEzj1r423E
jlQ5or38UpQCBucEGjZlRL7IpNfHpeUaOb8rZESrYrWDSf+FvqMmYYniD7e50gJB3DADOQ4WWzd1
J3UxjHa6qPsnIn2K5A/e7ivUtXpnYMdCp7IpEdspA29k6UeOs83oykC3dCRSesDj10WtZ25zI9Hy
JY98UCQ4D9F80hoymOP0BZP1tHVQHDTDzvnFXW2KMOuIvcuJXcthi0FGHWRGYwEq3AfqT+MlVpxo
x95DAUGy2u9Sky3ikjfhlYq0NfP0e+jzk0H7ZcabmvaDR2pP82Bgfl13p4zJ54jhl8tIrk5AlHrn
IU891tmZn2qMusb/YUUEo9sd/K+j3AvjhGk8HU6DESKph5/O6lsDDTnfnDhwr0mO4ETFiI/533KN
B/CRgIXg+fyVgxeE+hJZCayQmW3Sn6GhaWfYLlFQYgDEu0OvBynhDMvZN3ulM1xR6yKcH3LBW+Mv
tlzz1nYyfX+l0uycuKEgaoQvbcyCso/K8YhIr2SQe2PLgR7pwRmaLxvF0zYvBNWAheYAAQaq2Ogm
nimJYvG0f7aWw0YdbiZ3GJMarv+w//2GV9PgbpeQbH7ZqkugKJ0dADV3U4RgPKpfhmExWeUQKaJF
/m9EMpl896PYj1TBZYL8rl5Al8pJqoaNTH+jYDdCidgsH9Sv1/82Yl1RIeDtzSSVzSUT8qzbWvrl
r+RRM2GZ1nB8HqQReDuWi2W8LoGwKGAJepOooRT6+J7vjx/e3vKbcfnkTbs/zhE1h4eR3rn9h1pG
XCZERgGjuJPexy55I4QW1OhjndFmMy+dbuMgk4/9pXjI35XN+rpqi17PDBXGC54q5gRjssashizL
z4SxVON+uyjCAkEGhMPaA8ZoLll4HwoQtILnFy2pmcL+O+3PH2KMXRCF9n2Zcyiznha9JhI5Eb9v
UgbGhpgLYHItOUnOH63f4DBzmAfIdlG9bO1wdQs+v5h5VZbTuQ5sd4IFwAe0V2jHi/UHzCKa2txF
LgM6toOGiu0jeWRX+gDhMgAx6Bw0vibQMlElEF/k9K93fah6tqxnP/aHHMODFjTt8VdwmUlDBuB7
jZGjOBkJ74Nszvo0+8elziZ12ib+Pwh+AjBtk0pllL+bjw/rKfBDnUR8znfoTy+d2UTRPfgJsutS
M6rVMTnKJXaaaSU/NYA6YWDz0XtB8XL13aWzaOiUEn93LWZXFuDglo4F8TkH4+12y0A5ZwTpn9yG
Lcl9nugRTmekJXQxC1CFhhV9Xkd0OROyFxe5Da7/eM1zdGrtlBzu+pefhD17dej8ZCiz+c4o2SVK
a8BH/2ulfDebp5QnmcPYGzJ+k/MtcKBZzCac8cl7YKDm/En5DkNrVPtzgP1+rbfNDPEVag4G920x
78eGD1om6dYiLr2OyA1qPEggQtDTN12LLjpuPtFHnN6N/o3m4SOiI91fsdxQf2cudMHS5TdmG2uN
qoYlNgE5PnqTNhIQ8+EUWQJWYxpxSJvlTjgWWVHr5EC7mvis9NNVsTZGC4EojBe/hgqAXSHEBCPU
2kJtl+7eI3mngfSYULwDwQZ5uEFh21LoMwTrX0M6FBWgqO9JOlQlkWBvoxHG3PzkEJmzSX/2CR9A
GsZvl2KQxy9FVyUHQ77xWx0eKZzIqKfP9QIeA2yDTN90AtsuWMsUIfwY815UrvEwizwHtlEcyBDb
m6mY7wdkeOgsGJ+Kc7NbSGmqir0BWauYpotgsCMo3XnIHO/pV+8i3p3Z6qfBv7SKmiH8ssdQ9XcR
gh3KVsiaucVn3Og22ovGTIHH9dT50VVDxEtFUbgxgC8ak5Ms/7rsd0aid2aYS9zvadBTAzihh1MQ
tS358w5+A1fVPE0N4tzK7P80rvXdDrHpgcyQ9ukCmLLAK4MRJRsVcQN8CpKIS7lRsulwnPmhhsIQ
CimA800T3yJfCofje6wOtFYmuXZpgYgf0b2jBynG5GCmz/RRp56WF287Yot34jYGwJeKNU+4sYzl
bltYYEpAgGyQckebLo1LcSIap4a1dOzPaC+yktYgFRlIPOR3xQm8dHdTrNL5kXDQU09gBG2n74d8
0EMgZgl2sbocnsuTFwhVP7mO5OhmKPlQP3TdDVRM+1NyRaeMHDQWJqsrkfws90a54L2Ks20rUVw+
xYXJofhKuI5jPc8HBINTAXs3aJmJf/3vyJ2ciUhrkFJTDQM/0dnQcRgPYzDhtpzeFYeUt6Ipblvj
h+ZllWzvO1XI1VVlSkAQ8ifhACSBwSjY9spS0fJE3QZ6oYkJaNKMpS5RLO+TDtq2m30pOL9E3YFp
ZLFE3PWTA12uhEwUDKglZ66Bs2Lkl0/Sn0cJOc9vJQ4bqfyXO/alfnuHIOqi0PBpHXBn7Gmb/mtv
U04BuWFgfIa1hZpi3YO/iDAqi1nlYu5EKSEa4y0+dhw3/miuFne9oZoOulewjpCUOavNOH6luvo8
QBUVdhSiyCk5KPAY8+bToqnGFiOjiCS+qRO8LafnTFxeMwp97oeTKsYURh0Z1EY+dWmNLUM/Gv+o
6IO6F8qgsf8XNFbgKsM0xuQyMLeNtSTlNsbx5dP5DXFOGg/tUMini8ihD0exZLSuPXXpRFR8yS/y
vD/7JmzNv1IPoaQia94gpkXLzak5Ww9KW+5CqPXqO+J9fgnc8H5YXv3tHSyBiKtidIIDTHF8VMH2
cPvMrv7ciRs+kMKnQDMxJ/raWW86ykhZ65KdoiD6FvSd38AOcodv5C7UmS//86DCxgQvHnr6nSt9
vwt7DlU3DWjQKHyk/VPkQz/hZZ54/O4fDUoxHTzbOfU6Qx2VxGZp8XCn5o1X6Et5eK4SfJioAlAv
raWOIQIxYUXEr6UDmfsBNXPIPRE4DRvb/DjnEHxPprw/LafOvKzEKxVicCXLnoC0LT00GlhhGzuA
Ktu4HaZvLY6dtcHSrLkVfZ+Kl/jCephHZkELgjFQcnFpm3TA0V5RFvNpCoxl6vdNtC1iKcKEkWXZ
wb+SGlypoMY72olmdngTOxjJqoQBqo6x5Em6aQUjBsOnuN18QPVhbqGaXpEj5+cXao3hGiSGBSKu
Ai1/VH6FDdqo+WvxiCJJopg0W2e+sgidswIY3+l6w1Ftqs7tmdbLW7HmX+9MLc5zDH9MEy/Axvtv
/wEUnFookKJ9MhFw1f1q9/q21L3hKewEPHd/v2L22S9uSND6Qq4slGJwaJGd9ZiNdeeo1B1C2LQc
Os0/GjDV6ehR32KHywtsdvHkMDi26bxowvhuwJ+i4w2jAA0hGsvMsjMMkrA/T7pL8uAs3UTOJop2
ibQImXmofvx1ezO7GnxP4M1hLdnu5YEO70CkjEBQITrVrePxuTuEPAwlZ66oclmss3oUObbGqyJg
ktDOn+cZt+1kjfKWs7PAKzzCONUvF36I2LZBqlIMHq4mCVpuq9agk/FNuDsHWCZ7pF2U9btqaFQ2
YgjqGnPeQhS8MROxwUtkjYVpokebqmqsmVL3Jdy4ubuEaXRyfr2RIcN32fxBhm3KDWoOKnujOAEe
Nj/ie9X+lo/8ofRuBbAgBhgFKMSYJAmBZCvAYPDw6U/RheNqcPEaOQNGwxmPnp5xwhiPDo6ZZRlJ
KiOBQqIJ+ab9+BWK/HBJDVjopc6yneLQmLmzmGopvyIrPOlQuDWg+zLi7IqpEH537BvS0LPLEdbm
TJ35wcNNwlrRq7Eyza4sjAyP10ieVBzxAzcHuoVTsXxMo79q4JL+AvwS0hqoVJXgULAqHKGfrSDk
Lqd0dUkPPoz9TFzwm/OIfHoutnqVPSRb87Q4E4oIT1ApAQ2n6MqA1hMEjbqPjlsTmhn8BPGIgMx/
S0W5Y+QKSKdQwd/kNYznAIooeHe9IE6tbh9sT50ZRooupo5gm1VCD1Vhvh/gJ+VTF9NUi22vL6O5
y+++aQxlSGi7E34VkZCPBcjJB/jqMkiL37Ul5HMMZuRIaKmtijsb2p6Pg0arCxhAdI2qXruchq+T
PW766D5g8Z2g3WR60Q3q0F3AgICfJ6/U3q46pOS9ykZGXc77E4WlFMdrj31QsPDkhNtn4J4p6iMQ
QVtKyj75Ds0A4XpkjX8a2hV1SQ2axLwoL4rhOZVnVXyvgqcOEoHSFfkig+qAhL7tB5nCRj7nWcB9
5t1yopi3HJVIoFP/qHufz72mpXZ/2O+wzA5qQJb5tZjNoh8U1qOzGLEdBYmAAQY+0wf0JoQEIIGS
At5SrwqiymH+SD+AHKzoZs6YbWQSaJTw6P8VCaM9qghvmQwtDi/wUmevyxc/qxXLTX1hf4DcJeYh
MG9/CWf+1CdI1YBIEYrtnO63k8ukanEJ/BHDh5W6Ry/8geGG1252XQbuRFrg9mgkNduiATTSSQhL
naDG5yFza36B388+pLjLTWVWMDemmmSvEXP1crVDrxjUK8u/hOpypX6U/zbTZzf2tvjEjcB4DjoO
SBGCv3tSLQrK0+761PAzJgeHzNXMWFLzKOI/MnxWaB85LCMq+XlZ7j+A8Vmm7G0G/xCo6t8FUjQj
4Pc/+ygg5NW+f6s21VdtBLPSD4qu27OmYQeuc0tWUD/Hv64wGvtC2hmR7gTGTnBM8Z1uRwTsdC6O
XasnHpFGf5Nn3mghqoavfUch78b3Y2YpNZSEouYjsQS4DJSLXIZYIqXQAW/4Z9SUXrZ88Tr5aIM8
7QDIXsQsLMPAFM6hABnflHC3dPHKNxOREHEINfQjoGv7xt8ELZjygCkuowrGLFW0+JLsOTJYsqnT
iMPSa/y6NTvr5T2z0MqXW9YkyMcGYwlOGwxyu9yX06uJsX2LCohpJZ5uEBy/vgBgiarFrPLva/19
9iDds0H+fSDPGONfWEzh8Hz9ntA0fRiOgDmd9rhFjEZHZJHMNI1ILeTV08rhe3jZwdYGbnjYnpHH
affLtmkuONryFNvHKa9WD23jIZ3BbMnLViNw6/UmGXQfD8NqSfjMb0z4lbKtYCLaJyNr0MBhmYB3
MqpJfQmwkDL7iGuJUAD6SMkT44/4b+/SvKhOxOcYC8AFBExVKRfagNMeOgdkEHdww27O1gjmyAXU
trW9LjvRPxl3mqjE10QyDeQsqvz6domNhQoN6klkXzNYS8zvloNmmzjclpLX13ZSCB/V7KSxTn+E
KWUIoBxU5kTP7+ww71FXI06JjVmsydLYfwfenvVF0k7phlBLgdbb/XklIv09xFKERcHIQ4WFuxH2
VvDxyAqIvW+qHU8wxAMA2vqiBQcJ6oIEP4BJUWObCTa4Yl2qnQKMSiuG3TH0+mdkk+HfOuyUhqAz
D8+OTkEczx3kdryvpWCr9lb0Ql0b4kaT4LRWnv5bvr4UhCxBhbzds0e93pubCYVSnO3zwshKxRVf
5EEmu0V5zENKMXfB9VbyjF/QBkxpcr8bcOkhlqrxYPe2YzgaWumDtmjGOWiX/T1Xf3DjCusY4Ydo
oq/Fbx1jvcx2cB4GFzYOHeDGqiwbBoRlbH1YoCi0wg5rkvFQqsRKD6xXDPLzjB4eKS/KQUqee1+T
fppHswOv012GhZWDfpycKSZ/jUP1AUVvlFB+SOBrsH0XektvjTfNCZ1QwMqumHQ5w2CwbCC6yaUZ
poIxXRD2I+IcxryuWfDhQCs2k5xyXcFw37ocIu0UwDs+N0jKylqlXsv1ULwT5oiZCCMI0lQwuDOx
jLX2L+9zjFAQZ4nPdGeD7BgbvtVc1wHZPQZxSNr96BqXDCNA89cpS61vl+qIEbXV6etEMmVgVwLX
Gu2cYt2ZnVzNGB8tc47bAfwVZshVZERLI1aVDCg9p1IAdGb2VzIZjMYRKDOjXJeVvwxXAydRbjZh
HEf30J9OQLPF75gO0qE0ur72G8TBswmAkbPf8yMEg5fD/l+VkO8N5wrvEPQUxtaPZWzi/ToxZ+EO
cbSeaPcwjGwXzQGAiDxT88sj1WXgKaiuqbwENlyDjB6/2l4mDEqvTXn4VQa4nu7mSQ62xmyS9/DC
UAroi8u0Mjpu7ibNL1MBE+upjPdljsRNPNq27EEQ/C07pviSpNM9VdqHQjhAN4K+oBj5MPS/veuc
19y60Aw6t+EJ8nmvdmZAt3ddCDjlI3+FyQ4T9WDd/V6oRagc5Z8VSUebeZIBA/7rZScL2ZsI1vnM
i7Pyrfoob+hkm0XugXBE+Rwo6OMxjketNi1mFvZWK8YlhjxtdPzElNVB6f3DG8G+ujbk1PQtGNxo
Rj8WRhiCjuKtS2Z3mLJmnDMWbxYmqjgZNB8iXMRggbDSre1ckKsDB8X2WcYi0cREU1t4EjYbyRKe
g2rVMN9CD/vgw++QajpePXnkMVDpHt1E0a1BV2JqSF1a+JmksvqMzxiOlk/sMOLdlSJg6VIxiINF
HSvdc5hyJc4H77vkqHMsCREM8TQhXqM4Qk0BCMPf1FCvKlhoz7lCwztjaaXjMWxa54JkAlrVcYat
9tYuhA7dZZ7GlPXm5x9I+mrZsXeWHQZxOuytJoORnT5InStFRZDqNeZdXbHjT4DbYWfl9PkDSDbx
Ke5Y2IGJM+iGrjgpSGkBeZHvgHdaQuPLvOpnpexrO1z5EP+4PD0BEnYiifijTpVWIkE8AjlZau1O
RVqorweEQlzGJDDm9jff/za3H1ERNtrUannYxI4olQfUe/j4160o4UVWs6jhFER8uyZ9iWLBS/Ji
h2Cp8Bu9bZWjZaiW3TeUXar/o3j5gvobJ28v9lRClnsIkcPkjDse/ikDN7wTpJwq5mzAXwbMW8EM
SNMAFcoeRfYBTmZx7zwQY4voRyA2UEJUnMhy6ZHhTLlFFhdM+8k78hgdXYsMkRZf/8cXPMwCyk7M
a6tYuoj1shFphnvyCU/nYy3xRzhl7TxsI5HJAQg6HK7eJNxEmw2pdlKkz6LsPKGSuqy3Ku4Ovpaw
j5TfpSDBpXhObhvfxwfKBO2EHqJKg/6l3WUvSHGhOvwD4FSRUZweb0fWYNO4ZdExmoWXUFGpHS+9
5sbtXTzsFE5w1j21/8HG0ayB579OK8GsWlQfYrdftOJ86XEvo8EJCdNYGJmDdlX8JLucDjYTuF0I
A5NPwO4ocYhKaCwyi0fBinA90HtqXmMbhEhMjn9Z52nbWXNUZ0oRP0OMmyK+3byI2Wa4ZkqLG6rh
oBNFFbbaBSimf7BT+NzqU3n8cSDzHWXfRpTZBwtYcbC+gBwyggR9FXI4YSEK8mCrsBqbMsqgLKJn
PngQahHw4VeinZb77GhfPUoMWXyZ5LH8eOw7QYLiITJUORGWR3bEAcVLKKQuwP2+PnIT6FJFGSTt
8O8FIlpflkYnK1s052Ivj1BYaXAotdSW7EgtEDvl9OzX4uGyklZy4zfEmB4mi8wC2lwToJdWNdUi
aiKckOB1uYkohdDttvCE2u5oCz/Dza5hiwH8FkfxArSuBPB3n3NSgPJhMdQOVBKZOEThX2cSEATe
nSY31PktqO29JbeYQ7TXfUTSFpfwJfwjjOqXG+NXs//BeMlXBW5GDNVPoX/MfprwB+7FjyHwT++E
HCNJseMShHB0D2YKU7ztuZ3WKcE+xGGZpFoq7ANPfswbb4VmUiDxZAZggE+NE8r/CdsU1eQfON1d
4pwUBZNoWI47RYsnMexcLaEB/jE1nmaOFbf/rCjxgGtAKXztPtYaBqSHbAcYg2oCYOdQ3fsQmLF2
UrLKQBW4TN321KgxDnPOxBYMqzkvXBdVPMHjn8s62T0mnFuT1EaoTrQ55HZCLD/aONJp+taY6/8U
HbcERlzcjWB7hDiKCtZvPLTHMMs8JfBx1oIZGiP4H7tRFuHQWZLWE/LRqN/fTW4g0GMtUPsO2FRV
wPpP5iqokRXkZFAfiVo8RJe7oDdK+2mUrBOBiykYiB8VD1Bqmk4k+DRnMDYNdIZy9VpMJPnr00Vj
nGLknVWOwRjknBeY3u6al8adXztLtJa3s++Q5SsoXX91BDe5PrrD7qAE9Kdl8zlaJWfzKFNKdm50
jln0Yn65l4Hy1//S5wpoERXrIvByKSBlPd0ZyWNqiQGtGMhwJVydlnC0TY7pc3q0YhZWmJDgZHHk
pdmunw6fTQ2Gx7l2H4K/oTx0e6OaUO/PvEbM8SIawXLYyfyu5pD9nsD0EV1ptOcFQ4narUf6PYUT
t5WToK2QRU4nrbPCwdL3yDPu1KC5w4EPp/MbeKMdIq2t8/Es0IEv8kB6gxqXd0vpxif7VUsYWQh9
nexF32Dicj5sb/H65HG3dG3JdNB9hDatO5AMFl3e1z3imb7H5gvkdUYHJzQHW/AtAaBGtFQZelhy
TmAXrodviWhfZ9PbA/UEzr1L8FIRi0L5ntJS6p5tIUEEdiwppsqrDVRJPUk8Pg7n09YhOQFyIy2b
3qi5Qs3LKehgElvjl3uUIXdLNnhOOI4S27nfEJveaNHnBtyQ6XIkcJIdVgGzkvp0LUPNSxYJfwZd
tiZg93bi2sqeVrDFZ6aVY8tCJc3BmGMEUQ7TvvqRlUHIj+rrBxPJf8qrvyrqOKTbsOVuELbvY46D
q3na5Bcs9iIvXhngt48AmXUGDRjdFV7fu0HUFfDJMrugETnL7gV0D2+uvGyLgAc0MYjXVXRSp8u1
2VAlZ8Co5N7ExAlcxACNktEcJ8rj8WIeXxBLiJcj7oRlYoKdFf2O707vEbFBeGIGFcJ3VJ0m/NLw
oOF0ZQ/zKqQviA0iroe4r7YJwgaqqhEVsPDeRJedIbHr7lyHwxC+dBLwkwqOaT1HVafKoDpSJL/D
cbfMWWfA/c+8OA9gluB9qVf1YWqSHfkNAiZdeO2BiKOBUts6ZFj2RkmCkJwZiIyGinPSLWxe0lme
p4llOejCtt0alwxdMOL02oMifibMLiMOTt/vePngAAigT0fakX7EJHd880teTbAlyg/pqLaU2Md7
/MrvY5UpZT5ydVXX1UwNyo/hRW7D2teSG4FdFinjIY050+aim9jDomHoOV3uwClymz5liGMhAYho
3KJi1WOm4mT7JWy1nHTNoHC6T291oZ/cgSZqpS685NsEvXuoVFwPkFVLrTR/ESc8XXeGR5BWNZWl
OuvKe7KAGw2OMiyBGdNA7aEtSEnQkQK+iSpYTtLygIEc9C1/WRHtKXHPOH9hFcfsodfHxPZyBjdx
/jzBjKOaseZfohpZIbcx5FGrlGjFMxtWh7dtXIsuxpA61ZCNtyB7bNjptdHXmA451xULyh5RWSt5
LSINbZ/Has9p/I2ZDHgqgZpUAufn8d0TeaGXFqX7v9RuFHkdMu+/XnvR9bSAe/My3WpkxkJQLMb9
lE1oOi2n8Ac1B9FRgunznWgRX/DwFF7r8ouKfvjFB38pukkR76+7p9M8kX/pKy9cKA03zWlyPMXA
Q0a8RS8iHLcHJz8gtcUrWWswQnHoBftWZhBJt5ha/spwWLbj155SyhYWQraWuF9OFqoCxM7I3AGB
hpauCrfhhKZCOnJ4xJaUmI/LendzJZXOCOBXdlAyu7RMhH/jDZvs/oDdcMozhI9VGFmytU0Xzn9/
3BxkERw8dCgEJOcdYKBx52Sqp/1ma+MQggNg8fmDHBVMmb5ZY8b44wBpHVoQwaa+kc1EMQOg6wAB
DIEpmUgC/hDXnXsEg/uQGouh21Pcw9z7a82H1JlK91hECEIO+AWVtgBOa+n4TWhw0AKg6WCtftSC
7s+McVTU8lk9pHR28NtJyK+BH8WbuuIP8/hFHc7JajJ4On9G4JikwxlC7j/6+4xe7YeVGQu74UGn
6QXx31oz7npnciux8P0d6xUmGHBjbMzmAhIKmiS/fSGaRO5pQnm6S3nA4j31qu62Qso5puqP1rpo
E7ZAZCH5i3LpyZcjLdrBCfMVH2S3Q5ECrnAd/MGXBLcDASWLAQxeEfr6Pnk+MJqVur/0P1y2GE0c
5Q+kq5Cwqg+fIe8jpHkp1fThyKsvcfLg1TEtzLR+QRFERtqhnl1oJB8wM5KTSmCNd+Xlo16GFrM6
zWXb0G4ZnuC+NRUcxhAaB6eB+oRpAhUYN4iUD+3WjBIRLlw/O2qTwJwlcbtVTXSyQttreXYFh1ia
A3W0Hn/R93lmsSsMoiyP/HrUvJKYFQfJVrQd3T/hvKNhCeFm9bSXGkwN5dUdPF/6R17tv0kBy/Li
5Iq36c2/pXY6j4XYftN6j37YVT6z3DMkWX9Hb+bMdioufIrPR8n8d+yjMJIAnSn/jE4JeBIVTEfy
kiEFZs9zpg2MZcgrUjSKYy25s904gk56VWTXve+cAJDMXcb042Z8f/RxDMn5j0SNGQbaolcXHFBd
a+VHNeet35lA3N+bIEOpZ306gW0CoZu+72GOt28ilI3liZ6vAyqPvDLQeO4i5aX0nM0mF/3rdwQU
XY1p6L3b7oA/JySr6JddifXi0kHPvp61WbeGaD8mIIGGPoSp36oI4PlZLOrUq+r7I8OcnDVxt0LX
bXTCFGzhjy8LYDIfcE1/RPiwEkW3zYi/NYoYCytKjb6mgLJ9MUgS/hhSXZrcFO2DY3prs8sTpFDN
E9SXRQAXt833sKSBG2rBswVPGLnWX/igXTh6P45D+ZBjr58aZncgtWa9Wb3QesTAICfnBVO4yzpF
3iHQgoa2chy6CClbZI+a2/jsucikHFBqSX6py6/73m0v1fBLXO/ul3bbpfNOys4cN1L3y5/x9jaZ
eevR1u7TRgfy7nTzE6oW2YW4pIt2BXsBhOJN/MluE6+7bTDLpeOfKb3QnPlBn08JoGffNwbEMx38
cHWOWwUTBl7LyTUzSjkjtGmbBzprrsvP/QqKNinucsapOzf97Rb6D7jjzIQOKbdG61eNamL5DFia
h5Lvg6y5dTL0Y+SqjKqFmb6Xjubh8ZBOoFF0Jmnv0/dqUJDHR/P0OhnR65BvKT/b9NzaPCZH/F4I
SefwJCuSI1xnY0WPNIBrRsjuiXEdoMjUthHb/nHn0Wt++rLbtZmRpeB9aIq1/zbWvO3NhNectmuo
pBtI3+Ruc0axLqVI8KLYecu8dyQtOoglpNMyCJuwOREUfH9Aw4YJdPqsfHnCzwB5MCIpbkErncbD
Xv0NyVr7+oA7xjedNyRkOFRA5Kf2eb2SFE42nA2zIdX0gZGt2LqjOJ9Ovpsk0vY/9hr9zM7iJQ0Q
Kv4FEYZFc9Z2gzU2tjxSAqouZu2bJ1m0mxinsdQNMu8fDGSlZ/MoY0HFt779knM/6HZsot+Qh80n
GlArfYtlnfbXlCIzsxb5537FIuJrS/gGm4fFcmElmePVFCIu8gg853a6duI7RihIjfAujB7SNfDD
FQwCmglH20e1E2YAS0OsxhvFQciFW7zELT6Y0fexeLTBOQ16Ibr9P1JekgLd8zXoh7ECNhJmbRgH
pOFyNzHxXAIxK+OmeY/tfMMuKjOiziLF53B6wuaFLxPHecYEjysCciWgbqLTB6xAL77AIGaoK9xt
3QudWLDoK17WhyxrHp4pX/oQTW5C4bectGRERUQmLlLWuuyNPjqq3zatQaOE5b59fKo6BkQn1A8t
R041Ski4ZBqdPreFwChsl+jqPddkNW4cm0q/usvVtm4Q3l2biEgROLrWD6Yi/YH9Gngt6OvbutN9
FHCPrjxVml7olQKyOtAfTBJAUmItICmHQrd4GTY4Yy6WfPEI4pcG9hZsCeuOILZ2qQGxpY2UoKOZ
/lhvHQXXlrPNtxcQ/EWTOvYKBa9JmSjcIewGbm2dwoxo7v1emLNuVzO9Hd7dnWVdHjdN8KcGV04O
JAMs1QmGCSI3SG+P0Ot6XLqyqdHjFYCplQ0uTZTuQR3iRXZD/aIvC5MZ6wlbJ4N5pZL17DDYTqp6
QXc6xHFw0bpE0idL2poR1VxC+MTStBG4tEicxSOj5QJwe0TAowJKf7qVYs/eMG/6WQDyeLos/z2v
Jyr2kEtnkG+QPMkDaCHa7y6ygRgutzxFoFxa9UaLAaCjFYIblFckSdxf4tjLSdmsNFpo3PZjgh3X
rVyCIg11Il6fA/fMppjjvO5+Dy3I11AFVuJw2IyX1VcuwoSqE1CE9x/i2Cu60jOO/dBHJUBD37rT
hQIi9oSWAyPvBXFDh/EN5g/fP507PFUVAq63V+PkBBp8QDk6hh8R6oHHs33lzuDWmytsHxaYF9wa
+I62gcAuQlDptxChpj87YXoCciWti65kC9SfqynWxgAqLhUS7qwb6avv1diIrfOsyaQTunCu/WlU
kDWMAe7zUTSO/SonHNCkTjKPOTcePDXc0oHXYWmGp2e6mmndvuHon8MdqCLvaHTxGxssi29Y7UFB
hAA1zygH6pYDwMRmj5bju4S3arDZUGBXiGSbsLnvjPd/bLDB6J8irytzpbALQYEvwGoNtcHWaUeR
qvTBeJvM08S992nU6q/02AqEH73IX0UQCw6NhuGKOajDQG5YjDTwyFsYdOdEXPOJEORQ2TAK9ie0
zbj7QEslIrnngLtlpVxk1UvPr9RF8miL0tg2e3rHVlzc0mr3QlK7U3L54UX9OBh6/KjhZf2xIMgk
Fn1jUMKUqf/1pneWuvUbTBCMzbrrIgopuSs86oq+9eoesbcOLagarcOQS74IoAu0R4uSCQax6l+q
5KVvIArp8IKEsYneVhPCNCc8go2Md7D9CKk/XCtNrvAWkaD5KYVkqC+5EFbM7etp74Rk5U+R/7TP
V+sgMbz2xNYsQA6kG4xef66cJgonKm6A3xJPVUk0mKYExfpowaYjudqAOWkF5tdX3gPqhEJHhAKZ
pKmhPAlKhgwt4RBcTDBLn3UIQZkZvy23cLJm95cOpJXppiOvwISkw/zyh8xtRP6fceJnX6Zac7es
TrPCkYcPvGTA6lYRkKO+0LA+D5cxY71DW/Efz3fGB8kr7t+rN/5NKOLWGzRyWYiPCURJjyImioMn
e+2EsVljXO+UN4cImIUFDBkef0IXPQ61j4wxcaYfHlZjRGZrk9IcoTjM5qmfuN8tpnEptbmijTwp
lXtNEPZRsYoWtuhqrJqM5nl4UkApPqn8Ru9vP2M+lL5tm+cNDzqKNd/L3X80y/7osKz0R3awYYRI
ydAkWz3+ecSOejMPSZTMreZarlY106DgS7/YmHJSImXhvxFl2CcReynxeqlJ/8LQxyuokqvBQB9X
vT0Q7hpibze3Kn9wz26azpXhEWcqcVoVSjjcH/BfeAKGW39k2ZB51k+q4hnJpW8blmUlb2eRosHk
m0HKf63oXPr52fO1DfJUZqlkdbHKAEBijzTYO1mBRtNZ0iLPBgrJ7wfhLEkwn31zKqhHRqGm9xjN
ferHVmHWkvm650sn9sWVtiDZ1G4O0PNz3fzlj4IKPb5nFpewoz54x18NQR/lOqTyvhBOHcvEtcgI
50atNMGyoy9HQdMFiiwvCeOtyS8btLUwpwtSqrZYRIOnhSiEro9NnIIOnexNR6s7hR+fv1cld4X2
+Krygsm/s7cJr5uuaCvyAmiz1lJnZmfwd7aWMuxS1frGrF6To1sXhZ1sp9oKJZS9uliFJK4CHyP6
v6jBMl3STTsrhww96ZTsEROXawmfGkMaHZVZRrn7A5s/gwpAtAFNifOCjvFStQfhUuvt00n3mDfM
TyhtS9zbzimV8fS+umfsgjmvkEBIG0c60psBnvGqFOuIPHC8w/XcKRO2Okv2tcTGu3tWAMqeRCtT
IgULR34C7eNLjNFLTOQ65CBN8Ie1MJkph38qBloZx/DiW/r48DDgegRllKbrKIbiY+jwtCOubRNI
FR9WMm98+rvWcHIatubMrDTRgqi/cMkyZve3Xd3Xdh+rhzjP1oc2O0W+kJHizVUxeLPVgTJNI3w0
i2G9dp5OnFuFGlGDWQbWxMHCTxuWko0eMXeDrzUcMy8dXpQmopvv9GtnxnA3wAO4nWe8LEsUlwyL
irqdcpd2BKgniJzrK91k36zBUcNIKBlY7/0jMVmgrYC3Q3k61NjUxozTVhgx+HxkoF4S+ZXhkwoV
rostqWusauT8mPLTih6d/gLTbmCmexJlOnnJhH1oaoykiWg4JX8poKbfq768f7vXw6ZT+VEVnCLW
y1kMzZc05cZFKA44FS1rnQPWYE6HN60PzGnQHKJu67trjALOIZbjfFYF1LseQlTx5i9+TLdlBADZ
MUBmYU3S14JG9DNlAyGr2fq5eGoXYYiPovaHLGQwCZ6/ZFrqX4bgSjcFgfoIycPokWEzZTsSBegS
Xa0c470povEWXBiW0TY9AjBdmb3FlrxRdKZyesoPdgy3ab3hc/P0cpDKt/LGi9UBFD52Pr9lLa1G
hwfJvfCUphIrMhQj+53uTVbpIB9k1UObEheqi/9rpapuIfxJvWTjq1k+51HH1N7OUx3FIZ+38lON
BiUbYLNCdr3tz06Qp404xa4ezkrkApzWLOaVyTwb9XixUanpUZcgNqCOO+jDUk86LWHirtGId1Mu
GFH+l3xT38BFQxBHWFTfux2kvDwc3z2pKE3BKzEmMAj7BlWrwTGZIozorK9FyjvZKjEQKTC51T2l
7Q1pttNyEyKlztMChS6pTS3dXIOVlKZtIQlvs9pf+G8BDqGTM4uS6jnhZop7rTXalJOnaNSIXgMf
cZ34ksMPJDDe/c6G2gWVCSuj6JeNMsJBKRrtm1jq3WtybIhffQVknzZ13DarLSmhVW3nIzk0Z3GA
9vdAuy2E8EM32aenOdKT+JJse7s9RY+JLXtzJZZ4w6pS6dADOOTmURvNsEbN3D1ubj60iEXUWY7z
ht1JoGp51wVmhnSSL9crj7aW3YuAYozDQOrsTakSA3XQdDpRvc5cb2n1sPmJXN3uV0eInesn2bxr
lgWupFC1kLVyGtf3FRDNpztK+Ap/EPPfTCQ7PY+FypGZLhhQ9L78LY9ot1aeSCynutzO0rKT6OXR
7SRGo7XwU8WY+oGGCOQnbKho8YKiOvfM2tdAqTJNEG4hCA+eKOXVF4mhncVIdT9LTcONe28+WSRD
jC3SHirHH/VxXX28+McwRbFFULAAFptWeqRf1OVqUEMFw5q1xDhuykmgL5PKkrMSDf6vfSr7OLuJ
wtdQHlbW+4Y3yElvm0SNZ/EFkGqHf4oo7ShmfX9HSvmF/M11POms9DLu818ZhGToZrY4p9DY3+g7
R7jwk6f6/4Eq8AvoAKgx2ZA9Ret9aS0K/mKXPDYir7YxzOhk3PPv2hAynv764F0+7Ulnywyv/jn0
xFmTHSCB+r1+oGkqYr83D6T8EKw7y7EueXY1bePq+vguOSlBlGUaQxKBLae0Tm8R9VXD1wGsvv2S
0d88mHwNSZtt4m7ahV4GsXysoe+q5y5x5BQGFHLW3TNbTfyMJphimi7aR2nYD7udhlH7evu9CR7+
DESqT4SRiRRl0ZZ5fTxxzwbBhAqjbQVSt7OhXiwrPAt8YDtf7ONCWRQTGTCUKYpYfSt8BYCXIr73
NF1Aui2Z+5dyo316znWBAG8fI+QYYW/bgo1sBU6L4rWAoRPn8fGrOwnG5zTRHlYfASOyf3I3ay49
IrWlDr+9ChsfIqVt4PM8IWTv9X7LEiUatoSiIgruPiqaK+Ik987CkgqRdTwky+NL+slMNidk97p/
vp9gUH55toq4/FZRCoiRslaA1IYIuqGKMKdhMJlO9KlJrtLdZHGwG9HYm8q7ytifSWpJUzQClsdM
B/co/RDRfeehzEIHsiEggVgA/t3abYrukB5XPaZKTODY9Ffh0xLh3wtZw64/959M3x/sGVpZGtRu
Co2u2L0ICY3Eg28Dl8Hpwe+vjO7FEuSIwo6X5geFAnGAl20JOqHASEpQGNhvAnPrymqPVs4z/g1Q
GnKb6LzED280UVR2vTvqu45JnOY7tTxAcGbo3g1zzaeQa1hibp4AGuZUWWiGFTimdhSMs4t2wGR1
4krqFhbpTiFKgxxw8IlLXBQ2iR9DFWTJ777w6YeGeEEmwdAVLcC7k2lKJaxg9VztncI4JGbUzjE3
pQpiyYM//55LDRl7dawqvpVFVfbTjgHOJ/fOJkOLDQMA/a2BiaC20249WQgOa4tXub0okv9ZsloT
UGG6InHzY5BsTc5Cp+vU7ellDVah11bvoVdlcMTFCWsFrs2hXF9Mu5cKL93lk5a7C9oIqFtUp8Xs
kMg4fCBYTe3QIz+lXFizw0/z7vgVFK6Le42xXeBf9hHn49MfImIT4JCnX3S8Y/Z5Xg5bMWHw24KA
QkpIK5n8ygp22K6Lg/fdCFhujTpQRPNEhKTXrDvmp5+kvQM+zdOS8fg6gP9vLan2egbcAk5CoblH
jBpfHD9v0AE0yBvqVhy24EDuawwVKCmOdIvAKrKijRQMrH/LpYbH2L3Nd2RC/JfYC2oqyfJ+ToBU
+ryzpLoLf38J9MOkt5ds8Q/Mnxp5t4XOGsX+cniYPslVkTOK/axGGLCa6sVUnugIc86lJxHMUPIP
GNMfcG0w9NEghLRKr/E/g4jvQ7SJFtQyUmw8CcSYmtxmYiV3JVBIO2G8RhAVIsCK6YKfBzFEHjae
GUmxho+mRzD/Mz3mHjq5HnfQjGMduwA93MTY+VwFeb/C+y62mCYuH3VABepqPwkDq7p6RqJOkYRa
3MyM9tcti1ctfxh3ocIDoLEBmDbKdnzgRu1MxBThlCKKIB3C5rd99iljUVa0L5XIWIxrIGcuXi5d
ecC4ID+gw/1upl8TmZpHbYNUp7ennzYq7A2UC9343DvgW6vdjPSjxCkg652iPjJflnSKpmLyfLVg
FqSenm7spkq1KeGcXfJTKGNnudc4c7z9sbCmP6zSKpL9iWdGNDNLgjR8V3VqcD5FJIBU3EpPgfWV
OFZot82v3EzPrFoxDpM6ShGpIGs77y/t56CN8F/6ZwaaAuip6dSw/ksgQHax4oeX6Nb8D4Gj3c1w
Wyv1SqQ0LYa92aZr7tE5L1f3NgNUqFxgeQlEBIkKaJnjFBQU/ZxEQO6GYC1VyvMJMToKjnnrR1LM
y9MvTrDXG4ndM1iUYHPMM40ANl8DgWtD9SeUw9Td656mrC9k3x9Eeo2W2cGgG6lF0Ll1kwPMMED+
Fmr40gBuGfwMq+9my9d3zT8jXz4EvE0FqkgydCjRNs9hcl8YEvFRNy1BTwsLsXoD5pkG28Ap0Q7Y
JjKzssrPRr+9gRTkvh83P8u61GjhpYRh4/MP/zToSR8rKzGtjW6yWTkX/lVqo5hZZgnCPj9vCu1Z
1DRwKw64t+B9mBi79pTIxRI7uVyOz/rS4JfMdWwUOIxQpvR0hajnLuyTpR2WEBFMwCIsf4crtXm9
7GqQUD0aeAxOsr7eJLv5RIyJ3GoV2l860J/StCZ+HPlMIAlg4BD98exXXQg8bT2dasnJFH090kT1
IJTBdJAFY4jlP2MmLEx9mHI+yK4QQJ/k0/hyfI6lWWZsiI/OQxZYf7r3kL5PuIbe8jhRLgx5RpkX
1sljoK9s0i8AEPmR5Q1qtnMVmSp/W3QdOTL2aqKu3pMKcQLT4I1vd3lK4Jr6KAp6pArpDqQqSP6/
JkQtaLimvxvAFptiDHaCYxIGUtnu83+gwMXUQ0Ksi+jETwxz+Kg38VlXr2sE3xVJa7idDtkaHp+b
gfQI3/2dpPOLUNrGAgEq2lp2QmfsXFOmoKCrcH20aDDq1Fk5fzbyErejIJb+cbiQLBZJ0IYz24it
Ws2OQb19AnX4Es2XcHVB5VTc/FDUuGtSk1JcSzSBJrJRxyY+MCOqzzr6fZWkC1hTW+/v6tu3FnDH
ZcAdD463qZnG6nzxuT+cT7MGhjrgWhoykflOxpKw+Zki2w0woo45Vlcvuho6qlPvPE7vTEs70L8N
+LbjA9U+XSoOa71YUIqCj5RnqjmNXyFqYgatsNffLChqYB/2e9eDX1nRcGdkRXmg4FfH4B5vbIao
n7n1NJuUfQK1lo69nfksBOhuqkg908jHPSITyONP3OI0nFIHMFWwStPIkGEHNYu5WjysWwQ4gEsp
oZgU3mkhMsf7/rNJ8mb8GC6Z0ocLXh82N2VgZbrLSqhRfR3VjEfnDPI45CZPhIOY0LxF7ORgONqw
6fCM/WqIPG4/iF1FWBUBWWIUsRzn9EB/iBOoQ6PUqaf6L2urKBPdJPIpyrGM2wmE9kCrnXsw7JOC
Q6mZYDffSL5Q/Lf2TC8wJH9SJEZaiqrBV3jX2e/79gelnltc95MOAw51GKoC/CiI9anjsjYGZ6+4
WLJKemMoOVTWTB4OVQf7RmmKOmJYcfk9Fz5kbEvz/CjYmvf466wJrjZ8r8TIBJrX3bS971So0E+U
NpWI59t9zq6QcxO9XBfYyIp5RVl6LCZxpJvne6XR3R/OG17bDdUqTL2BowRrWuT7934u1dceS4nZ
lUy9ODWbaI5LMHTtFK1lZy0pW+/CjjN2y0Ct4UTeMIIAHNA7iIv0I6xbcfSjcBQFYzwo7SgL+esx
zA9s1QJV7WrhkuerI5Hxj6GE6xcee7rvFBSKPI9//0kG/F4gNNxFodlIYuOQY22cbCQvIeJnD0m3
OgBz2m9zFRxr9DDJNkz/2BqPCDWwkCiSByx/5OkqkfIqisjZsMW7TLZAcQL6f+fe6aoTD/UCzidV
K1W7cGmbLIgxqBahftN+rpqV3i9/cSTpGRSOoDF9ufYbrnUs0LFYRndS0vHCbAQaw9/6mtUOVgpH
PcQL5aPc/oJ3fD8Ilqio38pW5URgb0qIss4WClFXWk1mm5xFBZjF++1m77L2tmgGkpf3fRXFF4/Z
tSfvfL0y4pqR9Zbb2dGQSvnmVyOAxocnyb1ayldyRPOABC6soUiSrCJ8aRwk7TBKHrW5hSANEES7
qovRSmd4UEmMgLJxNgjx6Fx9wHmWVrJccFB7AeCVqGRaMBIIFHTscYoQSamXXOEbo7MYxc7EKeZs
f1fQxaVcNmk00BGArQWwvH4X+BhRuEIm36w19DPMdz0N3Bc556m/y+84XWUXMelhciEP1dHx/U3M
YjOFnIuRa/UWCR+jUIh5mmfdP2YRhso0LJklTTxSRIGZFaDVjMYB5FnfysmV5vRMHra8dDcb7VNP
nVyVGk+jEMHCk22GNbnCA4Z+3tCVwwTz0DXQCAOUUFTm8MNmcO6e1b00PlR1SnE8D9IO0yGW3Yj1
+QF6xZ9KaajkMpWH+foc4LepJ8Au8Oc1W77X/LXCQoCmRWCEMNDD8kxopyp/Ox8PepVPitYDvSin
3I4xVrJWTun+UVKmO10lYWlsSP+Y8ORfQEixcLbmwIHDjT7XYsvep5J+s4Nbdft+vN/0bmmmnbw0
2jcc0ayvBV7JbHZFFotpQbBC9lSufRWGhrblee5lKZgH+9gEjMSrBcdMsR+X7lwc7d3T8AJ06vAe
UBnErW2FTJVXZvUkScoWbk6ev5PCeBvg9tF2Q3dBpvdn2UT32+6V+/1WCKAeS/6zfzeFuLUfnX97
+K9DKicD3yXPw/dhLcFihPI+mc0035oSI0U4TZWXebUWBghUNNFNSo4UEud8x2wif6DuUAPbDA/z
S70NdTqlpH+k0BlLrrOXOSKHvUIHMOgj36MjhcgGNOHOYCGa/UYGYF35nDaJH+HSGP9/7E4Am9H2
zZakRANMKz3wc9U4EPzY7MbbM+68Q4/czMF5Yg7OEGBSdlCFWwd4t2rWmu12ETrWQaq9v0Y+sJrU
rT1/bmbQiWS70iKvobRSIHoofFJrFxL+b8Z4Gyzk4f4rXQ+s3fzU751uDVqoZMQqPnvP7ezT+LUd
k/wEFZeGVktkkTZXLUbN0YkoqGQhd8rAGlMjTmnqGvwdidjHTxMQsEilFNCEMv2XnJEl+7rawIu/
VAKCmCqz8hO+CHqXVfkRnonA/XdSw2wn7aZpQyW8LkmFGKGDzox2+u+tEKNl18EyXXpqrZ0u5BdO
dzp79bPeZfF1qRCbkreBQXJCZ/E14s29tDIKiB9vi2Sozr6KUfU5MDxg8r3ua86EXYVCvBvAkAeG
ovEaorZSz0cFv7Lu58vzsqz77m/YiTRWQjfRToxCapvQXyKa/RkmHlXkjeLs1Gt++hilcdTiTAPQ
KxEAKKSKMnV3Fxt6NdYUBs1c36FDU4XzxEGCJ/CeysWOF7B9f9zM012ERu22cgdwnvF/JWz/7ejC
AGKBfuCGZbAbzX41LF4sYSa+eWbK6axyZIbv+S+vOofPZaA8v0+VMtDFNGu5mS+HCH89tIxBEIBU
l9BVnmpAsiID/tJuPQn+BTLCR39y9zSDnqd0P4Lfg9eamepS1S3eDhqLt2iLYdc1Way/ggf3IAhC
TsdilOiIK3x7o5QIyHI3YF3OpC3XN30zExlL++DRh4blS6UGT2ZT7YvbuFqyztra1knJ1HEi39yd
9oxRbPFc/dZ4pIzUYrsiNEi8YPDRPixnU4WEJomXJztTBSDpSEpLTBiaCkxVgzpgHCihAM+BA5Pn
rMC6TlarLDmwNZfjhmQ2FZ8aQF3wD4+Tr2rNXCqAlxnwPKKhVbblkAJnZvwhmzcZTUazFZHlmghw
cRvAmH5AQHrgq3sAZj0nYELvXUvCHnYLRsTS1naOCxVFxhRKvR932F9lJ+ZJUpAdwORsxyxh3MtH
aWn51jvQV/AGDcUorTmI9O/rWJCR63iXmnqAB2LH1mJQsQeZvNLM7dE4jcIzsP2FAIVOxuMOzgUo
TGnt33iHO2Fj2zY8WISv2s95cBVUZH7qHycb6z0sSMZ4sDIdl6IWJQOzNzyPkBmuE9ccl8YdIYct
clqzqhJR0SJFMbtUR/bNJbnpxcyUKAjCIB8Rxscecnbez5DOt2rBaE9UUscMq/ZN8QT4kXWnTnW0
mHkJyc18/gT2/e/S6uOxSrYdpQtbqXzcttQezRRVbxORp0Sz0IYef+RFvY2zDDzcfozJYkDId3bj
oTlVkTdrT/8buYrhcxBxZD4heHxbmhvOt2LLKhbKZJkOZdR2aoWRFUNsStrUKbe3IsLyvLw/Bqm6
vNlg2/sMhKdCbeNIPRhdctLV7q61Fe9kujqt2CkCdJFpTjVcbrvEnzfKaOiv05JMcYJm5dhuF8NN
UJ7MlYEi9yt2eYTVNT4Ix1focyagEj/Wx+KrVVI0oqXvlOLK//32bqFqdo0cMUITHwvL8vBjYSkM
wWlZcPO03M22XTljrKgfzFJ3DwaDDISgqRdpD1fNEtpS6px/BBKPDhr8+CwV7MnSDRgCR06Hvz+4
tPtYRDfGtEPiDHhLdEx7j+osRygerBxvDJudE29lt8t6+vgU1gfKg595avB6kGQ9OSWQOda9yWCJ
8xlSrqmRB82orc8YKkYdYQX/i3HL9O6tWNoDHQxFDZ/8Hgs5oTjLV7ITbHEXejutjmlQ0nHTNKf2
eiStnQLfJrVCHv/QFTCBhHyKddEtUUihdaDUMPvgL6cuysbLJay6A6CXNqt/Jp8vlgrYGgJPdryF
W2DZPvfs7nTcVKuWeT03dqYqgi50Q366KPnaKUKXTNtxs3oeIgzKE2iVxx869oSoJOiLZTX3UIQI
v/T5/T5sG932e5J22KyG/8TouSvBsejpl5UIX7xynIede8ohpiE7LjImGuPReXQSQrFK7VmHIiyL
KWqW7fN0F0yXxBwN6V59wy/kGmkBYZeqUdwlcSjCpjj3eoHHGk+y0SF9ssubE2/ds/FVSAFS5Ugv
7WnYiABj5fVaegOX6DcqgP0xwxyar5EzBkdnV2ZjQR3+NwGCrTDtiuvq5JSexSdciBvxScBXJAR1
i0ldHFIMNn3Cg+7/1V6KUhlpYkLxTlgKFcXuN7AmPdL77vTQFBFm635Vefl6UraGpFXgfntVcl8b
yWtHqASCcrdLdIxkIQssn0UGDXgqpGAos0TfA88mf4aEqnWhjsKAl6UUVekFqPtqYIbFaY4F8RIW
1XUaOLNKhDeBDr9nv7+l98gaa8IuRmoVHZNcJSaDBpjzm+zUOR19A/6hoOM1U+0IRZX72ljp5OtO
Db+m3ddhiuTdI/WWJdzw56vu+B20Z3wrpxy77WbUt4AyZGFOdjQ2oe9Wu7zzPTaANQvjKGShoT1g
4E7zKjnvdPMCoy67JqLhqKUL/GiWM/FTlImgXRoJ2JoCAgvF7ztvWbDSjHCwWU2urg8pkND66S7f
SmlVXv/zcmYIOmV5nqWS0s3wOuNWGxw4/G+crCpXVJD2Ckm4zui1MloAGbw5RN0R1hdwe+V2v9Qv
GUN0W+og/a6KVsumeJ6OQ3e2WaWNZQi3Aja3CR33is3xuLT32HLllWztU44HBA1CkjOKZ1SMgxSy
JrSZPui+K8BLttvjW3JA3JgxzNIWj5JJXsCMnInZn2Lu5J1+HhlVaI2ju9zmVwN/KCu+RUtmSyVS
lHlYsuTALZl8rCY7dtpovNsueeiNDWqB3SStZpDgtektSyY3IHiH2R07zUnxwgoFtAFSjgojv3Bq
d3IAI1b1R+l+oIjDzkTARyohgz9t84D4AyQe+kpB4JvyJRs1uJNQNwcw4pS7cTtNMd3bWFtPIuSx
ocaTFa/Z8Uq/aaJd5oNt5uuH+UXplEn2SX+6uWYrsD/R0+eciZtHnE87F5DdDjvKXOkcSxUqEdNh
N+fA9YuZrIAviklye2s8c85cR5uJVRkjtZsdhKa31biihvl/VS//bgRGfxhxHsk043ev5vo/A4ju
P6902F3Dn3NTBT3ea8N8Cyh7DsizSHeTNvhLYxxp7eA/hLn3zECjMywIkXOKtYW9De7PDNJVJOvP
y+WOifcSUpSrw1P17VK5tz28STXqyei61Y1ZyIF5yOIsftdxbZG8zCBYjmj+FVgClMxmC0Lk9cRF
VUuibY4RsxrfZdcC64Yzl9js+kJKeBlMYh+czDRIQtEhIxLSwvM1+FdK8wdt4ttRNdAxspmVP1IP
1BJj7WslS7IfyerFqlJFdzZOPQPjdQ1or6Ox7TPgbnuEetK8IfWrZpkhX6Z6mAO9sX13QUwrXk3t
llZCIG4T5cK0KRqqAxvZ64UQrMA4oB3LJGzmwQSF9C3Qk9neBVVA026pAsnvuG/nI+Q4zHTh3F5g
uUP6o4auIabfEO2UsFEPhhgsVrZSImyovkC1byZT9S7aqmtAthA5FkUsFhPzj3fYd6CA1mLFPLF8
IiM3Yjp/IgTOueqSOVOXZeV3wcIWnYQny8Koxoz0qdCSUaqRdadXwf2oGo0hvGeVORO3Gk5fFfmX
g4EGGjorcvpiJmnk2AHZWpLmP5HqfQVZh7muwUaIB78Bk53tSiOChyFq3loC3WU9/hZ7vnJRZ6yW
ZsN7TBi9lxk9BySuF8T3Pb07eGn78CZAGxMBFyjxAhLiGwWQqot81fMjspsgf+i/cg/fPAF5/g2y
BbhjXkHif3LNCC6TXPDOykjcjjId2kA4T8I6PFqiClb2NBAH+a96MpaPH7pPGXcY/YJ2l2PuqhgF
ddH+1tFb0WGqY3RRLwGkM2sJKChumAzHXAkjj58UdibdmQ0BsOdbShgj/TMMKRf/SqHgEWOVTzOB
MOUOkz5WGuM20dm9fRGXCDVylSkvBvTR4MgjIyA80ViVezqHkP4H7PRNZ5E+l9abqNU06IBHREjO
9lcENur1ZfD0tpjYsRLxC5aUaFo9NFtU3GXcMND+d/BuoBaeWOHHKIhNGlggX1bRGcelnLXMaI+V
wpPmwA2jhsA8LF8jbiU/eU0XiukDJXBn+Chjk81Dqsp9hWcvlRgmYmPQtiHPr9w9WKiil+OWMfTc
U47r+crao500KRLzgBq7RA9WPJbsT7mlvFxLV2CbxGwGeEeegAuFgp5HjFUwZwKCmeQMgS8zDz+G
rm8GLpG4rvMsr18BLKiMIU2fxNEr0dF3DCYOKiwRVwKY6D5X+sDyxDIYY6gjWUrL7WMKY77GsZvw
k0aoxe6ykz9NeZZwOAu8sXypTH5KYgOJ5wd8AQESLo44Wh3NrNcX2eCvPbdEyIemeXk+7LEEUTaj
UUg62rHW1j9OLPhE+G9D40w4kqQKXQn7i4XLlnyCC0y8NHzWaFwieutDeq53TXMqLPvq6MThqgFZ
c+4YCZvPGX/raHvhs4TXFu0aXUMltMh7ZXUFcHZuUJwMu+crIR7EhBpjpeD12g5p+NFWN3vWdWLv
I6Xi+UaQyr8k1n2BoVHbVkcJDHLMuWNJz1Wfvk5NoDGjk5FndVzdS+1fHHUviYi2Hctec5bcXl28
IlpCnaMz99IvGYu9OHk6yn9CXVgh9faQ6m43S8Aka0OaWfS9srjjyZBHNvxKRlnbalwvpKWcH759
tEjUtx9Rx++NezhNM+6otTqLe6EKJza+4j+LR26QNDuJrHbyyUIEyI2DhuNJwV7vv0xkbWxwBbfL
iQH8tF4f0cWWlW/30loG7KIZEDoPIEwy+RvgIG+ElGG7FQssiLV9U2TWGcdzyJei90K847vX93FE
l0C21h/2OCNCSWiPndHcuswqHtjSutqxbHQHyOBmoWr5I3/4fbUtwRVVYXpjlZ1RnoHaFEXYdkzk
YRyOXocuTWYfRqdY/fJC6PEJ0CxKguSaF9r9luKviwZ37KzlYlq0KLEQRzUn3HGmyA3zEzqTlLC4
cgWfQiHiuketgakScIeQg8Dic+RO+4g+IwOpKnlBHjEueUaBHJx5GOtcP+XJ3y7p8pzdzKuzNTQN
w9dEqTFVpdgXF7ZsKyA95O4yYLsS4sRct2weiSOBDLgyraQS1EUKdVojvmt6seG2/WBOQ7XV/AHC
N5ML9gnOrtS1GUmb43V3yuYmPjBRIfs023OBIdUsof0AcqZUBnFWNwbC4V9JwraAeclcYxUAjzDV
n7mzlJdNEYGFRv6rouBmWjQOVKxCinYRMigO+KgrHYn5x1Gfs00CoCgjScprQXbj4ApmZu9tz9Nd
0/Pxu+0hVZ1Gr+sxpQlD8+e238XyfAau04cmhtxHpAISfH0OEhXzPoT8Fkzo10Dpi6dksF1QAath
hueZHH2qA92eVIk7H+jtmNY9Zegnwi9OeGK05l6WfXhz5P/fnrTVVE0TJFOV9U9VA4go9Ss7CrL8
bHnqmAZXUoJHjbc1mOfTeBHfNVnEizJUdOdnQxiTsS+DQUK+kZLEOjHFN1iKvUJM3UHLCzQ4keP3
6lvFbbqFeCrpnx7FXYLJvGr4wUq5suGBt9L2gfXad4iY78JlpYJboDFNdZHGsYAXxqn1BTpbLmdI
IZIQXRLb3DFUd5C3txXqKjBSG+x4q7nuUHJKL80VSxev60FH4JsPQKyG6NPniK7bTTp9DSlASyY6
z3x9RTlDcLVodaHaeRv7eeOKrhIZlP913munoSOUYPjZzMBTR1Zo4m8Y/IxkhoTQ67Wg++VhTEAz
vOywtAbKObTjgIZnLS/eGGaDkXQo3kDuNNAIsv7cg5/DCWyq+ax6356sGKD4+nZdbjGAxzbLXOSx
UK/LuzO9Z0AaYdsReHOduoBQAMYmp9x/e5+8gv1Tx8p2ch6pClxmYghu5JMj7FIeHGVqL0xvQSrp
Cf2W9nVZ4KiMAUYMlsOsYXLfASaQ1tjZ2b6WWYkf+99tGnRrSqzZmwE5aXx20tI4ECJv/FCReAS1
8l4Bt3GVw4dpOD6tT1UOCrlkE62z0zHLpRSutz2ey7nnYsa26p9/14a3oUG2idMP1IU8m89a1gzq
S1o+XDv+M5/phasoDEXBc+uiU/qsTkFSAAeqCoYx/wzkJjBUryNDhIVw6pdjKILGwWCeSIY5zK+D
gqDh2DhjA5PqOB+YP3VAVRfsSiRwyfhYNvtEhfOTjEZPrUbAUZa7cMZZhL3blUbJ67571i5FgHsp
rqw9IuXy2gcQIDxV0KnEJPwknkTtJpxCVtuUPp+bHCyF+fFbJOeS2QQFAGYMc7P0cvL25Bop6FRJ
1DmGr8BG8IDfcIKi5/fX/UCNPPiop6mpcFhRbWs6CvvIOJVyTIIJ1JrSG6IKwGVh6XZG+nZ4hGwL
mOQQ+WB4Ag2z1QpTbrLv181GM/dnHH7uAyrll/FppkYx5l9c05sEXJok8aBHfMU2D3ckLLfdk2sj
Euu2V/7OY/4uGCnjpXQBVnMe+N8KTg4lONSt8AZDOzZ/I1e/L0e8Zlv/DBazxilOGXp6g/VJXXxb
cfXg2mi9rb6d2YZXdQR/jVx9YL+52+9h10xgKRRZ6OWXXO1+LmHYEdrIczmCwz4CGk0SffwCeB8R
c2iJ2DuUYECGyasooN3DWboJtfOEQaU28qnfsFty6fRKVR4gBNvWD+s2YTMbNkMHECx1tSGGbbnc
lJlYGC1R5mfhS78tmiAD6Z1Cm1EYNlC9GAtLOjOZ2eyoB3jNW/3eeT4H9S3iPNkdNpdwwr/NTHRy
KA+KBvv9nreKynzq5nH9Xq/i4dbbAyeAYnQVlU4bX6225syxX8riLSJfNFs1J91qYRkSOZa6gxTJ
SrtrO/+JGugcw0AXjFRyoy74ApElAKdJJ6rp6PgNbd2Mc+ZyMRs5UPHAQgKU1xh6cwJACFJ0ss86
mYk9oylzoWhgcrEwKMt5uw9ehDoeINqbitDrfLYePd1StoMl9Sf0WRCuDjhZWY461inan3XzXYhh
8hrZwo7mA2F+OMwrMUxF3g1ocVlWeB+lHqp3rhu+yAFrltFx5sAlMV+VtIHRWnZavIAuuWuJ/YR1
kJRlPLgKX4u6WaKm1N/F4Sg+A+FRUeyTN4bnF42OEeYChm2rFDyZA/yOaewix6Qi+viD5sNRdF6E
EOQNdz+pkAYwUZEfphkLCx/bdyMM+DhlTIyZObCCSLkRNYaJDfKakh7TLVFLbtGXJf+hOrgJ/4PL
LkAM/j62il3KWACJV/XSRbx2YclXkDY1p/DxqbvoprPvZljHDt6K8xe6koY6VaVl/M6+UuVoyL3M
9RFsy7djLqSLO664FeJZZzGF8EP8SD+cmrgpsvtk/lNPGygQnyaY2FpMWkJQE3u+10CpiqHSFXMh
Y4+h6NxwibG43E0HCYZOBnZIdVzSrKy4TXNKdLA7FiPco66FKC4LxzzgewZJ3lsAjRYiUSWjQ5gF
6m336B+01vAf68oRSGz+RRCmJzSLu0o2/VbA+3ZVTVYQRG8Aw6Bd/0AEdI9mfkCzLCGSDVrVnplC
c5o5NlaB3vq4PEwwGgdHQnEPHad9ZqOq1RgBA8SR0kTFKSh9gN0sfja6+OV0N+qzMY309Geej4kU
cdzveWjUY1dX8OcGAMMpongbeU/kk1TYwGZFsOQnopk7t+sERITA4Fi5VFjM+caWGi8x9uedCWnT
wD0MI95bX25rP2xvMzKoWXr7DsG961ceNgPLzlwv3UC7M8JOnYM6VbZgVwhdOvo0bgMesT8qF76A
vIOICypstPhqiDdfuzpyPEZCTn17F7JJAhl2Ncj70a0vv/NiLabHOCZG4Oofiy3/+QBYl6bN45s0
ZogHaS65zAXsTMdrbNmVq/ffDAj7wvXLyxmbpzLsqQBBJXhrJg6is2IofkR/j/aXIe7SQuHDjG17
hEdIVjuQTN5gds1CFJ0s0iX0OdCzhfhW/00q5wLjNmfb22Kj8gIPQ+ks8aiA+AnoqnIeEbvtjWY+
8VBlAUN8Knq4r9RaEgb12rIbzKSHmvv2IbFEgAwU2lG3PLKSI3wtEd/CusHx3Y3v4r5LIE3WfsEJ
cM20xhWFip3WtCFwgwPX/c4stZyK+4wqFTp7+98oNjxa++VBEKRusYM2VCE7fIw+0hqtFXWhJ+rE
cyUtzFBDPpxi7oab8JOoksq+Fwm2g4PONDGfJ4tBxdpzHcGCYCpNvIdu6untpnpj+STgn8NhOJ5I
UqPkNAlakhhTWn4d1bT1eyZTcu379dYxl+DpSH3u1aJPzM4mo6c+2S2gREfEMeapmjHvCNiFSw6S
TBKr02GJcqcw0BrI8UcLXAimKZqaqUIELn/MSvfTV+BsCAYxpV2NmX7Xrn61Wsv5Vz7nmUt+InUm
fjXpQMKL05kRcE4Xn+2A+INYY859yZE5HcWLiTryV3SG98fSiO2QlnLgZjx3dW4Olqf1ENLhZX7a
xyWTSFEpi+/MmJafLF8i3828mGWtrHLxr7MGOC/GagALfNPcHhPy7B+CYvmpdEd72w8PS4yk5Eh1
/Ngx3mRISXuMbwY3J3rQRAGLa7rJSgvAtFpajEfh0qaxNFiMu77s5BUzxh0Kmq7gN5nBbUN4Gd4d
W/hbOMdHMCtse0DzPSMCIeFt8xXFsh1WthIpMJgyZfCP764JOFS+YKs+pDJsjms6kKyLAshKDLOi
AuUoPFeMjjToUHCROR4P8SFaBFtM+/k3kSzD9jyWpap9vmriJkxZ3gvGI7FUtID1Sey8nNAQSFnL
Pd7gewfHlf4fsi8CFhjVn5UcZMxuRJ/e5UabD9r9xSdawVJO0DACdJMnXB3+BZ12e0mhUSGYoTy7
MG3yri5wxkAx8xslgGyQeh6UBCpN0y6WGSLLcBXHH7gMWCvcyOR6l6wSZp8sT7Ap9Zlc9T/bDeW6
QI0IzVcp6uJjnNIfrMeV2llhafONZOQmcDcin2bDVRhm1BMfIaHtU5KfQGhoVof75BVO55JGQ7eu
yEXGcKOVDtzF8w2bia1kkoRb58WXnZ4oiGUO3VdNTsf8vOo5hUBFFR+/pUlEZRIvIKr0Ry4wGF2o
d3A46ZIMMmApnt7h9atI6FyQ0Buw06Fown1yzFxSoJwtNg4Npl+tFEv6xgLid63bvIDrqXmBhMrv
uz4hlQR+u3/oHVi3hdyKe6xWz7/7Jvf7HFvNyP/hDYUHvQoFUa21JN6mP0CZ2Mo5BoOwabRsSiLH
g+q2cOnM7TMarikq/VpGwo/Dw9v1Lh9KABVt0vbInNbBGuCYFflq/YaB7JVw9KOpv01/NKXLwKrq
rbIjhLeYggNKAZnLI26sDFw3R596QZoYuuzm8YFZkfOei6VolO0CZfMG+V2Fq61veT/CzSvo2hTI
BDgf0pn/ynUcB9pPNRwH+soZivi50iXcS3Pf8B+VgLKNDDg214+WGaFXzepjJ8V7Mqdt6vqSNjE3
D/fHgRCGNpgI21Eel4cG++Sy1W0W/HvfjLtRxOnCrRUPw2vL5K38T+iwI5LD3fygIrAHHPTpM29O
gcD/sIV+wur1YtX9GqEiW+5s8a82s7qN0/hkdRfBj+Fsc8GJrF3SIlWhA8Vb4daX0nnsgr6209nG
SPD3VyEg9KrHJLYxzMVfCnEGKO9d/Lx/HdUa9Milnm43Gy0ekF7RvVB+lrmAlR4MrXbZZIjoGT8h
YFgQ3CnP+hHou3XWPezu+vluB/7GiSiHq7BLGmGdSoKakqoF2L+nEMpzxsOotIAkClWZbxoWzjce
vQTKV69i8TCui1TL5BstubZxauJPD4MP4udyrMD9e6Oy6PJm4akHZbIrT3mS9bMS40hHkbafLKKF
K2Yq0UsioWZI9/nj3YiiNRFRKM0zdgM6mszDDHopfWJGMYot/5NHthbaxm6vlF++ZjqoWdtKsrL7
JHbaGcoVEdSHLlGJAom1vljYPIdnwxn9sfM7G9WGL6GyY1CVi+puinSbjrMbHolOAPl//HIYYBXv
Y4zcjTMO1Twd57V0QP2JvAI/8PDFPdsWX0dQ8XPmztRptU/YZ9KWUFUbSlmCBYXn9PhNqbJ783nY
8QaSWivJBsewXSBBJ6kV7d7rl6573lpP+qzLlVupBmeDyaxHap2i6mOEAiy+Nr4FdjpP9S1oVMj6
B/uF0tinIzOtb5d/jeuiNjWmZk/k8MFju4ShN2ThUkbnrNuBjYCi248MIF9OLj7wBBzPHgLHGGHV
Dq3RAw/3d6Ju53s2AsgA4pjbq6ROOtSMVQg743Sv3UguQZF85tPk1KAeeJYiDRjWMYLiTXVKr9Fk
dZSNrdhYAwWUmtenVDb9tsH0UtvbuAdKgrZnyiFbBpWelqIi+ZgKoQhBQk88SIEwFHbk4ITi4PEZ
+YvdRfCrSFanLZ6bWhXl7xru3viKg1mNA0oMUPrn79ZtoSYDYZuid0jF9EseGG+O1dUb7JZodfDZ
N5OSfXpxX5yPECfnmkUWLZNa1lo4tbSofMYfLYqZb16MXw20TCa/F6zA1jWSUPIFV/Np7uzwBZ/Y
KgoikJJqPwuBbJlOEu+jtBbS1Cx3OdlD1V4ZnQkLsfSn0Bm7mK689TAf1JmALvye/iTRJ7eNyJEc
9jVs1jJNnkNCX5SHeGZYvzicPgwf9+0VAB5p3tQgJoa0iIe06zDLXZupvw2pNK+TqXin+MDegEi9
CAigluYNJW77/GYEd5J1RetA0lk5nXzhyEpLWHEZK201RZktij3oMFaOfdfPVdsu+EQwAgGc2kRT
bRXmTqvRZ+z9ABKakuGQHD9xVx0dDLS/TYuU0jbUC/CSW7s48+1JQcpP+g5lkfbhpVPSeXTVHfgx
cdfS193GHx7agh0heIaUQ4X3B6x8SXnlqzV3cXVGh7p2EWzJruZvnMYMCHFtMIJzIAx0EsOWxFmO
n/VeglsxFrMq96YkPB6XpCHbK5sohsAHyNGuuQW18ET28un09z/V9pQqnKzKHt9hWS8BU/SUXS3g
25IppgBTFeQuI9fOUEVvlTiYz7PUjrnI7n7gjJVj2R77Cu9xr8r9XakciSrp5rfoCRq50Dx61EEl
OR5hgh/wcIAy5BAnD8OAdU1mhAXL6p5/PFdZOKOWP4XSuyKyFioJ0lVZKeK0QcwDH9VuMOLvIXe8
8y8Zj4qOgGQf5MLjeKZpGe4y1IJmh4Wg6PvtOlwfT3x7FXDTCsq850cWjlBPV1XIeYbAOBuF5l99
RZzlc7Sf64rDNoCYcvC+j03uyzCbs1sGqejlM2X5HaFBr0/Sv6kxlvBgnZ5ih17GxrQBw6B02JZx
Mq02BVoUs3zfDfdSLtDXnzENeAuTZbvWe+V0UOAmXnvJFX/0uI8LRX0PNjvXEeM/CbeFOMroc71U
3sPf8nln7ppY5VCbkGNRCEnLTuH7kk+Y+Gu4vcqsoNVgKJqjSoyMjzelIRA2WP1FQ8usm/W7vBdU
URjF4B53DJObEWGtYL+zk7uUIdhDtSeNRnKxRr0P0fnHIdSNWX0wRQOsubkdAVwciW3J3Iuwqnc9
oG7etKllkWHDZnFsBvVHzzTyisGaSeIKElwtK0wOKxYHJ8Mj5yWcm8XMJ9O6RnW4PPIg36SzSugR
dhLSJPFow1+E69hMiC9tDb/wwoXWFpro2/CDIlHdHmmGN+/0erad9kGhqTS6xYIpR1yZ9p4JmzO3
zx7xudkmiFhgMrf29oS5BvzTYTxt88OseqWoo6Z21USd0MtwfQJRI9Gmm5JMfiP6Ov10O1aNjDry
KhE9D/g6B3MevTMz2CkIlDb7S51e5QkM0a6Khif2emjn/ryqWAN038W1Y8MFRew6uLwqk+TBs45s
Gry2Nd7yIAqBPZrrVxMKz8bva7haHVebC8Hcc7a6diGwkSuGfvUeeHUCsQovJx4h9sYlGz+DwXcn
YIYgasKEoR7HpIdVvgoAf5cqySvBtVJ90KAn32DetD+kaUj4AGmlA+Qsxs7vBKRZi1CFHUwlLQ9x
/f3O/bRfMonS/gFtlathgCB4ugmCYoz6X91WSu84Bixn/+fZnIlaT27aGWHzFk2O5vZzPUJJxV5X
rCLbRtsGj1yQTU0NjOdSMYpr+LuYIYZDWtbquy2lEgvODqjnFNQzhAxRBdl28vLiaCiMpKM+kejw
VFJ5/Fuzge8cuYtMMP1HLJDwR9Q+ohkpPmQOx839SGsOjp/tnx5ruX7B1KbgLLPrIMkl0YFKXgFe
AhzgHtWO6ywHbjwCfu1cDmIdII9+TdbSDPzCxHd4LlhXplrGjWyvxteJvgW27ZDBkisoirE15RyN
Fe0e6CyoUUDATTylQaaAO7aEABUQ0YC4E6pWJDQ3gSMWd74s8+qV+R9IG/RdLlxbxLGQkdS6WhrO
iGQO3f3NEU5wC7dne15IZxnJwGsY+WjD+7gyGCPuV8HzLQxz9Qvbh4tQRfLv1t2w+3SN+M33MRUt
Vok9qr0ttI0mDTP7zSXKHKULpVm3/vTKo+fkCRoB5wYjic7F8JtRkcEwyDENMVod+WcxqbnXBVMb
/iUT5E0Yz/80WzJ/42JLm6WO+8cEVy91gI6TMX2laYRsL5IqeZ1wi8X054kGReKz0mO4y0NAaVmD
hiLMvpIfT/gBkCPjZZcUK5grgOgquYwRFgki13/dnYF6EbPHduBOFZScu+pEpRsB6Xkku89oJe/K
WmXRWicaWlZqJ5YZSLmKAoT9g2Lhz7AW618q8yRS1bM+5jeq1O44eIB2OS+onNheq482cE/wABp+
Idus0948stSVH5Pn6IZlhaSKcboxrOdIwJPSWoozRNhIa1d50h3jCMkH0EGnufzthHDIypDBIs8J
yaFeefeoyUXFxAvYAnNuWukc66NNoKrGZgT1dldB62dbd/p1PD64aXXH7WavPi+HO59i+LBx0Qkf
eCYfRrKASKCoJIGMD+qsQo4zeUdtfMBOeUm39CPyge8h+TL/yRBjjgH4z32NNUl3BXnUEkXfKpMB
Iz24zq5crHS39evVNHnLRc8rYD8/FeFF6SWY+Qzn4GePiqJD4qaNzpTiPNd7Pn8PNheYh4Tca39+
yinOQ4kps82J5FRksjrGp7CVvy1+TXA46+9dREEXOs+EUi2f7NzCcHACzbM15vmRv7+2T4OWWDCI
wqh8i5ga/wOsrn/M9RY/wLXhw9aUVh27YDvvWcmv+m3WguDZkzwL5cblSJL0P6ShrW3AtRQk2JnC
JvJCIKroGlkZfUg7RZJeK8fXYRNNoVNnqmUeVlBWbgPyZIK1yBPwROX+Rg6WCneOlOtJRNB/dDAQ
SIp701YHd+3YymgeNc8DiOM3f+T9nWjJ9cnma/hqMjK8hha2tX/hc0C7KL2aHmNmlCm9Kk6y9zpQ
58dC8t0hcWd1rj2nQ4hXfWavZ9wRv993AxZQ67M2EX4TRQ8l8xjgPT/pLTGHIzOB8M529Qz5+fAB
2zphUJ8V8ARxU2turknbNhbNyIdU1+ZIq/Tl2yKzKhoUYrWhNjXLr3eV8DnfbEeGl5WmyexV7mj5
HDESzO2iduUGgpi723aVl6++qzouP1gfDQuJ44Xq6hJcKuA7Q9cpWB4qH+0kVu1I1bzk3tgw//Hz
QSSjREsAAWQPEEVEMqeK4bjt7vkwU5mojOlZyhRfgCfh2NX7vK1TyK0CG4RLtJM37eeI9KrE/Tgd
/SEjJ92/E9oV8rQAXLHP118dXjtdZQNbHWPWwFiECoVQDIaGmuo5YR8qIJj9wKAr02SalaPgUBnW
SRlV+EokFXhzLFB1wNkGsPQCiNL2YBf8bRBJSSaFJYZOU289Yy2B5HOm2usPlRXnsMk6DwaxtdDC
6J31/6iPaPDtPgjlJO9AKXZ6bjYVZouwZz2hqPkzeP4tm5zbKhMtH7MS41Vs63Q22DXP8jdPgT18
6Fv/+3tXzr20tEsTQsazfOcz9icP5qC8GgSIfvq6rJhl84Fl4l0ozUYcgNf6kO836uOz1XuQrzkG
89Ssgpas6CG2ACxoZJU5ta52vaa/zjQhQyOJKxYUFbxUQtZunSkzVBQm8W7Fr+rG6aK8UfaE9hmp
OChOOeXBC5qyS9yLe7dKY4J4i/KBT6VDd1ADvsuAq6Vj42xY0h3l3yBCTMxtPcGUXZpWnJHw0gqa
Y2NqprEzhJaOlzWIvlOFxtIDy3gnnE73KqfznPZEWjmapA3MRZzlfg0GDxF0ninQXE8RBwoU1jB+
OLTH6M7+HjybaPNst4wTN61KwIMoqaXdNUm7NhUauD0hPZgxmvd3xtSvX/EafNmXc4FfeZnMY3eS
lR7hzeMXcEF2PMhvDejG17RM0DPRUcLTTFIhAwiu60wwTIRvEbWUqjWovHIoVQx1ug+xXM0L9sE7
4MbaB2tw2Ujj+HbuFRxP6HQnfrgzzTCpfsELM9fCvQQfxuWuOOBZaerIZdpiA+XyqxEyYzFOQEF8
EWKxjmmBgpXTVnur0uVmS7gCegUgGIIRatmySi5powPT2HRfRjoI6Frw6aFZsJ449SEw0TBc+iTL
6BhNlLd2iX4xKvGdpsgwfZ4Izdz1X3XEzRBmUHGk48AsOZuYDwwT9z/Skug+EBZyPDt2Hm6TVkWZ
XdJMc1mwMau/EemOAhwD5Rl494B4CypnJyVXu2sbINuGWcmbhK7vWNeOYFLyQ/leQWz1OdPhlQwe
dJ6/e64XfHKC2guVy4y+0F4LOxg7LbaUPPxcMXFT8FLXkrvGwea0bGJnWutAAjIXBoTvjD24Cd/X
DfWLaeFL4kmwAEhlTCovZRljJm4uxx0nGP57fAamzHaisAdlatwxXVKwwMVeTbzc2UnEHxG8yaN+
532r6hc8US1Lj9bTxblkKoYFsK42C+C0K1jtNhOwGSmVuLXlSz/z9dn7i8E6GZypbg4niKmRG8w8
oswFmCBlUcjEnOeWnNTdahwqjz28Edd0xC0Gufokz5H2GJBaYSFiXFLNv09kuCdR/EK8i9R0aL+G
5VNKug5c+0q9Lu9Nv3wtjZhefn+HpbJ0WW7AE+jzb7/zM2cg3HPKfeEc0Xbs71MnKxGS6etsFYWB
pCjFbvB1i6J2s6a+BSFaxg0R1CqpTp2scR6CuwT+raB+bNp0VQS+8W7L+DhMOpTEXHAnMtfyWcKF
rILhQQrkF9npfuLi/Qd15kAbGhRJpIqhr42A84VIwrQ0h35OvsYZxMrAxE6/grJPbpyY7SEqHf1Y
qRGPdZZAGLfzLhS0uIrRzBX0IkOx0xjm/eZMhRHj+fpd1a6ovSOPfOZAUgoYsf4NcTf3iF3vvKxR
qF3gaBVY5l3YyxsZsd0UpB8iug4VHSelflXuNrRngYtreRgOrDo6YoxdVfvSxwG7ROFkZteONNmY
bx1liqvYiIoBfp3B6VX+TQ7bEsXvBA1KyRGv5phqWz7mEHZbceYxL71ZFP+zk1EPBgv0LV6kpDKn
CwLZhY1zGXDNfdcggBbabUnWgAlegcAD6DQhd08dr0y2HjdHIS/kw4uTiaklGRVT+g2cMzj45NvT
kg9gxornVbTi089JchAqyq16I1UnlCwSZ/mcpTDx8ddNkBu1IkdQQSn9PuHYPSwdRr7hoHJgHVhk
8g2VwvQhR7gzRN85H9ccX/S/G/Yyv0invi+SOhHemXk9iv8nJio0oel4BzAY4JldxsJJOR0/M8dY
z3JWNnOvVFaV5PHGTcOG3IrZZp0An7E5eKk062MC/+t7Vogrq0XTbdSE0qi+3Ba2CdDf/FaXfkOi
Jpaq85+1qA/tpRF9ZbGTCw2ghU+LAR3rAHlcBshfMyjd95dgHMPpMckr5P9vlVFISN8jaPGTkkoA
oLK9DQdC/uy8NetmhcJtw4jxU33i00EoXru1kt9lJ8pUvJCoX3RZl/Ojulp0zvJp1jzq62nZb4Qf
MVwy0k8ljXHq9Hqx9Q+k2URn2HvIwmG1OqYkOtwIzdVhzjPCJvBNWs4fHqgv+NnbNkbFARQulwr0
cPfKt7iWIPU9uLWHgZvPiach7/9sGpHhkKsTwiy/0ayefxDTGV5DozIlA0qalIGYg1PjFgQ2KqoQ
ty0dCOlk67Vmsh4JFfE6Fq/IgRuFmg5+G8/CdT+pE3ur0c34E3IHlkzelQ4OVSXorzNk8HvZMqNt
SqN7J97NZV54F7XEewRynMeUjvHWNYHaIkGA/b4XbS2tCxjCHSk8W5NSe9Lq62talxALEe4O9Hv6
r+JrSCRaJTQ2AeH/v2szcvGGxL1jziaEm1prjqZXKBT+z/A78J6sGyzsPLoGuEWv1350w+NttVvk
+S8c7VEJDnK67LKn6UdM6RM+RLBkuVqayB1jbfasLKW5LqmQJj9RMLE+rJxW2Pl7t4qDfx99hQCA
ni4/mL6reMaGK59TfrhDYDx8Kc8eOiG+MjDW0+yruaG2YKfVBN5WQ1aMWAPSCVe+8cQ2o9h0uba9
+U120VcLx9yZXOIbjwC7fb8ctFw2HYauAfD7Etwu6ef2gfs4rDg6t5qy+M1dMVY2mVSOQ4aXFkPZ
pAJPt4Ssi8Pyq3fkbWHxNXK+EKBEzFLpXB5GAw/BCF6C8q8ml2eBwS/rcscPpICmkDLmv7H/XJSb
RxsWAw9ADqIrSjGcM8xloNVl9+jfk1UpeMN0lzx0gr0HosTvRIgIYkYw6FeyGlKL7ju193SfyHQ8
kdeKPwxSh19a2gWzFZyhHF6GRcn7m6u6cWQP9pz4VijSMnh3guVa21S+B6/86AYgx90gYi21K0nL
uq1GFKDb2wx49vylkOC3UfsZOJ0GF3bXpDbb7havqV73BOOpEo168iv7/M82KSVJede5MwkDd9Wy
bI0jOw9KgvR5WEl0p6qvub8/jIFI5qUYRlnoPG+C06JSn3JFYM5s89pxw8MSFWt9pa0yucxfCdhp
ahOovJySh7gWV8wbV+aBoK3qLcMW4HK3U5EYV8AmLao8zLifxnmP4ca7mUzCcijSy33aickLN4HY
zf5MSip1T3vjwswn7Qjlh4sOAYaWaQU1xpFn0diS9lT+lDsbczGXc78Jz+It5QyiI2+Ibgy5NVj0
xr4zMa09DffozGhVR9h9jlDLbAmqEosVX67zW8mzWI+jmBQfCJNEAgPg8vLuu+TsDVDJfVCD3oP/
bJL+/OA9gDMw81+ntDHXzoQw6hjGyZFyxtDIDRpO5kkJEScDvKwHP87NHVFLmXq8Xm/eafjCDMXU
Xw+MZ064By8wU5Fa8Sd3PYtzbT5uW4+x6WVh7HJfX2q5mrN93c9UDWe8sDH6PygT2tnG1LJdjqZu
lb350VSNsIgkPwdjZRTVt5CISLaTQ0AtXLD86wVD0htmdWFOjpFsNCsUfXMN4lps9KTqKqiGE2Vl
m5DfI6rViyj4DOK6REi+o6GTB4a7qT2k8GVWzlbJ3XflpnqNmlvc0jNuSimBHOaLWECYjERY1k0u
SuKRqfhweDEIY4ngEFKuN5JfLGqi/FFEg7cEpCEmZrnXJtsr7HIi9bN4QyKCGOHFgVgud032O/u5
vG8d8bgKdFVVG+4M5J2ECQogCeZbObmhU0K6uP6BpSRhNVj2zVOeNEqytvXldZC7D7q5ywTqM/WO
n71rt965SFrltCT11RAcYi7GQtoEzoHsld4hhYn0unu/0EfWwbVMuQAjd+Q95fkaepwNw3hCSLAT
WV9HN8KTUphAlc21blH4l/kyi699ctUcQXR0cCfM1aYvLqWwMKFPwZJJ9sPi4czmtGOLVnZDSRYV
XzycFX3h+iNA0R0DA2/1p3KbU/oeApUNtiztaeczkRWcGhFMZRAkXvLwJ660c8LLSm4jYpv1h0A5
vp3+z1kSHZ5k5n25GVnqYkZjk5TGEgWCyag68JbHW2jf0LIYY8IbIv8z6ZdIAKZVZFVIpwwbUsoy
4941nl2Q00BSrYdFq3BY4wGd/1YPyiWvdIaxwYIOCES/F4Dwcg3bck4Re6QsC0ENZiS8cpnQE9OW
hFh78z10Npu3GpHEVo7yCoVLeksQB0YnkXA6gH2jbz8EsRn+SPE0NBDAkf5dtPBGn1K1E4CfnKT9
mf49YQR2lMwTzhOoyP8PQA7vZ6i+UfYCb137bXO/gn5fQtFwa88N74SfMJKQt172Lk6f/JklECX9
WiVHhwTXkaGBmgBOjPqw0iCtsuPO0upoPsVyPdKGNKIyfeuuE3nn6A/bfOFpwSQ82r7iVe7snB2H
w+IR8KrcUVz3RVC2PX60YbrpErEaRcVJ0a49j0W+tuEMYxhods2VRLQOkaPXl2fBko8hpv5nQS5C
M7hOsXRVg9megEnn0stEghWVWhpKVesPT3eCSd3FUUxFjOWInKi2oOAXSaXvjAznvomC7b5V2RC1
b1Gz7PD1OO/sZBVlK1CLfgtnHWRBCs5SHkwhGLue4Lxo7yLRWS61MLkgSoBtmXuQgPU+244Asnhb
Udy8XN027jlit0U7eDz8xAHJFyamYMh9JO1focPHDVqlV2Xp6flD9WmLrxO6tvK26i/8GvNRsqVK
KjPfOoCLWMpfI8aK3wEISd4gopZ5eH4dAQW8A6wNIXlZxPGXS7x/fU7FN5NmY+bNbX5ZzRbSnqav
CaQ072yToeGsFiCrjaUL42euCuLH36pbnzcIvAFZhPdeiQqUXSsbSzyY6CivUASNQeAMfnor8VDh
nwliYZ3ssY76e8AlPZegoPfqEtDC4f5MIs44Ggs/71q8Px/DvZwzGA5snYbeA9QSxwfruIOOcQAi
oMEzHdWtlRWEJgrOTqDjDFwY07UjybFMpahedthyo0b2crU3Rl7h3M6SVIVmmy22J/uGVLJOq+/k
75l0EPn6cBCDEyHqm3/rvQMGYzaqW3UzI4kLclqipAy2OK7bfkhPSIgDDBrbrGJO8HTzsIQ+w9rE
tDazhFH6kW+HmLAcCepAL2jz+VoUM9Gq4AaZkQyJSaqclLcGqg6tyXFrJDY/XV6kQJJP+qQa5CKi
DPX/q501FJP0rBvvqSeixYM98HjMBuxCGjwt3kTZhKJPb2ocMZ3TQsyPnSwjQEy+G92kJEBI8lou
gsXoc3DK8291D4vQBv5cELW/ioBGYgF3gnQX/yi7YebQ3RlxwMWM79G75/O+xXt1CZF8Q+WUthoc
DN0ezIG123ze3vJpJqDT2N/NyBn+mRhmPgA+Ba5MPTTpbyzjYyDlFufheYYUffq2LEpEkdJSBs1G
/uhx6k8iVwUsO3zIr3nS0OzVTZXvyZUUVP4Mq3mTiYn0McJN9PN+NZmbY+wzZCAQPXv3pxvNjPEL
DtP5VEU2nL0SZJGOiK7AD/gyzDH23TTRcvGh3mITUnR2d8O/DMu87b8SH8PNPvM9sXoGFRkEB4LO
HZ40/8oURHgC7HLjGblpcUfT4PNImNBvqhYXARAqB+Zx5Zoau2Uhj8IGFg0nmTnzDWrw2V+G7YjA
BncamLJthOw0KHZ7SvUOl4wVAE1LgfME0gamlkMvt5ku7cv41B3wA3vMvsVWyllZPUpjGS8E6qws
ybSQMa1InP8EyqQlWXJhKUPrQgsK1GwaCXF7oidiPy6YPCN+Io6+uq9KK5sTeYCcomz4ymk7h8ad
oBvu+Jj5p3GjkG3yZzzp7R0N/8LwCszc/J2k5TmHlwcr0svzXjigDmXbeN8ZkfD9iAeLoWaZNFcP
X+LRxooEFuYRYysoBbl2x8Enzj0lFNSaJVp3Dda33ZvDeQyLNj3T4HFYabYRMtk9n72wMzDM3xE9
tnef446FUcHGEs8mnUbE8sFxZQ+sw2NIHL9sVHkX4SuDjsLP+a5g03QWSNjL/IQmZ2l93WZT7Pzf
3gSzXB1SyUOPLzkNDDJKoM7k49K6GP1q0O4ci3bG/3nQ0ASQ96Xy4hadcqEHm2pYVvaOR7iTnsUY
QABzczilQHf3S6BeQ2GlF4EDIdOdvobXY2EBx5WgqFduZ2YYb4rsdQzNvj6kzwkG6SdGbYjIkau6
/5DAMeNeb3P05tkNbKfQMaopU2zlVfHvdrytnKQlS/sQTWK+V3ZrxDTA3Xy9C5W/eWakksoixsSL
2FyRYAF6M1RS5PqkrTcFvSlDqRVoD0UDkRneA2RARzQlbXKMKHAOK6inT6Uc05W0rDRaXt1piG8y
ydQmqa2BGBzWanOtEziv5Y3vU6W1PDS21oInGF69D3km8+GMdIFigjuv0s1szggjQTwTHS3Z13Bx
RHaYoR24V5TLL+D+bMChPeR8v7U/yWHOoy6/oh6qg02etecThlkzy+G/LSmo0YKtWTSGRBO0nMnh
uydInrYxAy9mzUG/GApcfjy7Laf6v7nNIhMR5p95xlwmqY1eBDLwsf84sZfjVFIlMcpuNUloBaTA
HZSCDOCz7E+5TAn3XjV7HYwBo3HsgWUusa5mz7ZAKWuTWoqOy5HuESPSy8BxuEQp5cLPjGqhWpcV
T42mz9JXD/Uh3iM06fCKGwMp3rldA/frrMlsml0cyc0GxA5TtUQhzUhEkWnihK5vOstQWUIRlC0P
TSLvGbrNWcWL8l+zYdOFubFhyW9dhjfon001IBGF4ClReQN6hGFXluMIEQKbRwSCl0WSERBGBn6W
DHimPzkltoa6wAjMX35rgJfm7UfjOgDgcDugj53fOwXlvoVgz/NPcwdsxxIuiyppvo3ceLuoztF6
Ipf5uXvwI5tIG2fBCq6lOPqzmBSW3Xr77i/Mz8Z8NaIO1nIUlTg/bn5yelkAL5OtoUJybjzeM9y3
+eFixuQconm6KrKMWiUwTKUO4yzy+dL2zCCx8LA7JJ3aLyiyYxBMtKZFA9VjabhfzZ5sTWF1odt3
nJNft48twLpQv41h76tCCjvDQEkAmvyFziUJq9yBwEtZoToT0dc/xjbbfTk1pp5Dmvzo4wzhLeC1
zhNxdWysIhwcl9Sum48VL5wnrbGDRoqe/kjrRKozHgzeQ+5jmYptuMkWOgDpFfoLwqvxuhpqKubr
xdDBNUHbRVRSFP0UN6U1mG9T2rwkcTj554Nbq2Og3yTkSAD2ZH9wYwa3uYlEpLF69bf2ykOCEiqE
5azFR4hf2RsiQHFvcIoymo+FDXFiP2ryANeYslikvOQ7d994ewbUiZq+LQIEuaOkpjEjbl2IMGTc
RrPlb2T1Pb84GZUij3ZNol+L3XHT+kpZla287k8y3YW0UaBxqzL9p6+sydvOO1+gquBp6j1YLVLJ
f1Rb19+vHIrwkbpTh/0Wmn/6gXU/c+vFEHXwHNXCMjTF3LhWP8eU1BaIGSCtvosN+Z5wIoQ8RYns
165v/pVZM0VkntpfydHP04hVgsmAJRQ+zxnz55wBzxHrZA7DU0Wrnor4dLbsVX/BvBTh79sLk7+y
QsysQnTiIrREiShMkqSMaPfWcvZjoolW21o2LNzyRapB937cFNpHpCxdT6DBRyDi6J+z2w5v+NHt
Ad6eyeGj7I/mwpvTqEt+NDVqYBsA700B3dsKgAARK9mW8Moz4bR82Uvb5haViX3iuljUyQB+zF1Q
duAK+epcLDiXzBfZimzZjEPQo/6rh8v0fV0cg4o2jXyBp7rUP3d4KVe1gWGvBPD6MzxL232gqMkA
HLulf4PLiXvUBLTIl4g6DLbjc6Vliuk4vPUIM6t+cypQa6wgMdA5PbtgVePEH7ZI4MIgInI8FUFr
4D96AzkhQQMiGS0nlDuKJb/Y4xDSqUA3RFG3r1jtq348ZbOHJr5bPLhz1kZpIlM8x9A88gcX/NHV
0SZS5AFPg0Vsn5Sl3x/tWVvRoryCbscowxN0BAISozTCB5aZaPLhnlmQtjT/usVnKNGNmR4hm5DU
mB27ldijZlxRxWKUaP1w1sSh+GNRLagk+0fJHiZq6pX4yKhsob1MEW9bl+/FrSA2n8vRjFim8HFZ
0iBOMMx3r3Z7LY515d0hL/X+uwCKBqWZEW6yCPKRU8/0paBKAvZm0jO40YSLYZtR8W1U1TDKeBks
LCJasGU4CcvX1dsy/w2FiqxOkC09ap6dUZTss6c+8c3qmPLaDizH3pTBLMTPWBI2y2aVPdRVQv31
EqCIbgqbOavF9zsEJ6KSRfC4M0Q4FAMVD0pSoeEWYc910bT8z9lY6nMhYPkKukP/p/+f1qLuKztH
5nFmQmr3T6m6WYjxoJ6etC2YwBkEK8xWn6VqgdNevoDK1we/DwnMySHJ60xmWJNqzr+PmYk3U9br
xq/v7NKu1KTTHiBvcgW8Nx8MxVLhUCeRCzeqEzm+x6DCJZBrG9RseRvquAbejd2z65IinjqwVTl9
9R0YAHO17wNA7uAY1JaS9TelQxd+txd5A5pf247RRkyxtfdrcdUajlakfnYKcuZdDZ/+QUIZoPAE
xploJ4LLYmCoJjYXCd1XZAZjVQMvMo9ZDXbf11FGOALJi01sXcLjriW2M4WeRr5gkxmI2FQdnpat
tRToDZbHHfat0/r/6h7ecTjpnp3C7XqzSOV8odwn+gTcJVYAqfvjnUrZwylyMQUgs3oxPgitM2s0
hsVtzlj8Cgp1QkR3mCByilLjyzMkuf2T8/+3MdcsB6A+Zj1S76iZqb/fiOHtJiwuP61FWsMax5jt
k3O30VlU83ArLJ4alddCgrtEbQCbs0LnNqXrY2Xxw3/4Dwh4enTwBeLM+Cs/q5AqS5TZmVYo5BvN
TkmAFI5efPwrsjxumYrVVmp+Xs8j/xjbwJncZ/8fzSXiZLDscuYq+aSXQQnRlAsYpyudjm0WJD8e
RFD2lMyZu3p0FSWGR9AZp1Xqyq4sIFc/waWjG6xDSt3tE52o1kjv2NBFcPtYOFngvFMjIjcJBvhn
c3f1ZrF+6hAl3LGL/UZV+Fgon1FEoZAp25Iv6NfAQ9Ro1DLORNVkOGzDKGKL9dKuuqAvsOr3J7Aa
ouaeL/lKWwsgsEPNKR+DAQiuPg4VOXcZmXWEur/pu3Z6NfF9AFcqMHrgt4GVQvPifNWEKRY7W2/+
vuoQQcEMdQNoDGbgJjmJPelIgNPB5CaSZJ7d5VQZK1brDLczJpToXHFhBxJz1PGkX0OF0Fn+Tmuf
TbXWvKYor9QV5Yfn2COz4Dr1rLcWzucfzrU8ey7A4z22yJS9q6RielQQMgLzhXbw+6xrWvYA8OSq
3w5zd8EzUG0XOjLzaGX/wU6C1kou50X2SpnXs2KA5351T3OES8KuW5MfzXxFJkSbnb10cxtQRb9e
/RQ9rQs4ngLsE9ujZDVPvZlzV2uA5y3TEMX+YDrfNEGtV1AaqkPYmGE8FnwMMYsOhqMZt5lJHo8y
P57f2Cq6sgC+L7NBk4TmtAxfd1LcJwh5E0nlyrbz2WiiWVtI56y08mzw3/1lPqpgllVDAOYbIFRc
SXUlolXSdvjMzMc7x9rLFYmWTZwen2ZFfYPEQJOL6wsF4BPwNmAjwLkII5ROfjSEhncQlwAc0cLj
klvJ/sSMz4DnqBk4iS1lU6nUlVHyH5LVMRVyv5SHj1/9DL1B9Oth/OAXd6VTWt2p/tUYaA8k4bVw
BKriAa8O8TaPUPvma9d4eWz7H1b3rzfTnnCBpm/imRnyrYscOftKLZsNkTXukSVMws/Kg9/ehPt+
J9H8idytob8Mb4btCoSqlC92O1hyCgqxl02oe6n44SihEZ4rc3w68rpBnGCq42AQPP/4HPu3M7Qm
zqXNPMBmUiQtW4ZEFSlTXhS2bCnbdkfgmHpREng9DIPLIfxfRxh0CW6gPDCBVQdUelf2SKWjvXpn
Hz6rl301Fm5Bh06W9tkWBWbl8c+vnaK4g2AfGpEm39oND6/6rqT+1qt8fECuVso0q0a+OLt1IwOk
EpIOrFhf3adWKW9s7zfTlo1tybt19GiYxrOgYmFDzDTQ+Tt0vlBoH6oSLFQ/45HiYwAPCUX6m6Ie
wKAWu7FvIDc1BxFuz/4eagg/S5L4A4ShHvPO6y5SSgfckV7/VBlySujLCPZ7ldo6FwlU+gfJOdOr
iUryZuDb90TU00g2Bzpbc6R0uQHOyGSUXcfhiUxGo3NqDOKny6Wugx1YdyzEse5/X4rzSVQedQzZ
B4xUskZ7WtPN2TrXZzIjoBRl5yhkUkz05lnJbsMmisy+IC4w/jB+eTivkcOcPDfv6pZJN+lMlGXX
mPdiX8WpQXZzwg6NS53A8MjxsXKOXtSVdSmRRr6AoV0LdrSg6QdHiUZuawravlv7SLaBdY+67neF
cxMMwT0tqwMlCGdKnf//bn6kQG5otUlwgFgDsnh2feL/LJvRcV+rszvslTNcQXzCwqQVMUUKf5I9
1cdkRKwK1ivGOIQRY2F9hw81FUMs1Y1YZ96V197oihOxA129mpqyaKroA4Iv+nC5lC3Z+Q9yZYAt
wmzY048qvXKEK94d80/lGoDp6c5cT5Sf6NOAEx77qNxT7REovoVPdlulQSsAUScQhTFMkszYAhw2
HGWkwDV7E0BqYW2gBvhHBX6ofnEIRTnXmUMEMgWkr8pL/3j8TUTGqguyfsRleQaFFa5de2uAs7RC
QzYxNVDJTrQh9Z5+DVDPdmksYd4W+w5aInAr92+L0cpsToZKeI1WaWuzf12l09RJtUo7UlCLktx5
KlaOL/JSHIyYoiu5s6Clda9TsBXQxfkab8zXJQ4JN53i0VjtLZbQ12NU2gdxe8DfkZGKrelM6eJM
gbF3EFv8IBZJkE9kvrRyaxvzy+G/rtNPwj649Cgn5zn03JSyzkdMx+OnleHTTokYOvGZkSmvFSIV
wAB86rLLx+xQONSe41X53hTQXDoDQTBcqvlJtrtPqfLBojq+TPk7P2usIGdR4QPA0+vRQ+CHeUuH
ZwvRzhZfXQIxWwbNPNZCIwK0mz4CCpHG4VRXuwDeB2qcPPRVHF+YITlMIZhiyCmgofIvM81gFE8r
0S9xD4jjevLVhpZ+E8iwVcazGwKinGfoGQGOpLbC6+ZDqSzlevNiNSwYc/c6GfqzIAItWUXUDPYB
wmbYPwXG9fZKZXVTxPDWdx+EkZeMP24t3sFxF+ZsOSJFL89/uU/vlR3ERvQ4MbzUhvMamyDDJH4T
4iEGkKFGYGZ/pb6OEXK6324TEo/OYoXLflEUWmdsJ9ajZdNI91HXV74M7CFVGA257MqUy9NGmRYE
vCA1oopM58XTx7gsXyWsW3NdFLB19rHOdWueTf7NIC/BhzcRZ2z1qia7+8FPQNMpo6Lca3jvT5zB
sG+53v/9J2J56FGn8rCbYXjUU8wY/iW3XB/NGrebPWj1jW52kVdzUtlmPWi37DOy9XQoqMheTfTx
OHnesU+3jZYbEQndsaWyK++P9jAVFNGLg9i7GmX45Rw13cEQWrMY56yjYoiIzlLLhkrS5DgLIkdT
tP1ppXX5lYPLAnYEvLmSRt06NDrfeZyQWJkOzZqsUfuZzsUAtLaMRwxzM8naLPebV2by01fSyT8W
yyIoUW817UfTfi0PdEJ8fYSQTKKaDVfNxC+iv3DQA7XUINuVGYOA+qewp04m7Ejv9EjFrXiuoq5b
e5pwuXD8saISsrSoj3pQ8OodyrBm86HX1xcfOIMdSOlYB90FP5UN0efMWSDyH8+QRhmjnO6XHwBb
r4mPanvFS5A6bLpR6vk/f95HGC9DqbuW3qgCJy37+O3SUt9fuDu6EjnNXIG2Y1i1F9gloGDA82rT
jIWZiwKL8x67KVthdd4Th1seFGeMwKPxcWhMq7wcrc69F6uhCvSVVlJ+0G9RBeibT/111qGQkm1z
IR9/Otfv1mT8l/fN3NsqZmZ1svPUF+wZROATbtCkTF0N5bBCYSysu3SRIT86+xjX2bTtwrJtbUW2
bqLX0KU+XPwQN0v8PdtcUChDmPyhDcarMXf6SYsrMeIFWjlRoiNvf3R5oQjSGiFvSH29cEyoTsz5
DHOhqXAxkd4JytVnWpyV2iA0tORj7lL5Enzz5fg8oetdIGD47FYcLSO9enGtnB4Q7vCo1LRzgiAj
jkDHResmeTKjbT+W9aDI9QdBdvRLaFMZgt7/UsmYxowEdYGWsHxLkWWIfTZKaeKgfFsLSn581Nuf
Wf8iNmWlErnYgqS/TWg9b9hfzTGL4Idaec4mJy0aWZM4xHiTEHbLFupN+MRjsqJXHasFjjdJ4RW/
LlbnJPKIPYx1mbh0WHd0FGGLXJhUFjwW2S8K7GdR9T2weUezYGXNLhHHbnJAwpfc/HOhhiRyabiV
KWRtpBNZGMQRDrVdvD1eWNye10hFupzOhdUD9ZPzv8HR6jZ+uDPkoujb6+E9oaK7OjS+DU0/Opzj
q9SCEspVxHf65xR0qczXKYdJHVW/XNEt6xzwfGzbUtrsXGwDCoOvkzAq4wXO2a6zhY+4qYk38RuM
XZGNvH2M5tY0sj6WBpUMM0pKPhN3+wm5V83doQ/vm8RIVsWgzbL+pY9CF/O5IWdbbT5jQHeFuHOT
g4cqp/USUq6D2R+gJXR4D4aY6vk2tTDT3kNvb7L624//ekXoaNNaXqKCnlRDb65UG9TnA7eYs1CX
0Zl0rR/BcSl2YzWLytgZik0clpF51vFILAv4SJ0b+lchc3+iBzQEnVVk5CqHy+6IubJDk3Pt4DP7
CZrdSphW9+0zNzXMbkh8ctKD1eW3Ozs/DLKOhY7HmKLmd4zazRmu4yQOAFJwy8Jv0GvpkT8/uv8J
IbhsNwXqqOxij/H9gdusWuk9M1xF9HW6HuB24MVFXFOkTdvtNBpS+vvoef3JJYsidLNLyLBSnmp+
MxCq9ljN9Mshiihf1vQloNzol5Z2DFOkHfYFDaXGfBtznnvb4SrqZhMgemRw5AEpQflQa/3+7yMC
XFARScCH0rsaGq7AnXM77pB4/JKhAVGsJC11hBeisoDIbL+zYI8CGA36tgLvHIK1Z+VTMLKmPLPl
7aA2i6F4HQnWMiYtVliGkH/i1x8SSjEcRxMY1tCSY6fFH8xvEQclx2Yp05/3VKw/aVLf0alh/qm/
E2EEVTYlKBh06TO0o9EE6bNbCRzQ0zfNx6NIJSkF5qavC9PaKUaI8Fit3DHCy6iXL4w4QdYEQWSa
umHWPur/zjf7z88bwkXwIG49wilASaP8kpmZm6+TLp4C3qM41EGUrOK+pCT1NnjnRX2nHcm8wMU1
deDpIMWiHolclOiYY+iFh7cJuSq5vQLGwTgG4LYpz0U0de0jXnMQ3RYG4uaJKQ0Ss3fusNTFO/EM
gzZQWbcF1DLoW+9uWlJOQ0dR/hdyp1cd0amRoiCz0mcC5BjV4PufwLwAFtpisjhUF7m9rnCMNFDQ
4Ahh2Y9UfwKh2mdgihIj6fppM1V0yjeVH9dppAZi3Qm160io/AIyta3jmKrhHufvKnUnVWNJ+krp
v1fLEf2F4SHKvYVfHa+Lq9ESJIcODekM6qG67ttsOXxCh2Y8mjR8TbRsaq/FaR6QON5Mdczw6vQW
x3qh+miFK4eVL3q8fvy/roz2fJ47WyQVUUCyWTmIIvcjiukU3kDXEFMSBP0sYRyf76UB4hhb2f49
qUi//3mYx0CKoKsXprLcI7t9yZHafPAqzpfMcif6+jZDZOalGdfUEOSURFn5qRo1Yum7D7eD32Vs
ZG7TpYVFh6GnpUdllIKGJ7AjWiPcEylIA8N7Z4YYObNHFW1i5F9DV8ecjdxNgPviE1v0Zl60Q0cs
dl48BpX4ydZEjmpE5WSF2NOasEUeNAUXFRM/H1WZNOcyDoGmAKdGb6ejm3DovkpSedt5WKml7qsE
AZPoOzuigcNTDfRywMzOAAfkeqsBZlhU+bR0Ibqy7hDF/DJGNrKTkkjVlN6bRbIINImSl5RSpGBY
FEU7Ga7wt+qDuVAzdyBPzkmNYQAXpHFqDXhFcqETpTadVeXOzMQ76+ijhxFwOZOj8+Ak6s+R+hN4
oVtJ4zLH1pAjeVjxkJeBIevXTQXAk/Jq1U45Az8HMAhqcJIzcbWLV75r4StxHMNSwNPe+4LZkrPp
j3j4r9x2BTcIAiwfLem+kn+7CUY58+FE5zXN8JObhlQqhKTs/umEaZ1FG0i1i5kCJCzWOdLSuaVB
uuUocAKTRLzKxpkfr9bFZzIUp+pGNpIcIgSj0VtcJEYLLrs5AhHaFTWlxIuIGJiac0P0uxjXGfPp
1qWWmQM8uwwRVWWRntx/1yBkwGK60Bai4xs7XrhwEXiiaa3vkVokwP9ywqZvQpJ+uO2vkhLGaT1L
YAIubkO58zxHBWJ12HZy7L1i0Mo+0nnNbiW8jKhDDtoek4KR0FZrky9I6XYY2Q1RRQZQVDxmBLTZ
qNyICCj/MEF91Hzdg3Aa+WHGdkRmZMtat2Rqx+1X/Z/xusJRu5xE74WNWsWwSoXwRmKejgqkbWA4
iIR56Qfz3ZvqiYZePEf/9PYKoa7wjhsgnspJYoU+pnNBSPRDcEUdk9sAnELe4n+prnP0C1zqjT0l
ws+1hNqtET2s/a9iPEtPXPiM3GSkcbKiGE3yVW86u4Kf94ESe8xdJcExHGU6mGNCPlbErLJnZVei
Hq6zXWbjkqGArSI65/ZNfxduL61BE97XRaXElwCPhc/zvcOhOcEKiDidu+Agm5T5qSgo6ghlGOBo
zszJUr2O2HdmnmEBKRoI2FuNPGV1UJcgvz0/7FVdst+F1VthZbcp2x4YHvLOHS3ev66j8mS3Z29f
1aTbS1ywfWsYBxgc6F7LiIXxVZbuLVPnQPinkiPll3EF649dwdmx5vp402UcvmU1dxpk5eFyCKDU
JrB3gj/J3vAOyUqh7q7xdGW6rZDyD8p7ZF9rV6D0HzLiwzDBk/yqJk97ZlgPCjsXq7NJ5k4wCkGs
m8IhzjwstzqXLowQoMZL1xEtMdKB+QeCQqve2p+klxLMcYc6v1kD7/sn0ear9CMe7j/X0iYmsr+8
Qs0PjnuSo2ay4MnRASAHVM0mKeWIf+lnIHTQbujdQSKLXwv5ptd5HuVwn9gpYsO7/BSeemTYWRSX
etMLnqAAn3ABjL24yxPMDc7D8U2BjCK7YypUryOqhpJnQRrSeKX0bfNYATctGcKa93X+3Xxz9mN0
ftOYGbzd6E20ryAYTTSxaIzfwvgmVN47MOEDWJ1De4ez3p6stmX2UnGKq9Xq0RVqW52sCHrmLkgu
0zM2b40VWzCnZWf/Y16PRwlrS8O7XANi4zFwkblnJvhj57SCMd6Sq8Fq694r9cDYS2xZhpc9VHbX
5L8lu7UrKaRXMrEs/tIFlPTEC3xIr0LjQXw7r+Ubrd1VbBN13ax8nP+Q6K3RYOXADcRCaawrdtth
gWmrAk5zJP/m8YwG1dXRSbcwEIMOPCGkxZX62SD7gA1B9/CBOLACWgoRk4xHdtRLhSL4jZtG7uAv
0WJpjwJO6t1kkWmPOqLASPwKUnfYlM/LxPheqczQk2LM0k6SmaNQlkfAJLWNI5aX2I9VFzj+Oc7L
enkFQgVQTXpvMXCsAezX/bWkhB/sHLnX/uTPRaAqJ6kPr2CYZ9osi6G1/5MdJVhbUCAu3D6RpG4P
2OZCftVtFJ7pt7oPaOukesDugJ3XvCoY2FqWMpAMVWDSCsU8yOmlwd6f3J93OqfbkzLb8Y9JIQyp
9N4p9kuPbECKAqQsrwXpLvCFTGCZl8967W/xUILlbr1lBlIpL9hqVP/ou4Ulg8WAnNk9DAEUTJj4
QfHLw0D/oWmoQFnAzIYJa8ikb/JaArEUvmiYu8bk+awhwvjUPZ+fC3QoBlfsWhzIWbCijPjVzhFX
W3m2v3A9hDMhDZ+C5fTH2q0SltAVW7T4ZFGfQxm+0ykAeF80YjLonWIDF9Gw44ep0uTDuNt6ewCQ
moTD90sSospPf3tcnqRG4IAtcG3tl3wx28/MnnvZ5plfV1+TOURNb9m1MtD1gcaNIAh8E+bmcQHo
51MOOam80qYM28fg3vkJb+1jo0+u6nkHtiF4cDeS8Vh29wA9+qKdLXKvUscMSpXGOGj4QOq2sXDJ
zThZQgVlIgkPq15YljzBi45LJou5MDlhpZqCP3jUjnfGJMqUkc/FV+m8GWROZpZMqRHWnInfRzQD
/4DUpyQwvXOSRV92OzoZwCmy3eOmPSOKFXME7pitEchq9DtUSdNqqDcYEh2frPQ52KS+kpY8aE3s
2rEZqro7x1ThvgT0IvJPUp6F+GDR+tjjAe0th29yM4/qC1eXkPEy+78WTNvcOL3M2EF/pSGhFnvL
OslqbJkvZdn254fIc2c49WZmZya6lZ3mYO4KkGv3eVSIlKrDmieh/MME/hQOiY2UIMZGy9cAyZdN
4mQ5Oo3cI8e7I/FgegfJaRX1ERwj12LGlrO18YFV7LuqIa8pdlEwitl5SFCrFHX0uF9+dFOT4wWv
OB9MdZyrz2EbRwLBS74RE8SGnnJOGhHz1gf5NERRmfGa5D3Mb3eP0hTA5fiK4tkbXSYFRhk4lHR+
aV2qKVuRQIhNIX01eVVAwtG6FjsfOk3J8il7sWWLy4JchnptZZnk8YGtfU7zUKrwZ506N5YXms9M
wuGT3M7xiwUOFtGFSWFPG5WtNVH7/qsBi2AqN6TnO9OGrUGXYrJpH3pOIDkr1XZTTUrlA5lEmLSn
X3wQEM2ADngUdP8+dv6icfBGowy/cul8AUjrViiujmRckTHX+s4f3PeCk8cfnxqO6a/2p5GJfcBb
dyrz2HkQL5vrybi8iCwKdQJ/TRki6BDX96ulQaieysvmDgoVr5I9917pLjR5J6uCk1AcnJjYieuO
zqXCy1KtPqI/3JxJY1+d3PC71MtRVXzRLTc1DJlCiH4p7mJXhKbw16Nmv3+afH4Y5uTt/MJMF0YY
44YDjvpSaQRT2DRjh2v4/NkRfjkhqGF1mrzvPRNmT732UzuUJEl55KuBB9jC3XAVHOJPXH9+cp0p
h/IJGMp/v1EKXeU9kcxEe8vH8eL5xGlDcb/LscMwng+rQmdt69m3X3AmSUQ0jOnqF2fYnKOgF2BB
T22f2V+f+XLYCVYVj5+FDtFinmSSXpSFqumnMw2IIq/GDiHiGyOOVshZ9fsor3YB9v9qEjo9BOhW
8eFYo899jI2RSmfN4u2IFO+YqXTeOvdN6xjh2obYs7rH7b9Op+0yF/PXJxhYEEx1q+Gl10+KCBYm
PgUJ+MZVktMbZ0TK6zmZHpTrkacNKhXAZeSkTCPAqayWyz5ecVy/7JPewfPmOy3IKJSwTqapD8CE
R5NzMWtlq4AVJbTvCZyrgbNvVOED1CofCqrtvYLWtmlH+1r9pE5IY0QuHgR+0OUD8KwhsdZsnXKi
WQhmIW1lGnGmQ5wGxigkVprsux5ZscbVdguXWMxmF6MAWF2kIupMHOUEJQhiJhRVOakWbzUhndO8
gpjmScD8EzDsB8iGN2vmbqa4XKjSS8n7IGrFb6MJHCGm1rGZegGgoUDhhhoa/uoFM1y5s99YA8yO
9jzsoshDF4GdqJiORUymGnNPJbOM+Pact3xK81VzaokajfrxuK2iJiRO3ZgY0kHHzgA3X3GaWh+s
+CHrl518QHMhQATD64QPC9et8acP9p1ii4hcyLsNtWI3o2XR063jtaELtS6iqz5EQag1qGasYuGC
wNUzPOwW3XwSEnT7rNoaTEX0x9po27Wm69tPIGW6jrMrE4xFca+WOQV/pzMkYtzjFqfFi3XJQ/25
NaTr4EbmT7DzbQ3BRTGNessCcXdX89L23RdOYmLm0YOS/0yoPIEuXSvZk4cO3Zg5uorfo7j/x/7A
4ALDiH8BLwkWAfKayAa2sx6HtrItD0aVCCFszi44Sdok/tji8NsOB8+Mw7v8purTqeZClaGejWAH
irBxLpGOlbXOJ483NKuaclvTuxgQBYdp9pyZBJnEY8usyFC+6YO8c9Yp6j8+XQG1VLomJUp8ZUNM
dwkGhzxjqKbRdzd5Mi8U/04yc24rbIaBjEOSRmxpQ06aB6fEOezHyFDfnR7NsAEu54ckyDfc5j1r
FbQWmLYCGL2hqBRfXzxABYNJXncsRTOBc/LMSw4id79RrPl7Lue9osseNNZ+YsU+nqQA9ZXHMxii
DWGNybmFw0k9mj3EbUL+V3Zlg+OEQMxFF9KgpstpPNBSoxEoPKbgE5/kG2vqf+Y80V25AsCzZY+o
lqy349BT+jh14kuqVVHSqRqmSZjGVcbEIKVNulyKbptWViql47ydqsW6Q3FDwUsfJzxwa9tThsG4
QQJPzAlfaUHoXy9cnm/jZrQfU0OSHqV8eLtU3MrqGzw6SxW0CK3YWlFdjYRiEH3RioPI10BpvlCF
dvSrvSwh7y7azDsyIn7tUSI2oJppfwwplmH8i9GJKNQKCkB6WETNXoKqLmWO0v09be+VLdROHHS8
lIoJYMBsEJzjCqpUFVoG5yIrm4EFtdF5j4xZOJ2EsbXmrrlj7rZqOcOvrJEomMFQP5yxKHv1qFO6
RKO8t7gHtMLEu4kzi7/XcYwbOuLSpeAbteOGxbbQmATe5XG1V794zyfLJ8K/WCFLA/7vcBuIsIG4
bjKkS+TC+Z5a/xSAMwXRJ+W4p0VTCfXj02cjN+OcOWJ5+rWhfjXlluooDpSRTOrWlVq5X+4iS1wg
rV/9y0WqsrWBsepGTj4R8YrhWTEk7GM1EUiJ0MuRzaU412Tfu9tX2Nfjo0DuzSpJ8BGpg23sCK+3
EfBrdyGq7JBWd/5wFvdYAAp7z3x0LjN8OEcbtzYeRvII+ItzZuDml9ZmzPmFgS60V0GnpEpPaGik
SS92pgfXwA7UwMx9hGBgWRuTfqq4djUIN+bok//sQHayEYUiNysnrnehT156O8Q/COzHfPynbX1V
FoZyGZJsP/9YN6t8YKSVxZDPRz7ue4dxLmffsfZfgAeOsNUcEVGiXnlNzrRdA5iW08fK4PIQkTDO
2Db0vJCgghf0d/ecHyuWDMBiY97NVcQQfhG0qIMENODgGTTsoKwYn2uqil1TrM+YDAWdhgjXO8T8
Ke748gjpOognz1IFHOLF1gsMWoGQYZId25zBwFH6bDHMS5CRDxKcVyPH6W1NVOT/v3UthGlDFdVE
X8BwUcQnHfLXTzAQMoLaGV6Cx9CXEwSfg8BAu511h8NeEZQJykzN2Idcsb15hQvjJEdm4iulxOID
U/HpN959u/apHElTNMNz/2GFXfNg0iiTNHD1e61lB2ixCBz2Q48CmwUi3HwU2JURLNl5BQ3zMviv
5Worpua764F+MvI/mXh6Xs3brQXnLEnX9AN4pa4K9NJ7I+oLBJFSJmUwsANweKjEMEXsPsz+homA
bg16xC0w4mJ1+HTw/8Y0N9DZQ2UgaSRqMYkgW88wYxBgHuPkFuz4A4uMUuMc130DSEXehiwmDDVK
ap6W/q7Nm8YqpLARx5ab2y4WBG/3jvupaAwCuGR0EDYJjCMa+bMWheFSQr0Go503S/TinfVsYtXo
YAJKv6r8ziEgVLLVcOyaOLUc/8llRpqavaTsA1OsYMvHnPlGFXWh3eKisDgUlDkRsroJ4hkyBwJ7
5S+akLj45QJyYOw0HL4tO/63z7GkxYpGjlB6aGBO4jCtD09CK5p0fEoOX6Pe0smCWBnBoYDyg4HT
G0D5BOGuwjBNBeluoxBX+q20qvuO9JXPIwLB4mUjIMeSGDNEqpA8rDKkHCxgYZiwuZVfQ+/jGOPw
0zg8sIViqHONF/VTRlKMkF6H9O0gLXeYZ2bVWZn/NoijFymIzzEVubzlsmL1qYofGOBrOsVy2fyF
f52xxfwTul1oXHBlSiLrN3s+Xsj7Sxk/4XdPT9RX9xGRvC5VUzbOommsHjNRfl87PNkIuP00ASpo
UZ38jkLefF2IeaaCd377vjTzvIv3OKs/LhbQ4LG4xGL+89u+Bn6PVh8mYkRVtRLWrbL60x/q8m7L
eaju61lNPDRrUCclr9w3j2ByYHgn0hl8IuzePjh6Niv7RDreGVIMRitJ5zjmrzzhoTfIM4PU1kIO
shEV/uhOJnjLHLwHKlGOsevYADmP5hUjRkp5//R5sA/M/Y7uPWk7e5e7UGjZ1hIoXG+CJ+KXndyg
SB+71vmJczyCEIfobdHHUZZl71gIWL2P9KtxOB8FU64ErHJH24hNxL8t0kJp22NTDlFCz3Ecxtb6
O6lpCyk4P43B0Od19evEcDubzlge9uKNgqUVt3fhY/dbPBtVeJA9jAAnjb0zsuEaAJ7Ta3j9ZG9W
ann7qvpGofO4UOMEfQ8nwbv7PKNE57iJ+nd1Rt0IbgEG3HOVcRHCXfsQCNNlQERPkTfGR2D2rAeP
GEKHBiVHIf1u8jlGuwk9MP67y24RB6IG2GJIKGdj2U3AVQq8lZk1wfGD34DQaa+evokhvNXmrdEZ
cVhBt67WwlTbwRpIlXM4hV+r5OcG5ZW3xS4kP7TxOb1v2q6ljWprLaFJEILk3qJC1cn08TRSDTDD
LH+d6589ZU6E79QFVdzi8qBS0JFVGOCm9Yjf+VsxdhVsB2N4rikLthp9T3yLD9DcklFolxioMdc1
smaFrLlYIDpW4YBPVlWOh08m/h3vyOzipN9Bx+50+2Jq9K4n6CG50Fu7+V1VNyY5rhCLzx4PN7oy
D3I7OK/gt8p6n/HQRkJfu1q9ePZt8d7uSXNQ61slv5jNEORrpoT2n//aRUPLQT56Kf/1Ege/gQAX
RhaVxlFnkKE8AEugmnZn57oXyoUOMI69IYrSRBxGqzQk3ZDpndUVSSb40qP/BS1oK+xmsadcHdNs
uzHvVigQOF8MjodMGkLemJO3dHvgB5jR95HXrnOBC5SEfg70jhiLAfEZimN6ZXUj7b6K5msuLB3/
ECPIcIjG497iWTU/hOm+XxTkDCV8xIoJR00bB/FfZx54E2q26CTHlYYN/ykai1PY9T9xamD3+Hr6
xB75W0SqEB9U7n8aJXwziOYHfPG1gOSBY+TUcUPzhe+0doCry7hlGtiz38TQjng2sBKr8SbkTJIg
QBsG+NRZdlUDJXfBLAC6CN6NB/y/p4J4cWSREbwNihq5whq5Zx5rzZYm0SxbZchNT1jmWMove0JZ
NUOiY5zpJXGnwcLXgvM0WGG8ECvVryrT3a5nHhULYQea5Q0mFqaDJMXWM3ucyEXHeWunhIZ0M3J3
Qgpr+b/Sw8XhLbnmPJO11HDXXxS/YsgAHbajUo2ZMXTVwmkaWTczkTAJOnyk7Oc0b7TBMLWsx0Th
qWR76KXNwqATrAgAbbPX5EhuxW8mWkWVD3fMA+HgDEseOOWGZV4QWBhHAsayA42+3yvrJTh4SMfq
/uHf3lVsCGGFIIsskvVVEj9FyZNze5rb5G7cYqjxyPt2lsiR3S24k8f1nlUie7J40QpWnjBo3p4E
q6w/Crg6gM37ORmRk4AXGaQoDVoW2101mrwNPU+gS9VMBmoJgu1bYfHcnzSXQbHVAXzA0oSnZxnB
Zo2tFv6GsrCPhEbXEfGxBqPQfKfIpiZiZMI4jHT85RNl9pn0w4Tvq8UR5nxFmODSl11UvtfQcrEH
/nxa9IIysDmxWWIvlVY7b9bOVNT93iAKwfIfElwyc9j0vjKeXXBKRdOhMn+s/HdI+c/ISb0uVHHc
9W7W0qfgao4Eztz5wOG4mhDtOGphPPPYkG1ioibVfCHmJbGvWQxhoT9Ru9Nrj6p+POOf9XNpqvTb
oSfW+Ei0gg1QgssuzzwwPy49IBiN7NU+2Ym8iBNRIUWOo1KKoeq4m6Wd/T5zVHTUHFM9s+Hc6evG
5hKhn1iPB2lDoVlZS66bv0CjI038JI4ucWVqWiKGRkmfu6oSskDwyqZNd9RdccnVuQIGET6rNiBk
osHfzFFWLUuvI1sLtOKFTNpWOnkRkSuhEfpXrJa4ClP1JxsdQQxsGc7reqQm0jb0U2naHQ1uWDJu
vD56fOVB4haZHmp9zl7fFjzfzWVTSVnv3ony7vedyG8hzNY8k7CIKpugusaMxHYNSLMMx2OXJXkB
WLJl9rfP24Mbn08acMIaGhbkoY6862ck1mk2iCPkjN/HhFkhb71BkL41yKfmVaaOseZUXawVFS8j
tDn9YNzu8/52EYKGhRubCKzS70Wz2ClHqihSU0cuaObR/LyGkT9TetaP1uG1BTycx7qnxOQIywau
nirssWmcsq2+yS7dZwqK/lX9jIiJif9k9XuUZ7NFmHcH+s5uoKS9W3uCyQ2SWQNBRXZvakNrbVX4
bmXlBpwnB2nqaav7qY0s27ywviApwElcTdHES6Bziz5hzUmh5tjM4ilv8/NyAh8YMb3guKcaSHev
DWpclZZOgZ9UanXrlPlkgr/tXq+DD0CiZYbzJVZ55nIYYpL76FHmWsHO3nV7hmHFDlcYPs5oEF3h
ehjIsSzFkYZbpKb6yxUiRvSHBM0zdj5brlBLy3PPxB7SD31YmWepJZT9NEb3w85Vel4W5rtXM/xe
dM20jj3GywhlvcIGmBuag31HFfhX7tuViciJ5Xmr54gJAjPRDvghJhzIJl2cDorRtlQzwr8A3xdP
IFmiRGIa7A3azBfVfxZ6D5zcy6As85F0rXzn5MLR+nrQO4Fes1lJUeaxcKwcXAQOl+SDYqmFy8Lm
MJ4dFJZhsWHLMi2iSyR4DEk81kbePHzpRS4CnoAsbepwMaDq38t//3nk/S1ZNkXrzAM9imedn9jU
M46fQNF3B/IYHQIUUeSP521/ZS2w3skW9yGn9qacnWGuSsGGxGCfTw7PCRRcmwIG2PGCMNXiiTvs
564fpPnbPv9AgKhr/0crrqhoNHWP4NkelUOu9ZwUHiJaE7lXxA80qQlRpBBW4GMBeddjaVS0lByC
yU/96r54j518cM/HCM3xB1SI+/zPCBCh45sbpSVymk3V8L5AKRXSuFRgNa9Ih0/aOW82trwTLf7E
Iq5WoR368MLFzl7W5XUEp8mcqYEf9xXE2sq/nPFt9e9DL7650iN1Ex/t2qdcK42jvC3N3em7JeDo
YQF2yYDzaRFwubE4hDWARJlKvSsGW7538DfrLoM4ER2vRcXC/v7Ws4MrY7nIKajMz0nxg+NpQ/gV
nrdeH4ANhOjDkXh11Vx+63KNg+8lWsZQqGKmGHB6BIiV1Cg/PbJvRXB9xEhmmSL3XERzKWGeevPb
+ecVg/rUenSs6Y9xRRNA7Q43P/lmw+1oldNPDt6vIVBOzThbzvdQh5ziE2+vsxKk6AykjeAxUEIJ
TySferSz+80uCZCS43qHQEV0GnnYvh6PsP31edCW4oC1sMX6gDHeTntwNmzOsxDtTXrbqAddI47n
XFPri84H9gG7CvicM48YqHxV1BymCwCzpEbpTatswIO6ZeoXR7Rho/FBcHtsATZGnS7kEnhRpXZK
uh4OVo/VLVPx9N76yBUKEu8eyTmoQ4K6R3wvnKrO7e2/TIca3kiqu8v1Q6lezaafSu9lMFnTiezb
dE1UeaNL0CtbUA/4qo6Lq8vUx7hOOttYR9ms0HoHJCX5VD8/d64P8VZgLWTk0e+lDeCZ/CSEH3He
6fZx5K2wNEWAtYUkFel3kZQimF3aqQ1Lkk1bVuC0UEqWrux8MH+S/7GaFTV2dVZ68x/ARiYQvsuU
kTdjvckra3DR22H0jMHLQZvD9j7swroulI738uCGrb7C5X+RG5+k4DJJ5i+pQCspdkaQeq0g5AEq
vFhNWZ3CL6dATkW8PvSGkptkI7FW7sJdgAbpTuv+4aHC30p3YEk82V8dzoEbEvJ+liZaw6WdkDy/
aNMEyfsNHoq+c4+jgWwvHmd7BlNkKOIkIH1T12/A4H2kVYbp1khKbCcVPnY4DF2RZv2Ea1UkCEqm
iUrIlsdwHcf6cIn5CIiXpTMBdwFdyP13C8HpfkSwB6LwvJbsEuxjhQvVfVZURzn397U3Tymvl4Ss
VmDDOBDVTKaStaRKfufZNodZ/5toc3B1n49Z1TDktUaIw3LELUoMbkxHRY48ixcgqT0Pyh+WeQdf
eOP/6erPSoDM5xMspBemlZt2A0+B+xHFE/8LbvQUJW/fhPRmofBDHMUbusAk920o+ZhtCoblZJql
22eAuKW7jdAt4S/SheDfD4f3wPWgpoO0/JNYREK1qH9pl/LzKI7mqUsKcFKgemQK7wpZYEHcPb3p
uHWEeGEDbfwVehO8oqJihbsLm2c8UV8DQgitXtjW8RttdB18K7dsd66aDRUwnW3vB3T4NFnzv88j
l/SErjIjAp94jdJKfg7ZqGvjUwfIbmAljjsw8PWEMx/oAw3chX/SiIibw7EJFHn9SUEqUiFjNyfj
T8KprL9Tw8yNQqpkRws8ysH0+/DQi8kFND0x22BBum3i43GYUS6HbKnfURBIQRn6fJThRscfmXOn
gnQlFAejoGHPV0Qf3emMUGf9b17csMY8XRYS0BXKr9kvvbCM/fIWC29UwUNEDOgxIcvCBzFjEmd5
AjFu+jDa3hJaHyGhJVNw/6lvNQL882oEtqmeJdaUNg9dmuqBtpUntDOvl0p5J84V2p170Vpd2DF9
Via+oJfv+3Su3rg8USCK+YFj1axgANN0dh2AVtbfE/J6y5eoo/o8hErsu9rzawoLOiGW3AGrVxaB
apavzo4YmLR3HiBGykunC1cuZCmVsiPYAtr2UdT9h2HD4nQjGglEtkgwyp2yFiSvUEEIQn7UT/h2
PxxsUP4pzDjPqPdR4RAlXXur15QHmMuQYv3DHKKGBo0F+KMvMyqod3jB+8403bNQLzTbkatD+MMp
+ZJurEZH93eRbAdPI9QO9FjeY4v6m5IJhkEP3D8BgUy5PJ/X3d2ZpzFxW3i4z6/R92Wesa0qWhHB
hHdnKHIwXQb4QWOjsB8aP75oeIMfnYsC0yDiFcw//0c9X1wsSC1j0gxrNF/aPhxASZZ2SDFD2Ctp
EjPyMefZyWTyIg8MLXCgTvXJxADBYpfQCIlmOTQ5E+HtqM/OxnlmNjsemBlujlahK/S3RqKrEV2H
YEXGSdrExfKuxqfG5e4KRNBj/X1O60kkz0fEQVL7paVcXzKi9tYZ067GilN4JL0zmn/GL1KbDVo9
12Q5rFxc0hmMO4Mlr1qJQdFhuo8Jo66W771BU0/TTkY283bNTZmL0fqAUuCCtKzWiFv4RfBgz26G
Bdc3NLCic3WyFwosi5XZzgAefAGkkTkL0RdJ2USZKEbZky/xOenYiripmAaPlwr7yGG30T1L/XMH
5Cm3RACJWphhz+HZUoi1Q/g8fYJ6W9Cn8+9vAYhiFgZKaKZd7bB/mIgoaa7YseH1zx/gwApIFD+X
hVNPKLTYL6V2J/nh2hDE5QE0G0XckkoMSImY3WTJFW1N7jHIgRBjr/wjepbaAd6D/9t5kr3Zbcj2
OYkkDtc9L61AnSkNrEO+tlTIflKk5Hw/s44Jt5TgTdOhG7G6uIk50P0XvwFW4E0WobDS68qVbX0+
9NWj9cCipNP8gwZLYVGlQXkOB1Oo4avC/5cMJM0zkLyY1m/vCvqhPH0IWXrnzL80zw0R7hAw1q/9
1aSBzHyafV5aA9jRY9nuDb6Tlqr1SJASGV3OR7gVOgDIYY26zowo4z0+1EK+mAferCPHgoK1BoDe
XrwmNIdZOTH/VJfwqSdpleKHDb4RGjBY1IKfzGNf3B76aTFESORrkpfvsVWExIORSfpBFwyVC2Q0
em0ZHvVGHjLODJkViEHfoXER52NhFgnXpU5+4xEYc8VgkylK1J5eENot0X9Dcsrv8TIVgy9OlKqL
LyO+8BVnDTE+LXXZEifMwm/DzV1QtIjOfE2ejTB58ypLcPuOvXe2ZrgIwbWFuYeR9v2ebPCam3/k
fvzKsa+nzsCY6mZdklkm1KDUENpWH9lW8yXRW1WaKnGgJqib5dHMlbh2WQ9+o69VknF0v3VmbkN0
Tq/5fVt+jVSyKA/Hvi2CXaesCS6Z/OC9bdbnCpHy0BApAgE2NoUCuytXR7u6ke7ZWvgAs5gTiYqf
TSkcB6lf56hsfPdMNjvksnRTUF05k4vY8qoimK4XITySUcNh/6Avrdspnt87zUcE6suCcIR0Kr8l
Z67yicfMETL9VB7X0l+ARM+gO2xO5zrefu5y2MR8MWgtv4bkdsF/QXhLbmi2+0t5qvOidzKK7Jj8
dz+qtkwproY2onS2b5J2uDf/LPpyJlA2XI4BZp6Wnyp8fLhpziXBnmLwmTiVBHGllWShATKuVvFW
BKWE28y96BV7jIFMkK73HqPpjqjGrWznS0lq8nrx4FHBR8KfN6yR5/xp+7PHyMoGTkF9T8OhTWnw
/qjjaJk/7xRUgJKn7SaPpSkzrx62eYjUYtlPB+N2HYh2shlvLyjgoQ4RaISvjhkmSE6okL8NpK7s
hEAbpiWeVYDfEz3Xk8W9KhxX7REJSewxeahsKJAcvqVMydEiBzCD7xHb0/jbn96vG9TTkKaQzMyX
3WhtEz4hXozPvAD6ElXTmkjJ8M85gwzojL6gm6h7pWmLvqN10neq/qMHacNharPFmlPAhO00ulGH
r/fHgHSg+4gXMzf4TM4ckNVal+MxrqALeXv7N9EH8v1X1Y9FQi/XHpNNkNpApLyTgQbAUubcERnm
cmPA/mOvEbmh2bI+IFcxz/Pk8+8WeBpxg6nUdoYVZVkZImFcczEh9KkULz1zS4E64TwffO7IqL1e
BdgKSBE2P7ok/xASZ9PBnGHME2vmrwQTSqISgq0j4swMekuK5fjkLWq+cCLVSs1E661GxmB0xQUE
ylpo6EpZibKMH8uNd24OrHNjqZHyj9GCTIAECxwxeQ1fu7yWT2VV3ePCcQG+fsBKg8yPl3BpewAk
Bki/Ygp/lJMKvo6ddU8rpH/H9zroW1tZ7JqpLiRIOITQyCo7SqphwfOeDMycMws3e1Dak9rbIrh4
4Yx7EXsPXF2FYIQtmdJpZvLhEHeEcnbNzmsb+gwSrukJy+Vn+SeIUOUHCoj4tYxKwTFz2JYKyuyJ
sUmnIOIFL2Lrzlv9W9ne+T6UkQkM1UTNk8TDCVUsGMwebFoujd4u3/6Ashn13WndY6tp2myX3/sh
3gF/hk/hgx0zRAyHBsm0GJfrThL+P275U93Z/L06kklS5OxWpEsD6MwbsQFOUWvnf22NSzMwmSBv
psl/AZq4JrGtrI+OyZKUNh9T39/OeoeVPOHfaX8ca1UtdkRm3VdKj3hNZ8UkG3VbkX6CB409bMOj
8wxuf0m+ySQQ5cxnuWykU3QqYZ6qzK1FQT3DQWmnQptcck4QviszgU1lmsDmWcmubRBX64nkmW8G
ZLmf289grYuwhpIWDMOKZh+FYoTTujES8mXrtkcqKHtPz/X8PFad5QbkIoLtLI2gp53RwoZIOek5
S+REMnZac7B3lAc9tDV4WplpsSiFwlSRz72g3gOf2TJoCuFeshXWwnBtiwWYxeJKcJNlxrq+1zgK
hUS1SWWXforW/QY7LIqNUnBzBar2tRRmBMhSyAVfNFw8hD8KO5REMDJYHX7XUnPkTuA+ICBIOUcS
NVdgRMCsD7vtCs+0zGHFg32KsvJo6pXN+xEIjrBtFDOwjo1nl/CrGaw2iiom22CXjd3yTOXVQDrJ
ydbFCe/UJFQSfvi1oOl0tR5xm1Bs6rDessCaqGeDrl6GnoAYuAclJr3LD6rfpSH+OmnUGFGg8fJl
R6xbOooQWeQ97jEuPlTZPhLpWOQvIAcTovFUbuZbgLAfjZWCtWxFRAk2PYnsi/oAdw8AMTO3wuRd
Z5Gif7J5eIn86CkWJdroAmHuakDzi9aXUPzre1EIfilLzcfBXNxFeCpZewhZvXzqM/GEIDRSmXK1
rfrvr4CY88su1fih4W/biPf5zOyV51kIVDA/0o29hCjH3YOefma74jIMnOVDW54pqP0EincTg6pL
Xy66UdGXH9J+z8hUb4EPyWZ0Q2rDob2vit34GWRDsjDpccQsR9lX0WrCllfILiFhNAJ7LKu0A4Kh
do22VL7hPnq6UdQgIMZS0dO7jMfAUFxWGYnMuY2tDjtDqOqYkyh8IwoaDj1lggwj3mOdgZ6mrkbG
6LAJRpY+g6I/jdw449Z3IFXU4uuVC1tA19/c/m8mRPPtZ1bV9a2IR9ae7h4n7mQ4zokvCqAomn6j
rd67QUA3vVfbVlCz3psMc4YkbGPBIvr9bS5NZTaGGUPV88F/1zBlwQpnc/qnLedG4t2a1ifYcXe7
Q0rBvWxkWkgU9pDD3dV2J6NCMxw+rY3BamLY2sogGEwxAuHAHZhTOelku6IhTSGyqMEjQzsEkk1i
jdKWlw+hoFAYgoY64Tl9485GcDwELIActNh8+tzALshpxejsQ/IRhDz1g4KlIptiyb7xvEQb0m4s
lzRvrnYQ/FRdQiXB9L+0AKbREu7JmcF5Af0V91NKcOWTCAM7CTfvnkHs0Zhajw1UQmTiPn6Oyzdy
hYr0XNg3LdJs1DkO3/gQdSpWKVwCETbYsqfpzdoce/3PImG9ZxryA20k6hRLMA9ZVuahaXcDBq5z
OMoOjyqOZl3ssH+pzYf0YASFIxI5EesN5hlY/BHbls68GGYvgPdPj/m6yw6a/jIp6GgdTl+G0Swb
zEk/aoIl3aXwG5GjTbkWYrKQ8HKmM8dL8o+Ljh7MRgd9W3fg4KKBVuu54PFVBqz7Nt9ZSD2ob42w
812Ngx9pE7AdGlaWhhudMBFybSUyWrOQ3L4RMDPqn2ZwWaeLT47IMFVAqXk/XM+JpTNqPFMb925i
VR8ORdXLP3W2jtT+mMAY65qriRokk0iw4JARowTvSFRVl70tsSvIZtGcz9Q3jX3ECiH42zI/JPO9
UeT+pdm12ZPFwcdhqgK0x2bf3g80w64yBpYq2WxeLnR4lGXeaqFQI6QZ0kUKhgn13PWGhA1g9iFa
jksb2IdKLjUCV1/146e4LhcPicJpBJC0Jys2yA7tO/xQMeoInNICW2xO9YWmtdTbdja/f2AXww2e
vX8hrhqXFrnTfDmrVNR+GMqaLYgIupeEUIxt1srw6GrsjTpjCESYbCE9WULYk3+rfMrWzkTkh5sq
wWkSe+4ysLbth/lyAzwCAkMaiOz6p6GmdhUHemR2iEeSJaTJBCjcjX40tdnO63E+AeDayxz2Nv7Q
8sVM2FRkptFpGffO7mOOwrCylg4pi6afq0rMkd/vc0jwWRosZs1DGLNys0GBollt928szZ4PBVh0
k2g2Lrsc/Ok7ZmFdCrubv8r9oTu5+2nfFhCOcM68hE0ICAvgggO5f+b06YK//Sx0/SEwrUcpZUan
YIeCEshMdwKiZ8A9Zh6vOLr/D3tLX8w+XILK7BLBvlsrTkbZpz1jOyNW9IZW0Wpy2EY7ALYWTLSI
oXaWd9DTIwwD2Qio4IX9qhZeqzdoE8beKTgVyQUwC4bJYlRB5r155Z8nDQx0V1dCHDQNvp0rMMYQ
zb/TLO9C4SFbRiHjxBDdUpJe9JLeWVw7a4rL44YGaV0kk2QP1dyNmSsyQWh9BcBOK6AT0JIe33L6
g1Euyg6HhSZx1eSBednwmCfxuLGuHqWf11NJcO96Klae6FixKnK9+Qt6tuQJNsquC0fHoYJ4iU/A
0qxXtYAW9YfGy7F7X3LbRozGsN+lREtKImr09LTuSAWQ6UuVwUihfZlHpiZqsirlrHr/6JbGRtw2
4WsD7roEmyIxOe5PgWsYj8R85dGreKMg2dQN6quFk4t/bOCphC4+bzM1wI2iRUZ4H/veubAgNf7Z
VZwHMmzYNWxKW80OzvNl24L0eCC2yICy7vmCsKOhBKZ0mgH3sCLOnIzaNfIJ/gChmBo3zefh2dm1
JjUdLuF5j/QJrG/gGQIQY+hD6tnuyTkPirOgdACcJy3BNfoNAeGO7Yriw3CkYC2XI5n9OOp3czfl
aHbwt7UIU/NhA7Hlz6QnHwrCsK+2iVOSOoivQJjl/0NlugS2V7hvMyYNhm12B4fPtqONGleF89Q5
3oLoM7MXPn9glF2b1sqVi8mktyTqkxQZh3eixTrC4tsCkHT1i78I9B20ikjGh+yGpL4WwYIsw09m
gOVuNAWfCxG7vNBBoxVD/5uz6odPp8d3Azdy4KBJ8fwTHQ1AfPPn2ODF7+fcvU3hId1cb4F57Loo
paw5u6y3sryD7ScVb2uUe+wj4S+dGQTFGQQwkVvtT2SiKFriisXEFV5TSzhNlYgrmkFe0YhdfSPb
HGsgZNM3eKWmpmgxjhh+Iaeat8p5tOgveoYFP488DYjrIdflmujJdsiwOKicoQZeuqIqCBFiLeDa
B15y1Wc0nZNC4xCBjfwrKiNBT2K5BTYp5/AYuh8HtxE9fi+U+NbmZo9VCiWNld5i1DXeUU75NuGr
sCAqrmVepVW7C4426/aH6jAsCDtQgzq9Og+pjTPmNHu3hBL0zZjLk+gIgnjjP7ATvJqgcrp01XTv
Bobi9V/6OdKm5MqJ87E6kCHBtik3E3j7gvLu9iqrS71BKirhAlIMjytrCwexXHi7XAOnWNRzacoF
pF0QeaVS/l+O4pnJGAoDpFY6opvk/jB2Emp7LO3lbA8NT8vLCJlkHyKvrNo5Rug6d145e4xZVhQn
gr6ajmujNt5J1EbCx4v9Wn2EvFBpqDjx3r9cr51Zwi6Wnc/NAzzmOB1JZCIG1jSdc9MxPVDd2B1/
it4ecWZ8z6kNePabDdfBq/A4w+SA5/WHH4sMPQ1BpMGwvEfd/CZkh4XBaOunEUOEr0rV4xuIigrA
g8CcWlMqVKVGuz3bZNCW5vr1Hr2b8VwYz8Yigb6rr87ovrMPzPdTBpYoAeajASkEJH67zzPAn1RU
zyLFE4wh7nvdz59ukgUzHw3NAljChRL8h8L8Sh4kPM/ozm7rGJ0Iw/3a+aPO2eYafB7no0ViA6gc
dvm8O/be1mYGSVPkjBbCMNZToht726OiKjnpD6izpf7NBG+U+HBXPUHEfxdI0bFk512a0XemUfqH
hVz8qcn0LfD51p26QuhGnwQzdzE1cMYyNiJKr8/0h3to9lnPiHxBitY8YZkOnja/HEPw9GnjullD
LBU44jg3T7uzs7ahgBl/nQhYiK/Xl4UG8mkR9JuGh8H+DZRwf858nCoyGKBsWL18lL/A4cTve5jS
yrGwGNTxEOMuk/aDtilhcudItRSx8ioI2C/YJJ5pE57sQAPEaJ9mVfS+fTzExKLn9MCV+BT9cRuE
qdrB2t4rs1zB5mHMMdW+R+vhOX2j27ZqPyWVXDOH7Xl1dYOSIU1IjZwm0WJpoaOARKwFypJCeo1Z
rzGtjNhTl1GNZow5iXKAscneMCFuiVbpWLuVUIKMr3o3gYlDCMWKLzrCsFLJqzHSz/kvmwV9pgVj
/UnZhJ5NbvpdmaUx4anU7bP8Plc2b9Gkgih7ZgBjVItX/4/Y+KS0QqxGx4vZiq3mbwKrt6E/yQvT
slfaA9QgCCpLw2BA6OJqEgnc4dy0JK0GH1iSfcSn5jDRIvwViiBCpeyZJtWzQjE5RrkqhuxidTli
M9ehZNqO1tY3e5PQRhCNrK5XXYsN6OCJVDLFxRplPCdtpGmwO4ABSVI/WToos+gOE/oYVS8Cr31K
KK8emJKeupgMiRpKy5ToXUlINKA0OFfF9i9FdKdWKungetSXU6dhefyhflp/oWeVZtmsdNgmJLQC
FhBsdv7RMyP4VdMKBna4MXAfI776KRAjuKT0NUDEJl3BO7qoxt5oETJ+E3vd9L7Zl6NdZfhdfo6g
LGQ9odnuluJnJ0/MwaoNkoVzwUmn0zgm4Pv7+kuUEXnt8+K9+Bb7Yn3P2QJfv5OHUrCKFxfUuPWo
+vnU2nRhsLa/afmtXZ35/fmk2S92ZCIwzuv4K2cBdqQn+sxCPj/dDlhICeSwObinKAlyUikkpcQz
00/5xZD1aS8nkMwhKpxa9RCQHqrdER74pEcsvbo1tABIqLDe9R/OTVd6z+wcmsvBniqfhWlEaDt1
ZzHHks5DnRekQwjXGUdVLkK9GF8GxEuqrZGSz95Jz7hc7RMco2XfHSSi/diYaf8hnafymeB+Fsuy
T+YEC9Kw37msQ7cSvb9mEngJzZLSUTdtkPRFYD7yp3NCweHTerNKbW2dAbNV2grfcp+VvCDmUDV6
thUjvUvFkZimkAezuOqQKqTbdzj2C5+7P5sbz+LhouLLiKuHVGdYpIM6PFRNa0QqngSoP0yG9wzr
zSVWaInypP3IV/fmWSUb5Y/Lq3k7kqZBSMybO0oyloF1DOd+KfPpmy00u3sbYTD2oaSvtBvmGUnX
FUiUwWfFoOSwuuka42gmHb6UJT7jAehmlloEdKcAY0XnVPo3Npr63hfXHMibe006rJXSGDaElZg6
dt0BwfBsZUlb6Bqi7GuXEPxXgd1YBdIBEoUdSZ1/RAAsM+zsP8r4OmvVsNTlWLYm+YVanIzC6LoT
VZ0aIMFTNYSig0F/qho5xg/J2dNKlPOlFtQGugx2sUt6j+Q52Vm/txEC9pR6KvQFJ6Mlk1YWyiRW
iJtxHE/eFO9MwpSsX9DZvMww2lWoimd60YcB4kdxxFNtzyfqJq12Latd8RKnYA+d1z7Piq8TPEEb
r2+fduzAc+5QEg2M19/HRXJYLBkPDeiZKLLrtNEtDI15Z1KuLxmnOtHNpqtKPWhwN1OheEGa6dB6
r5LMeVvgDxQi0KDWKjAOtrVhzilD3ciq2FZPVjZ69n6ItmaVt1h9f44TnUd9/+3xRGNN7/rDHAUZ
Gi6s6EpeuDxMoip/mz+dScpSACrD/nCraFFQUn9idrFFXiNPKcDdec1eBoiaICsLb07MK8KMifur
PxLKYDUGT8sT+ER6wWhBiQli0Q+Xqvk0Oq5Y0u1lfQZrMTrPvwVmil3uyFqviXP1QFabpKcgA05g
w7Q1cOJEVLxEMOu7eB3cdAbUiaOIXQpBJyVHcdTz+/kbecG2NP6xASMpJyxOCb0IFBpL9/vZBAA2
JB5bt5pJ6V6aQDfZQcF3oXi8O2O8jLPWrJ3Tl1+vTBRSVTd74+UVOAspoD30BnNirsYk3nhfZgR/
4F67PlTxgcUtiXM3tNXx+F28YvKRLVrySnOfymqLJ3stSgv44bhU04zhAr6QtrZhBNKYWCBtwsIf
5vn7Yfci+GIf8Xlwz2UicMB0tq4fyn9E70X6B/I6o3tGGbhcnBmzlBT9l+XANWGJf0hjkZJH/5Aj
kkepOTFKYqitcEDt/l7dVcvyZDPH/Dk/f6SvjWv2x+RfEcpVO6vZxG8mOLh/Ad9kstgXW404KsV7
lGWMra6bxvBI8CGV04rKYfBnHnlw0XyV8DrDErmwJWuSXQL4z1BiT8nmGT2hNNK9hG973RDFGh90
H6+cVhaRTgKJbhvsKTPXqlFhGfbjuTqMM1ScTsBNFO5BvRR+eACMOeWIaXnF+x+tva58PgugqdOr
kMB/jx8i1ItGl3xPXpjpBN+vo2qI87B8PaD7I0UVmeN2BubYd9rKaEGiF5yNF9b2QN9pMHcHuLsL
KN/pG+jKve5o5F5W5N12Tpf6LxkvSF0qesZ9SYEC+aSWzuBOFzq/LLTXcVGuDJHg3pm8O/gpDk9x
dvGng5rjd1yLH0BjtsYpRsG4hioS5FsbesK4Cu6ef+8X/cqIjcm+E7zAa01gyMeyLvtbWghRGj5j
a86xJS9j4dJRLHPe2cB2RZ2XFIoWertn2byFXfLGfuItJBTjAiKH+EKG1HWsCwKZbWN64U9CCfYL
r6/HgEUWXkInI+RVGHfADbwufd7Hupi+DS9ExRKXwgbN8vUEFpgg0EP6L68QQ24k7MY8nBSQZb11
mQYhjrOZ+q5zNdbsNdTuwFoMuxiEPWmNh7CLQjyInxmLYAK8cz7YTh2f355Knrf6AzhYvphtHr3a
JdmEWRjq6PhUY+gMf6borNcJu5ojuw07ewU6Ad8GjZlIGa8G7oMybAUeUjw2FzP6vdKMSpJwv5aM
qBxRrhHspYlSuqTk/az64bTDrTHCjVXW9JxnPh26Y0GhdPO1YzerElyO162x0Jru0DlsI0LxZHVu
SWc3VKOmZMzqTIIfpwfy5kStXZuKS444nQv3iHlo/mE7+KmvCDKET2Uk3wfLfZs6AqKTqdA6UwI5
ebYe6lK+HllLZWY4up7uvxiNFbx/IBYGzAx30aLHf0WltYJxpkwLm7o80gOV2+N006w0BaXsZjUz
+N0V35trzCZx7LdncPAD4Czh5ru74Nhp0OX849SQYxXWpdfCvfHE9M/ZxodWEVFcO6WeO4xdMQkr
l0m7Bw0vkCQn4UAozUwFMls8/pWKa2seZJsjV3Fj9KKMsMdfNy7x/8eCzdE7Kw+DoAc7uhzgmKaY
dLJI4y1ajBPCbQvJRpOZRGSBdX2nM3NifiAWn91bkJBEN938mOPsFbuz7qysOoytZ6x2AbLseuhH
0I5OSlqYHgJEMwF9oL/DEWDdZ5HhBzgdAcxhSlZERM135kyWLtG2ASeeFZvpeh0Mam8vntiSMIoX
0GeV6cOGIg4nfDQwHhZftn6bDpGhIu6YcK60yI0O9F+CdlY8QHywEUzabhsTL7cZWtL+UFz9RPKk
xxKvKYKRZI4KbjLIlaTirpSMPGhzZpMkO2+Fu7MCkWlMWBQP9n51mGgBuGVFWUl3Re6Lv5bqMlUN
mFDYdvS/w/33wvsV2Sa7z7mWf5Gxukm/P6M0iupu5UYsFSlZOq6YuwMPsTvv31FDXwENTWXdYtiX
DG6ei8D3/OCItpvMaomaTysUJlMSMEqOzaXumoNGQHNdfLzSrDWjWQx/AhZe/nBCpfyW2TOQTkGu
sY9ekSBf3AWbDoNU8JcGVYtXS+0p4WccsBr6nmBPUWbiYBY/1hHrdGQ1vPXKu7gzOY5zOD1ZSpOG
rT5tqPU02eVcsuCHzTaGewBex1NZ93zV/zB+VUxKGDoA3lzOGAw4j5abDD/E5BLGqDruBQ72Hyqg
vWTn3iBWuf/BgFE0Go+47ybrUQzht0DvOKqQURz1ZgmTBK5P9r3LGcubc2BLTzOhh9/iZTwMak45
C2+ZEK+tUxU922tqh5v7DEoolbM6slZZBEKwf2QTlOykYwoV7QM+xlDUa3AMX4bSt+RHST6kqijE
VLZlYziQdM4yqbHAUU14qQUL8MyHi5ELmO/p4+qwpiJPO+9UpkG+qkjXy+iScJrTdAGv4qGuQ238
qCKCqyh4Lp7xKkUiJ6+Hnj3/5jrAGnjL2h2nEsyetPDKtUn2EKG53hLX6g7YMwinKyGpyO0Mibay
a8ww16mO6Hco8twHTuTiprWwNdub+AqTcOsWGVtNtQ6oT09D/q3hKE+jeMB0zNaLq5BiM3xuAEGF
bDOxJU0p5TazyVSHeeNuKoyS2aX9pQmztkAYVjUiDE6WMLVoUeeSW7uvVdaqffM22Fu6wD2ARiVG
6RJrddetsid+7QqCGd2eTYwW3U6DTR4hrT9vW61zqd1RyCTFVt3Q0/ZGQlHKlH0EcVcEO0NTZl1S
0Kwh085wZkJNv6OSkb6yizJi4BDUB48+1y08X6eOIaUyDYdHPLrPH51deiccLoRvZ5Ts2IZatcq7
Te2ZQRhe+2Lf3hrzCxRroBWZDiJRsYecAj4vI1qw24voSnXmuwODLrmYe053VcscnjB6rlsPkXW2
U9U2CLBXu718WtRDz4tvVodUjYBDNaMOqCbuw4pumZ1O0llb/xlnUGocE2mHtPmVUp2O0KBS4AEZ
16qQ074c8jYaagHCyWwzjrGW2BA7a0zHO7x9PNWmamME7rLStqOueIDZ15M5XMApWae2cJa2jGUq
evu7w6wRPuBzjr0CrNlZH3fFZKeh5iFG7t538QdQ26yhVUZEtgWNp5/TjToO0aH6U7J0mBUfwltG
gUAlstcx+l85CXc/Mq+9nOOCrT3Y4t/B6mjuYBY/q4II9gfG+cTyezmQucXFqfkfY3aFICqmAKB2
2k1n12h0KzTde+OrSIm0fq17Sver4ESqndBB7UK6Nje9ylu1S106LHor3vmsQ4YX9w7MN5QbpkHw
M2NZWsBrubA/DR0IUjeO+KJjEJKOUVq1N2c0iLjcYdTW6J66WXDk21Ind5Okvg1khilHT48xUyo6
7EIHa+p3X/oVlG9cA6X+oZrHmxJj4Q+bbENMDU2WF1ta8qFT4UrydjsZI7iwECIVa5553Yvrp/oa
4rquETCAI4sm54MNhhbnPX/ziC6jcKs4JQ//+Gwfg2YguZl2hBQfokRAl6PugV9wcryKRWRWpgcM
/xqNYGr9SbMmawiiguEdVdEdqHKMIT2fOEi4K7XTICMps3LXsTequptNazwLM5GOAgt3Y6iZcmT/
8AnROHSwUbUzs6tRX/e1/yG5DE2a7wghm1Wb3IjD6JW+d+IJPrZtWHxOPgGMp6NJ8FhoSsLJt9Ce
As7Xfa4HNHx1Uxx5m2modKZCy3PRj9i1NyBiCp0S5j7rtPUdmc2p4UxtmdH48KQiTH4wIdOsZnkz
RW/XqWsMpt7wnrW4nD2rJFQdQuUK+chcnst77qhJxlRyAnitXWRqbST5eO/PipKafsdWtXVANb0A
XvJyF82EFw2BUsajvzcOph3gOfw2J+SyuyoHHcDqCp+teueoFO6qmY6pcFTkYSbQWBENfasxHKSf
+jTPiwU9cE88IBn9vcMjj4R9ySRbuo36NL3L4iH4UI9uKHei9LjxCTEXLpvmy76xGygwDRSHjXNg
z4nkx+Dfl5mXSIOJbybXXVX0eIWKv5HzbDf99k/hRU92vOMUFBUxPdkRhzB1/5aZUMdhuKKztwyB
StFw677ZayTLrZibqnDW4+LnkGvwOq1cVd4q4U6jorDn8HNR32s1GFMzdMcZX3/UH/jdTAfDYXwd
TpreoRxkU5ePX214nWw9i/twB7mHWclZE7DaJBucZJ66EM6CHCABCkWDFBzZNc8PvCB5QQG5Gnjq
1A/NBGYA+2O5bBeG2Jj6NA74jRvT8YEhBzv4ltCHReX3cn2A95fHaywbSrWZgnxDQsUCNnM8WL6I
HBKosrc86RSgfSGIRt8tTWodvJ3kBwWcNduLzccQPXotycDMGCv5UtzY6pJbc6LjM7MV8rCGo9L3
LbWyUD30ZiMBVfJ5eTFvNO/jwgh7lSGdOJpTUASvlXipouh6o26+y/z9G0lu62tZEpkCjlyQlE0q
MUIsgXvlLdPucL8aah8Or/7W+PCA01prZcuzvmp6zjawT/1+1HUD6Yv32ADMBAz5ppGZDaWOVFkY
Nh8NsFAwMPFiseTg//xqc3qwuW8WyFSW6I0RuaQMdTSZrTNkZKBV0RF6Vm9yqfDm4/cdOJShguSb
oUU6V0SOvpoBdrzod+x+er1Deg4TDbmtZjkneUGrTB9JlrAhJF5U+gmJPsO+VOCZ3EmVX3UjkmqD
DRReScgT3kvT3nBUhGDZ+katjZmCkvrLPi5TS6MuiyGMsbrcaxiDXxpWTKZp2yOkLcmc+h0L1MsL
xPivYlP2euisXkxRW981luKnDuiA97iTnmBR4kk0/oO9oKUxFn2sYUnCvcf9U75gtaR6ZVRYHXCw
4iq8ZzMOHf963bZ+VnCAdnGuBHsS6aw2J85UQ3zVtpGkzVKssv5fd2H9ZFSV0bL9okNfaTHxwyFM
giAqL3Atsz4OQ3ZUEXWwpdJG1KQZ9e0CbdcIKG9oD1UULEFT7Vko2nuPaScoF++RR1gaTsfGwDAP
EsRe68+DU1OtLaehd5AJr/jH81YtM2ids1efIsXIiB0nEP8uHBZfMurRCZRxGg46T8gzD0rXNWgl
vQ/YhmBvY6mkZPhivqWwd2m9eEUZVwJU99nLSwVfD/LhxhVCpvfOiNSWGioDZoyT7e3e3VPMcHXv
XkxbQm9VHFHOjEt6Q858ZYMQ16u3dLx4q6kulauUMrt6cNDJZIfsyYlhA3BnQ6Im1tOPn21OZ3h2
/5N+/3CpbLb8dtbjQ/v18cePQNotYeHIJ58NBE0ui56UMy+7SOO9RIVXguFA6fAFhZkGToV8s7yr
ohjMdnEvRfmTCyouJspXf0VXm3r28ERkvfsWcjA1H8wdcQ+ywAEV7kwhOhfSxhxjigoKKcUkOToj
88P/+WQoRs8WIt8MDEwg/mU2gqjbaxYQw7S2AofTNNax5o8R6cTu5i6U2cnRuX9FReTEdnOLoDNv
euOYQI/XRoI6gndP1DI2i9OJeeKTtQUR1LjbPD4Kwet0hUFWtn1cfnyWLPWVrQLhnzSfUa/JSsof
ZlG+nHsVBpyk9KbaRKpjrdhib/scBqxuGZmHbvBWtdf4u1FjKokOxjtVW2PB3XqjVQ0s8Z6mW2jL
voD149bLifw2uKTiKxUY0Uaibg5ztymLO1Lpuae2Y4JAHZp4Xi//m5CbQGUaibYX83zT+yFzVwD+
e9ftfQCs9v1BZ5YM7XpWQqEekXrKwAcGe01AFGajnmVv1B+tgVCv0GBGknRSvdSNgWFLpOZyrPTk
V6fAT2isDBoso/YK/gRGC/WnUkuJgy5pgEaSl2VemogeCLq0GoKg520/aVYSh7ZWPMmnjdLyq5J8
dC1SO9ng0telDv5LfKna1gMkvXhkYQ1gppjXAYgs6JVEWlEe5r+pEgYIaL9KewpmefEVKWw8GlEN
jgSLN5T/SoetohO98UFuzSx/sN/3wTF+We+U44U89j/hzMqN8lhW18ffOWxR5t1Rue5kCzrVXyJ9
9+pgd0EGGr7TeVZ3Kh5B69c5e1cYSvdKGUmZ64VdxSpF5+ucEijDKa53oJj9hFH0+uN+QP8IRRLR
Wg+KBoQWXL8Rgd69Kp9a7jgnKBhSkH9JoyIU6J1TgDpmDwcC1z6LaHWcaN76AAZGO+/SkOH76OCz
JTS9bV4D7BmYslI8Oic99invvStbv3zVJNqIK0+oYe11amLCD4tEbK6iAUIrOlhr0pE9j1abgVpl
dorhyTDQ3YkF902DZtiRQW4z4VNCRgvixeYj3RODLT5Z0rC6wILOUfWSWdjTuqnHXJNkhret+vsA
xCSjsvwdcWyWJl7t+mAHOs8K/GK7LXV6Ug4Y5PsuB/NHuSz09hMHZvaEkHizQHP89cg8EFTWfcef
sSsNJ7GhmU0F5LG/QSJBKfRf08TShd6DyRgE0rMxRgM/7cBICtq3KWTzypDCtnLsVADM3mgqwrW7
Rzp97zWcuJBtvoPkLkJnPFzahNiafaig9PUje4zUACn9sYMCkIqxGvtS7o/X6eze15o5QAsOGpv2
2K7X4QV8ezALui/HnI9kN7afO59/MKldUxQaN62t5idFmNU5q71ttAoeKxEe00lyj0Rkoma+eMHz
oPS7uIzb37pnbMPnZQcu1SVlV6YWqhLY/L3uYW1lhwpzYSeIMGoxybcXtduelcWEUzNrp1sMkkZd
aS7luoKjgCQaO8PdG+GjG/lwf4WaHUJYtSIl8BSM0FpgV8jR17/zpO/BKSTLXJK305uyiEjDoFRB
jqNiWWSKDxEZpj7v1xnyBYE4+HJsh/3NPo5lejHzEBMHIWyCuqFHYi2l5gBV0OBCCBptjczVWOKN
Witr63fkZ7+txM833pJvPiYxzDX0GtL2UgYO4WbplSug+8Rl+tOcDO9lSh31pXAw1UvjKI+BWsA2
8kO0l401ISf+eSWHH5T3ZHj36KKDkEyzCXfetSqwmkXrkTQh+sNGuJRv6iPyZw+HUId3cEpBjHd9
Gh+QOYtF5ETnjI+sBpJ/gU9mMITBaA8BjcPd2KQS5fjt19AwjQf00MAC5ApUW+aQyUonZEQqzS7T
O436pQPXzxepDkt+bSA8D9qOJMdsB5ZoBXNbsRL730XK+GegC2GiCHv2gPCC/YiZaF0Km8CTR4Ao
jGHr+3BeOFuHEmpVVNaioUC6BjgHERcPtQIM+8P8mRwpzlfW9us9+wlHOmPFiwr5WrWul8ZDaz7D
pHN8Zj3x7WSRZahSi6pDlbZbCtmYDXeOFwa0UmVF6MgzSdbOz/ow2FRwWO1Icbp5f4ndKyt6SCTT
WwWnnupbo/uLrjygncQQp9ZfbneciW8aJUOlzsqiTlCb8sB/+i36Vc7AEJcZvyor01MArhoPMyaz
h0jTctNJcOYrh+ooXX0d6BtQYHtAl68pVc0nGuYbp6f51uw5x//IPPUu/v4akd4OSx/Z2cMJRWYd
vfgm0qCzLo+N7YbgPiWAGbtTx78hemPI7zwEaMcfrrAPGexsgo6otslrFBtVNEN/BTw6i4iF26dJ
Sy0W12rY3cBLtEH9HBMm44h66CECbdMtPUilkezBYDZ/MjV1y2gTFNqb2fGNiJvDIiNXgXKM6Mob
YBxziZg8OulqjEZ/V6zEbuUhvtE5tqnSWLGqJtSqFqFB+pGWd7lrz63l3XinuyK7oxYMTWuJfHal
uQz9TT6njnkyBT1H1vTV1+RYQttJv3OrJXX1/PMlGbGVfj+mgrQCqJ+6fzF+AZO5RMrIZv+cRcaQ
AR4pGze5MeYpcrnTDCSDYVNTt8QoUZz+dZsg08Xz1KENxumGZclHrkcSNQjwN02EVlRdM03Wcfyh
JJhW/oJWcmEhB5OapCjwNBoGLdCKNh+ijPt15sC9OeuwK2BFYJaYcLjVgBftKB+SL6Xncm0l8Yc3
hLaIAag4LK9ynnqVmLBsDeIR62VGLuMQKRkc/zgdzPbc6ZwuePJ/fYCJDNp1prHlpYPxb3XhElbF
h4w1FmG1tb2wyh400vpsAEWIo/7t9CEby8P0Pj9Yb1hdwPUbuHcLTFDHAfNfBJQsPOuDaU06OxXp
S2HVwsW7lfPiEF4HiIwb4NpsQOSbAPc1QOjKlQH0kTulkb3LAQfM76CB85wTmLZysXohzpfz9td/
vi8E9ThttLISaZ0q8+ky6sVqm4s5xqCIwHnqVUXF3MNDSpNj5K5GP2IsLwapMqQico8EEWtb1RRV
ceOV2baRRs1DKgZ78Z+zyIga0rWfjxrrRtiasBiwGaef5jvVUzepDQMwbiS0oOkaYDdnMszglBEQ
+poFnID9f/UlcYck54nFwu5vyxyAMkOQL8kmTE8y6eeFNWh5iErJORShgX09YCMbLVK4CxwiU3So
78FQBPnVSu0V/AyIn+GY5BFiiw9ZP1wrMGVGXU9Ow1Z9tAHT6c7gVfThKJ3t8X4hOAdVhIHlF1q8
Z5HUjeWeknzXV3P1fzIOzsnHtyNoUaw2/OHZtJ/5hcDl/FKtxSD5zWkXeCPdzGIAyVuHf0BFyHOT
N79CZI6xuTGafogZn4AkItyg3Qw6jsKNcJCDcl8r9pZpOz+Yauq/w39qk049INlHnMH65M1bQ5Qt
/n4d/A3F04EsDu57LKIVo0BTbNBlUEm50yJNoGRYvZ3aytafzQO39xRFkl2tj3LYR5yE1OV+yyRw
v6+VEK7ghWhBj3j5WRNQMGtSisNF//TMQydUAmO3DnvyQharXScDDEBIHk7rQFommAt8Qcmo6wuT
NrQvKYzslIbphIIQ5ncir3hYUC7x1JzxUjfAYdBffETVz0zNoOFDtHww84UM9d4cldzkOX1DgaxN
bTjDblQAdzqCeVSsm9D7GBKv5AUm5hx8V4QNyUileCC/5/6V9MxJWwEhnXNKESh/CTi+cEbsbJ12
DEBzMS0ZEFMRHM+WETMLeA/0ihzqwpFWakbj3zKy4q5uf7EWvI+6dQ9vACbsnNJAC3PIMvLnjQ7x
F7JnUpnc6cLdslBxlJTCphytKyqpJoo3mLfnMtf4sYX5PLf/SpHC5YzIKuWZK80RUPjYh1lVnjiO
JyAOYKwIN6rrNz+RqZVcw8jJEWKapO+dt0CwRztGiUnbDguU5hWL51Ag8yC2ZlsBopoIG9/U+m/2
NJXtNHvvGU4xaCK+b+lJFoQQohmjEhsM8woI1EROEZqreaiDgpAi6V8ED8JF8+HhQMGs6asxJvWN
26gBdBysLYyffjbgiJJ0sPz8mN9piQXWqAb+HMsU8rlKdHeNTcdqqtgL9jbn0Kfuy61HeSV/mso1
dDiD4LZJwNhHK2bDc2nxUpna8ZmOa0E/OM0DY4tzeXLHHGfv23knDrmr1Zi+CYaH59ws+h3y5XLb
FdC7Xe5dNo2YPvycHZ8x++AyltxqZ/g1QddqwwF0ihK5QfRyev0qHsoSLFqu+wzgofB1ngSqVCqQ
rOO/Kz4dgfP2NZLSid03o3LbqZkNaVqJGB3IlVyRYJgA1H6XCZZC5zOu1ukNx4Y/d0D0+6ZGhF0A
6x0wBYRS+UPnTnyCrBf6KIagF3hyNW4hQAAJe1cR77Yqsevk9dufRc/Kdzi3Q7xFJ3uJk4W2ZsKD
vK/ZhzMBpgoLb8RZGE0MlVOL3BAquQ9ujUWRwjrSsu8e67OWpTSmy9/ZlBa541rdde7cJT432Ght
h3AfWxoEi0+o/aBjJWTaRvT9NLBMOIAh2q7bHJpQj5UZvQ+oH/zC4DW1f703Q0XVXNl2o7i+q9D5
yoAJVJzuWv4dLoH3nZuC66wPjhjnmoJxVO3YFeup1iT4S7HUggkWk6jB3ywtbCVfJCJaUkcqV3WO
Kq+PNFEfIEVAZ9PdkQpx0UX4sOWK+urqVcupBOmNlL2TqbyFyFmbXgTH8arwj2jUFVTub+zqeZDF
gN48G8nCc/1DLkFrCAU+11XaQMmOfwP9s/bul0+mBHSjvJ/R0HUw7QQKvwOigS5QW0vZ7drRryVN
boCG6GDRcKgw8n9P/S0uW2CHyznUpiuV1qNsLD/HKKT4wKHRnOz3AXJWe+6iS1nkAUYftmxIHNpY
bag1ePu5O5lB1eRICB/19lE/7HQGWigvNGkStXrPNBvQyH0QaUTHlkQLsmFC/oygnqRXQ59vBn/4
0zEMOXu2NGckl+vgiB16/UdX2eZwldutoqseHREWsXixjbQvEvI54+Zo3eeltNZd9sNbBIz0gEtk
Rw1dMGC/q2iBxkGXxeTRIGCgVBWtucXgBzVAruGfCKhX5NHPyxP6S23BCYIW0sWMoFar4tJupb2k
eutAI+t5MNC5PR3J46U50CggyH4oaeisLv6R9L/1nF3NTaFeY3NgqVrAnXJeF/M6r5wanFbww1As
YzwmU0+9hkxtSQbzOcWaUAiLRvS7SccnsDbQO58WjqWT4GtgBgCnSLvRDJpbKLWPzF7IN1geLXpe
Bt2qi3KULC54SXxFMMJTvTLyWD8BeCZ9mbsB0QSDUnfqQx4OP5wZSwmvxgX5Xpwk7qw0NaByUmRd
Du1X4rv7Xm1E1WN+5ARGzBTMkN9ojX1D6KErvbzl/AM3dRBS9YOnZ60Hg9hk8jWZvs5XxzvqJnsO
YQeTxeWu7/yWSiHHAck9u2Q1a7dfOHTvlDkaYLYK6RsikQoHluD7PCuajsjagHlHgAsbN1mdnIsb
9eNRnHG0EDvCzhTGe2KDwxtRUq7fXTLlplz+HQwAyhtHl0vkTUQX9Yb3Br/Khqkzw1cFUV02KMn4
PDfcSbF5B34H5BV7b/8x6DEkg6nthVIhMPELeIEeJ5ggFo8SZH9aEpJsckIHfSNqD4i0VfU8tZal
2Jwypr1EYkjgTu//p452vVL9BUpT+ikPWIrVlg65LMYirFkAGz+thKoNs/gFZI4QphrpWtMGNWRd
z4G4kIwdAIokLTsFG8va3rJvTQsQ9Mxo/8JT14NptcrRzkKXVYnL6PKDzCevSGbm9dseWKDIARc1
m7mv8O+ymb2roUOhWiAVgoHfL0ggZVT+0eAl5ALYBqmMZXvRIXegcz26gGLza+1sr5UPcv1RscKp
KYvk43AstwTQPDjSIMH5GPW7FcNQCiwg9ergiPP5ek6lyrDtSNet9CACHaoC3vazsqEHFCzr/3vo
SfToUtWQ5OqKAeZSmejYPwMXuVsnA3ExuCCsBxkfiLn2r9zeFnKhExU0xRrgWafnVQPU7vIj1IW6
cq0ggLoVMGvwJLaxjVIru8lBW8XZ4p4IEnTScf2xpX+EmBixrN5MP+4vKIhuWty5hwHIo3anEPdp
zIn2LK5pczyBUirWhVHFMVWRgq8iQN16AoQ5978iohtJDWpe/Cu17aSjTXa05h3KVLnkRfT67Rj8
ZeGGIACBJ2hLc57cgLhwPVcKrawqx8tGbc40J/qXmFPq5nOtquPPNAIuWFCBbMLkYSVAsebk8xS5
7HWVspAZZB8v2o9+YREXGVNVChe8rrKxT37TaVjIAPBGMiA1xan9Iu6yXIViAHTVo8vnU6MbWraz
Fe9gr1D8IClCkdabS7ggrzwCTLqP/hrCTk1o9W1x3VzdW46d79l2GqWCxJKi6mePuQVEMwQYWRMc
p9nrts1Lfv05N3OZRToK/FfPNROrnwN/OUEC+IPuzCsjFG7/R8XjkcRiHhnkwWgjcwgRiM0hwdhp
jYtkSASq1A+/vVkBC9LDRsoDQ8Ro3zNWpD4+pWadPPksJTiEQfhHpxKnZeFGQuTp9Kn/5CaI+bxW
hLHQz0aKK6jgIOZtO6P5ZxuNVjTQD7ApU80ijNxzs5lmKHu4Yczt8Bcjp2n6LEm8r1x9LFsYFE1k
EDcClN7+qhEUOAQxZiX2BeG9izDLwR0BfZrEcBFm48OIkDBtAqO4yrMT4wouPjgs3Q/Z0AmZ1ioZ
eQa9cBNMw0vWLrJ65p9E6wCOfYN9sxGXBHEDARlpx9soU90+AG5M6+TWuPEOByk08ex/1INgdCTW
q7H8BVDQfAWfeNiqUHrp7wwuhsPHhGFjxbUw3QEO49ZTWcowc6Re4SRtL79CKvTC9imGPZRkp4/3
I0NIcjthtwjU7Jv/XFhHik7VQNatOlhl3m7xNAkzU4nWDKCdM+/TevdXae/3pYrGZWf8uN9OdGiw
yem92O7ck13YscAdIdxTjhKdQQOkQBmuALmRz+8MDS8r4NkYunp8nC6xwUEZAM4LC8pdA2HUiLd1
cDqL0GHEGPcAeCP+lfPwuHMlfSVuH0XggWZP/uiYNT7Pge/BIvWnR3rfv/Ag/WCPz0BvQ9oQ2Odt
mZ5CO7Luzjdc8aTFu2W6L18qO9fgCuc3ZFtpOQe6ApmMxe7ubxb7FFzb8hIyfZg7aGPCPBJLceOo
TetkbCZH7JLXL3xHzc17XgSjF/sJNM8F9BFrNH0fMOj3DCGZt9TQMf2JJbuBPOyhFYo6fZSpmRrL
/EfsxdtpOKOBgpOnib5tatAklTM/KGthbBa7R5NUiu1D06jCx1Ur/nbtjHw20jLf+J4nDQDrJQOm
0mmKSyNAYlco7S0tbu6eAQ0S9A7j2wqTzHGwlozNd3lv5g9+UXFYjnMd4DNwOnkVRm1xJA0C4gQT
ksi/K9NM4fdN72oqYYIulNh1wDTFl4qIRs5RaknGl8YeVvGEldMhqKgsGupf1n/+iLz/p4CxFvn2
3+VvBj9Oy4OLFyL+m8cddP7ZoQq+BhgP5OImQIe+aiwdjPkR4x91xjV8GuapU4nM3yb493laIogT
RuqqNdPib2fz2v9YJjQyhIOqJJ4FOS3Y03BG4wDs8ZN0fFUO504d9ozH4Z+8jmkH4mnCPC6G5s9p
NuhHUbF63acZyXCfBNDKZMJlY/LhfDtSeAhDJ+Gdv9sLZwNuf/f3IpqvIAe9bqjDQXMtaiND8Lka
/bSvJaB2uemGxSjEHnPD7+YUZeS0jOcGto074ECfWZK+dQWXltHYjqpVHYIZxZL8AIZ7Jm0wGGj+
+YrzsdM0e8VQkOYAszGWeDP+0iudIYw7iRXKH/RFezZbgqYTolyoFdPvL4Db3OlqF9HiUe/hWSPL
7jVIhGiXd6vUybH72VMAI9wXmuwhaMoErKkl8Dpk8W9Eol6gdrPXSHE4zfmKvl1d3Rb9GBgrNKGW
xvrRI3rINvQVtz2YcILuOGphJCJNHbdG+K4+eYJcQVVry+G+jIQU3OZX+5QTvaA5ygCMxJcLAsHu
/+q4bMTbam/6SIeA3lAKh+1uS1yx7jeLT80DDMMhraAi9GR1uBk95kT/Fxuv1ShDrvMVkOu5ZS7W
8nCbP3MUjHDRMh5vDv5WTk6wkfLz2y5fPq4XtdEQudC7a7pSuQPgdEQOdPp3/uqPst0n8iMD7FgH
yYEsTsGixI/r9dVKexDlZOnym4U4d1YmyUnXPbvbkjomG4y48spjy6Wn6xivxYUYhhNmAKsXyxWj
b3lpXNAd9yKw/27ef5tXcCpuWSBFYKsysj8IFvvbnq+N3FLNrbxSnQlnMm9SZk92jir8jn1ucFb6
Jn4JeEqXCl/kPwxKKbE1ZmgSM6/eJMd6HIyeKIGWy/x/X0CLj/fyXuUq2svr8uMvyNgaloZ/qEyp
zmWShXOlb9TYcunihzUDn+emU9d0v8cu0qQyQYf8s4poUBqaG7B13ekW/9Qfq7XEKn1Bj9ae1brE
zbgmYHwaEBHUq9Umot+g1xOIAB2mo/rICJ0aeLFTLtN2ayU5qrlUc0c9lBMTS5Cg0uoJRGnLwQNh
G46eNCHHM8Dknct1Xa3Djh/+7BZINGN9LCVVp2J62gX+uy+RCJeW+UuVVJ+CNMmOB4TkGkoY10qD
GOcsU8R/NBdUlX53uKGW5spQRCvktvY4LjeRRDl8xIOg1ROm3BEv6XfL6/Pa8Ib3Yxnonlb8IOMC
8Sy2iSNKq49SKuA+u0vW4mDv+lceevAO6ojpURgSjDKaLDeIqqoSsyNsIauGJyoVV4SWv09Wd9BJ
9sMOXiFFruAemKRnak4BvLQvZ2Ss/AuxVgNzG8rcg7MhvYB1ixREQgsaqkU+RxUOf7RtCFTVHIN3
kEsr7ZeP5o1ZpkiUwI/kHQL2RxDfdVhJBpACYIoQE25vIprKguwOreVe/rVTzocMR47E4A07gsRo
JcxplJs2OQz3FzXyLJhhUp5HW+ZtrORxnE7HPcdqT2EWdIgZ+vfqtgUazXbbEpGC5xKGlKgfye91
f00ZCgObshPRVp0xCX1bEPbqygtxRizL1ttqS5TOnpnot3kqdvR3YmXsytUl0fuJ13+R7FBJEyRb
0ibYLZJx8yd0FVz7JK140A2JAGtzFedbcc/G4gD15UXDEakZWMZaNcHnMkF1Y9of2xllDPQSLnna
scrnFt3n9L1bJ+WxxcfPoEzxwrdwWl4cEaWU9QNQdYZWNL18LhYcknAKBQcVGMTSk6Uy4r+/TWJy
aHSvbpAMOCo27kXZcrv7CvIp3/C2+vxYeumVQRZejAi9Y7o3eOX4Y4clYLnTmo2iWkNJ9qhqhYfP
cDPudU+owJCdhvSL0P9o2cq+fXSsnaUJQA//uSasTsMpaYS/E0mqnwfYcW/Fw4IyTuVu8uOdA64e
mAYoYr63fy1y5r8qpBZIkH9y+33f0bBJUhjzoEk1ih7dYGC3pJo7qWNZz+7w2E5Ow8pG2Iyh4ukI
s9l5c643qg/LEUgrsc7InftOoSogAoGjQ0RiHO1w2ZQU47RhsynXedmMxWEPC1K4fxXyyu71gCbc
ur3fezvclb8Xwcz0E4IAvuZ1PMY3OMyGCTB6pYNDJ3HA2dVZMxy4zx0QGD3RvJahQsvbTlJnV/6A
/Uwl2heRot1GCdjcdCQ6OhCXl2w2ApWvQ2aCAzXHjSvYshuXMyyUCsAcyxy3rH2KGt1bmRjNRcuq
9/HipUW7jXsop6QZ44deYD4QkTCuLzfXXa04VXu2qOCAFOlToSGBssak0sX5pjxDZQ18CBMsVpsm
D7jwcXIHW1ghqaLf6iXqRYTFStmmL9uAQiBxf7Cl3AIAMbapkX2IQKS+cFY64KUqVL0Hws6K3J0O
VXOWwzixVctFve0QbgFfthhhS+jU6oHr2QvRsO7OW6YcJlG5G7Fwwen7300fnQ0NpwMHSzxdqAq9
rxVml2e5brHl7ZMNKGMoFYBGIHJEmVGumnl9wZPQxvOts+opOl6h/GA2qHS3ylCbRxelZr6NT++o
2B79E/Of0vI7Y5TDQSeyAuiGunB5Be5Mn5A3c6RmNkGbNWeOA+czLnbgTNI3FBnVlxKi3fCdIMH/
5ikohgqEeGUASAl0UXaRSxDw1BgF3CFSzL3KT3rLWLLutqyuhE8Hjzx3Z7SQ7VaH3xonKCEBaxo0
Pxx1z/mN9LOiV5k5ANE4UOAqdnIoxMjxDei7K/evOikU7s0a0CPFGfTeWXMXgFMmeO7jrOuYB0JP
xy35Nbqun4MrNJvaKoru4vpVZFbXPFtZVBEycqWAuYqumE88grD/BVK/2IYl4Myl8P/U2qqHyKzr
OTBTfdXh5m+Fmp3FtwymncfDhElv4KsLdMe7djhLalKsA9CXIPioYwe/U17B4uPhNs1mEuPvdUWU
0pv9AhbG48KM4lz2HzfyrGhVn9HOrQLHkH9TOyied5UIY79s0nNTFzyBoCzehkmHrYXAE1FrNFmO
N290QYKUhPkOgX2ct4uwDF70KO6eqUJvC+ePHy1xszyYGVujAKvkSdKH/SwwLnZt1A8J2sAjdR0K
cHGwgNfw7zGZwadWDLv/uhiG9ny09gwVO57t/Mp3FeoDkWo5NmUHds4kTjELkGMYnrOdx5rvyhvs
/QpSbNyaaHoHhxejTfN3pFsxYnPOUsPmi6GOmFZmdxy6q0dmpoVXeFWTdSKGVEcUgqwLhzyFNIVu
MVL/7RLRtTAo+JcX7JpWmAayCX7HcE9QUJOCEdtHDcXB48xBwBMIu1YB35AT4afMp/cvC7eHZNhD
jPxfmL/Cg+djfbWr545Vj3JV8ECuy6v69c5o2ZpFF2m4t6ht/7uvGt3AwTUn93+w8j2fyABQwv1j
tKZ9dbmaYsmXirYPz6GShGnKbwkehKrjNI0t/R4tAudPj5SS3/YjzzxXcBUk2EjUpA3qMKJZTEeN
x0eZjhtK2hRAjDnOmKWyRbRg34BStdlKE6hiq6VJ/EVBLiAvrhoUjEqO1LKABAe5gLKd6J76tvON
nXUY8GCtRmpie5Yw9WF13YEwNC1Y3/HIMzN+4c9LBPDpumKcDabXMc10T43HblfitivInlgPxQuQ
iQYzsI/P9ZpxiMp3Y0ZbBZH8rWIqjH9cWbNxW+Vj+kZaU7ttJMf1MQeJHMIt3IwpcWRjLOCe0WFr
gjKcI9jdAiGRigWLcBxDx6/j2ZXMgUQEmwU9WJLTK845/y5sekGd+pQVXT7XQY6ukpB46/stbog0
piEpCzPEYSIxZlv1Qsud8egpV3iqvm2RrtyvERd/luyknzX18kMXffbstbFratGeRTQpJbAZAH9h
Vy1DbdhkvyG2y6514AgTQP7wnjYYWKvnGRavPL6KNs3wy/rQ8CImdOQbOIcz+D3YlJzav5C+Fkhh
Wcne2yYwutcPCNkW+8k6dccCCC6gh01cpVsajgppBFSudOelUdPgQcv0Q7EEhcxEN5e9cJAnf+TT
9ie5/RzkdCz7ep9cdy4bgnxjjYd61oyNFwCtdK9hIYg5zeI0gbwwcTI/BNoKBuNgHt4uGx4EqODQ
GCCG1vY0hGSao9PHEphdSrchV31oexH854oJRIUxiyvTXCbjMPCW+o4kP/5b1wVeqVdxXwsNBe7C
NV63QZtelEc8S/Za+4V94rfL3L2maWoxtaYAMmaYAJIZCeMeIQoJk4N91MSJShsVSe6wL/TaGpWg
ONL08QoBO3Fntn1+Gj9FLlAaYQsbLcI73VXAzjS4WmPP7URjpF07oKOP39cWbQHn/DAa3xJl+j8H
P2J7zCp9nLMzrgAcNWXm7M+pE4vQaslOeYDd217SwTSCaDslYWWDHaYyw9O4Ru5cFp4gwrL81jKp
W91se7YKsyNEYdUFJefCN3hqTeocdw0AVXSxfOrIzFWL4GFKiyRrsAKaQBtuigTyNod9WyS4IVA2
3yzcFugRusfi1RfKge+rh0BtonZDuaPBsVJQiKI9TWuKcAjJcR/lspiKHlRyZOXpHedw/180mpco
LnY8KUwZVh0lYIv0aqedMt1nUIsfDaCb5Fd7e0tK8MF5HznUhdWbccbZhHDI8plSHy2Lr1EEmaUG
bbTi/ZRPLsUIuWv67VoV3ODqYEB55SA4XTjPCGgTkujH67XiezxGwp1Aw173LitD5NuGS95xhWnC
eksyCrHvopqwLDinx+0ZY8nFSCiFDsYX89mDuX9chgNqHYDg6agoAJIqIrZ3mspPJixrfds25HBp
H1EtKr80eadcNGikX0J+wsy+gITxTrVKnK3SkJ//efAT3WN3rY5tot3G25Ix36A/Hlq4jEe2k5ya
NnmZqxH3C0r6Qvt6/GRYvJ+guD5n4++cyenqE/i05hn1BhSHLUwyu6bHtDsFAQyb7twMKNsnkkRM
s7McTYCHKY5DiLj0AJh3/p9k7fWct6/sb29N69pZMqPCyOZRecENqlIa4H5LfjgubH4HhpY1n/yr
3H0k0j+vMiLGsBoPr3k5JnuA3ljGhJydwzswImFdMvIb7P3CQIx2bu+qCV0GbOcR9aE21TsnZdhr
tAbmaoe1dXQbo3NzjU74Y0A+umdH2htUKXcCf1QCcFhlZMIdJIjjfGIE4+Gqp78hQDM9MmvIA3Tr
4S29FRI/qhRVAx5WtT3CMhofuRPqKrHZGhTXSLSfB6S5VYOiUmx72TCIVKW2Om/o3KigvQlE+skY
GvrJEPLyhQ39mbb2G40gRWyJcNnpqdBpQrxet/aiTmWx0OjoUM2FXqKp9hWsBsXjFVuwveUDNDpB
28N+XZRzH6BKRU1vHMPwHmjSsbo5DFZfQvlaMr/NQiGVVaVHhYG/wt/dCwpnZZ9Bb7Sw1LBv/86O
B6aEq1EydLMuaf6j0ewtuGlsaY4fM6PmI8G8FEy7tlbSibi0Cj0PZ/3VAMMhcue1e1HwoQVePkjz
j5bbIFsRsruPAjk/bW2hcsoegdOE6P4xc0rZGuXlQBFU44WyAwLQsfXFBRb2pajpFg4p1L0/jtVi
GHweL8if+mRi/CAunqdhZL3cHdhothvQSTidVGqRlfGwkBVTTXfYPl4+G/xXjvbfF3MTM83zNbCM
Nq+IMO3bBmcsOGl7RKTFtrbUb1lHh3MpIfTkh4GnE1MBalo6UlCQCRF0YEJ0RRg/HuFVZCratufO
wlSJiblAOoM7ZKwevIR0OSo7Z/8imzF2jfsnMXAaqNEN0czHiu3wi76jWGWcC+MOdGU6q4ljFwTj
sbzmRyI2V8Wcv2jcbkhLR+TDDbRFLlmPoHsxVNWDstBBXBu/5DN2/Xx86RkFqS3fU1SdggNUZwBM
CQxaxw5RllxEWsk7oZES5aUxhIKUxGdAoK80RgLyqn/6ARuu7VINanmNIYUMYIGNM2a17LMLVFNX
83YirlTOuJ5GFKhdfnJ1fmm1GYV7hCgcUOiaH75Hksr7klz0reGnMLwy6yTQY760SSImGggQquNi
0pQTo/s6kBCNjEzrz/rWzF3paYxx8yPNbgqAXECfRknL0A2zNI2pNgKu+O0MKsm7WmAKFPKncsj7
xr7xaceJFcJ7tRsamNuhWta583XB7IJmOdGYnBKiMqaGbwKdMyFSC3wXJIx8MfdIZqc+fGp0+F98
GKjCRSeW7H7biYDjEv3LZ7SRys+gLGM6q8gEDJpdWGq5EPTkkUkXkL8nD/Q888jZxgUtN8/BXkzq
mw4Q6CS8b5C1fpCQkBBDDjZqT951uO7rNYYpV6tUgCXRZ8jgCIofIzBWCkKREbpluK/hXFhAdy+E
HQY8/sNQEq/7mSHu4lrfViP0RSYac/NyEcACe1Yw6DxvM8MQTXmbRhABaFotU8+D+7b+i5nqWr3N
5IfS3Y4q2gydccxrDqbST3SlsS6YmsaN5oEMV4uWCm/8xG30NQUvDPIiDar7+rL45sFY4rxwN7n/
Nb+sj7VDgqc1/vREb4kWfGNvCbFTrn1ykZwsb1z4fXEOvNWtKbJw186AYbcRtKcGij6nvPskenNv
cdiyeFmaeg6FONfUZaCidsUb6rR+AEkkNDkeO4JUbJLssxvTvUANRtPVk607OzwtIybB6DeRBuxx
a3+5yuJd+ttyEh7xaznrcgdxhoyKfAshPhbpTugE17g94cDti9r4UVo8buFQKyC0aoBMuvlq2JgG
P0AMX1AiGwVtvk3tfw+ogihXACQgnh+qT53RKJqKaGbw0CtDHY+30CcULf7XCCZBOL/qJYxmBjea
nYPiZSl0NWwQ4r+j9VgbIPMBp4IJdrYdGR7AuAAvwDyd2MazSjHusHPh56P5NXcNEqfsQqz9MdD5
bBH0EyM/6RVHP0HJQ90/uJarE70NMH/WAhDfsK1aV3MH2ZuOLisGGqeZcX2XtA2ug5n8tcXURDPm
tGo8jxX+hvTKmLLEH6RU/Ruy9KXcrZsQMb2z0G642drcTcBF5pMtlB/VI219Tpnrl4y9eSupnqzM
N2uNNHV6rphRyP3KNYZeF7TrneC0s8A2+4WnloYZ7xgV2JtUIJUakpJwgIUuCuXDnqe13vmredTe
3sly0MxQZ0Q8N18d3JDxeeJNbS8NrBVxXZmht2FPFGeibaXYSezGFqwrTxSAvJ24V4tFr4unujnq
G5EQ8W/OYldHiIdoaSPCQu1FjZrDdohSYGWNI6tAc4LSFcTEhDci9X++SWCurfRgZhFfv4L9QQZf
s1ANctjAcipG+pKuO0Cy92Bf18UenpbUHxKpbLibsdPG+BMyc5pQRIbJ7GfVezkFaJ96KQjGLBwa
gfpk5sE1QBV9x0HYXmGGwyCU81/+5whIchoPKlN3IsJWCsM70ctjigxrkXbA5+FR/ib2V+ly37c9
kDVCjO+d1DP6ZSWLXkp0bft93WPaXxlAxbZwK8bfuMjGjaqYIF4hkkAyYzmlFDLuQlDjtS6L2nQv
qIgO5IPCkckQqhTG8SyUhCPJpWlA3Ot3ez0JndD0XRKzDXEtof6MgkcektBieiQY8CPVvwmQHBJn
FplYKpdm4QsLi+TTk86KHPfFdUVCyia/2qnpKuI6F1668a761PG+Gt8bjvYbHg/XwTNGbN5htJHr
mVuoYoQRRcvUGKjSMEOTOTrljbMPnpMDvf+KcMgp1yuJy3CNdqr6haom5LjpUCzKYQCpEkMbaAKq
40cY4vBFpLb7a4cWDqdhGvlfCWGfRd0tvIxU5Lp3eZZrIAWC4cUQmQUDNkizZyMVj+Tien0mYI15
VaFhfmJai8gc0k0s7Zsf6hMRWnlua4UF2pD0f7hQ8v38bzK9YDqnpATkrDCscgkRrrMMTJBCnhoy
/NAth106xWkwmCo6Uzc+uZky1qL2NuFCV3B3207dLyOy4pAeJVYK+QwHtzIxmjY6N+ViOBksfLyG
ZeRN4mJSwrRDQa1UYRbsLL894u54F1KG5sK0w5opg24P0MRixLm5Q9G1iOW9vWlevkQXyMjRqjwD
wc2KJ8QdQNOZ93PO12dq+APw+DcsqbAS9IzZYFFuQiWLuhM7ELwSy/vFoQQZPjTdJfMOjxiMxlcc
7YONlLO1haEpTyXMOGAUr04ayDtEwv+TkmT8YbiRKPq61AhHximybe9cQkuiTs5YtZojf336Nvef
IOr7gEhl6TIHErMG3wLnUpuAZo+Xcqv1QIret+G9u1+CCsdbSVe02wnMxfCVGbDM0k6Bx+yv4xbU
Yhcabn5Z3i59h87BX9aatKosB+AMUThV9EAarpfeh5ef2w60BjKkAY3G8qPENWzEPdCTALH+0LUB
aht3w8TizrC8XfRB+rRkIpLCgAJL3btNhQssKVGeSBeZ94uadXVTdkm76I463UqpiuYEtyeA8uMy
wk27XMoUoVEymBBQeVQNl4N0ZRMLlxMg/4fjuVZNWkIs4X/r7iGsViQcA082wx8ZOWQmpCq72xOl
qfWYSClpzePrq+QrdWpPIaJDKvid2D2wkH3xfR9a9k6SGHCTO9aXWJzTdEqwTE/dMFaZVCh44kBX
+zDn8lowNqwEfyDiq7n0r+C0i2f3Rv2z7AtW3stheuvZkvJoCHrItABzfV/SbEL8zVRqZUdmOrEE
leYeTDfoleyT1smfBvK4cCZy+osit3o3uK0GravmGygtPBk97EhXV9j8RLAyoUeG8mSt/aqkGdOe
ODRuHY6zcEnbqfnohvgChajnUNBoBKTBqqoRufdRaAX8tgFQbUfSBwJuhBOwlZU4v8pRVsZp8qx6
mlniFRwZBZzKq2R3y7bn4R6ha5xsbv9aJhsCw+c5uXkFdHUtgmj1himTViPWYXU09wZAsjpAqw1R
GzY8oHneGDf8JwCYcSfPmL7KLgbqQsk1ToG/dl8T0bgF6TgY1uF9W5mEX3FxUeAgdRGV4usrRELj
52wcYg7fQpyD67QVJuDXo6tgBR3DXF1fdycx8fcHdsh2U8FI937RO2ex5n6KrTAr8B7cXJSioFVD
cangA32anYq5xnCkzFNtFgb4e3cb1yf9TJ/zC3hlRxODwU3RCq/KO6m1RYSnrFKbQaWczc6Psm5P
p/3k2IsuXWdsqkNPvA+znecpuvpJb8Sm55FOpLqPKcrI4xWUHIdicdzdVMBzp+mH97Cxn3+XvcVT
sniPJM/yA1lgyZ8zPDQu/90mbVO/lgGzQcvkPh4zU/SS0zwLs5bQMBTJCLWl8NuqmG+GQv7TtQ7a
ao1Ng5bLm+wbQ4qAy6M+rjwfO46WxDJ29c+xyR3/gISBGfXlagbWBdpXzyIX/fCMOjRH6t7c4LAe
6tjsFBJGJYgYjZ8pir9brKvyfGEiGjxzp/aJr19NNvSisunMHxIJB8YPluJEt+gVCp6GCPzAz57C
z9+A/ytHiveSh6mm+8w79QAJ5wa8kRLgrzKZlFVX+NQVP0ZVHb/4B/kOEd+TSELA6mmPV7tAnE+F
e0WoxR/cq5u/K7o2Uerd+xw+E5iv7+NoudmwdDj+jYB+zfl2VYKJ37hfrDCYorgxANaqOUVkiHQ+
7MVwDGOoafHtCZ0YUUWpovuSSzle8p/ZGRRGhm262VQ9agVF2TXb8WnNRT1uvbJfk+6j9BmFEx23
bpgSJInvA9tYveivTnN7N3JoZMSl4NvV1xyOjY9qpX0yrUSbXJyagnk/cV+MH3jpka4gF5Tsvbof
2nTvrX22mXh7RAVgK4kpHxQHFd4RFEXY7RNuKjNikfQCll2tNskArfsLkcUWxvaCSkU/Q2pyziY9
grJvodZC0Z3KDrBrldJmeh+h2pVWHwmRZTqV/iE+MrPG6VBrFuDjrb/w3Wls6TNkz2yBS/SoWa3A
XwTl3aPo3PoS378lAQi2hAiz6ZpuIyZ4/Vw9zZSx5fhiyaGDOruTfbL1PrsOUkn+EQK38pVO01ZX
9ZeU0REstTlKtbC55omCNXCwGc2AOCk3uxSiGV66Z+DXYRnnER+91WBoQpBfOUtjUmwtDuKUbtic
st7uKJfYW5HpY3ETCmGvbhqmABXl6lGq1CVHe6DlUcfdFZUBNnNRUlT60zq99erxz8/HLxueOR6P
PZlcZZwqBH3Usg/Hs8Ngid/T1OxVJRm/ApgHSEI9vTedpeh7fBqtkGgRrNcxkyVd61HqNWRIvS7S
MDvwKmZ6bGSBv3QOAOcbMXgzwk1TmOFnyFk5UoBi9w9xbqqoX3uM+iFMuf4Mf9lAB4zHpiLENT3M
J6f4idOwIjHGYd4UsDVSeEH3JCOszaxD7lXHZI2iUFgBosGiFDHreBzuaoMhFsQsWyf8c7QSifl+
pvYh4xjRNK6BJGNgYcX6Ui4t6X69jbdAXY8zYOlyAoyLz1PIOSoP7QJfIW2Y6FidhDKZ8fiVxZvz
LJgm06jAU6Lgc0TENdEQf2s5MGk/0zo0a1xoFO6XfLbIlXghI5AezWADJWinbVncMjUQhm22PpbE
gTzC96hCBDUFjua4fGHmJYiD6PEy+R6fRJa4gdpxlKB1qvYo9tt3rXrqihulWJHn6RE9XeE0lswJ
IT09WPk235ff6LraXSjQp8gTia5EL0k4wxqfi4xXe6op5ResRcT7l2XXGIgqfGtTSVpZCqgHF3YJ
2fjMk28lXnrf62aXaCsBWCK7DYzB6o5XNnVVU/uhiXhS0jkBNKTSj7uc/Ueh91Pz9qoQUiUU4U2S
QpaKr7Af+b10goNx/9BLqzWN8cusM1DGDM7x40MStGdqTsvUPn8EMR6/8UIz4y/hLQFuXZ4w58Zi
WFRvH6xxlw1HZgG5EMjGKuniY9lYgrSfmerD+/s/GU+FYr/oLC1xrt9WHu7ZMHYkNiAeqKtwNtKT
HDlapzTc2pGMhwpKnc1lquxZAWzdkk87cw04mTqda0xyDMMwF+crNxVv+sKUfVx6B8KAdHm3Bxny
EDsPg2kXTtdFhAm3o404H31cwtMnXwVge3VvlW/jrXeoz+e9240+dO2clEyKpI/sdfsA/EWKwsPX
GEF5RgAawY/8j/sqxTpc1TxXICxMpa83Uo832k56wTLb2xO/Y/ybsEqc8tjZOciB9A6k+Sd2SPr0
9kORdPDtZKJuRWg1M7SBnsf/YW/XKnjmQlUvGaj0hAR8UfvIJ5K//QTM1g5arW2uWhVDV42PZK2y
0OoYvYa5oBCi2yNXo9BkKxKeHCjShNa9vNuTw9yQ6sxq8sBfLOILuXtUYIvC/fkoyVBPVSuoTMGE
6TVNBdRP6bvWuIiWcTrqfG/bAh/z/N4rUc+aVOnvDz5irVAMfPd/jvCLMj5xKnO74RfhDwbTFAAY
dTqJmyha3tuRIP/76+4DNQKNzZQpyqpklOEywWC/7pfqD5a0MqBeAHK9xfJAqqSyQg85uDbk3n3v
etpfIDJK4H9ZA5oO3nd8KsXExShEDcLvECWhhXWd7pj8E9c9lqV5zy5JBk5YGuES2+P1dsOlpXDT
GJCdtEnZg1oLSIOiDc6hdBtlpdnrMaDEio91Ksuwf4OM15AemXHp8GSidZIu1oz20DwoqYU+6yGM
OCIqzW++tKvvtmG3Zkr0cnUdppIqWHUkfLuOb/TmUnfcZtD3Zhv9ioJ+dvFVxPwjBppVDB4Lgueu
k82qPKXCIcsAHE1cy6O2Zl8TA1VIeiaTNkyrEopzAmsHP1GCCstnmKWx8TBgdghv2Ch09J/Eowsv
4C17JVQvocp47o3UL72xboWhx3uF70Gqxg/GIYDNvUGAvyJS5UkettiQDjNG3mZy5AaPapQ1eXc1
X0FdIVIFJqqgerDKJ/V92PZXsB1+dvBlWe8xWPRbeejckuDDkQYqyXsrw/I7sYMQ/B8IiAlrmtXT
+VOJzYxfgr8UZk9yuFa548xIdJSwLQsojBZ6YUcZrIdJKf7mkypA/YEo4g5B9/9AfcTEKDyLMI9n
gI6bNC6BnBTbiiZ8g4YUDn2Q/sT0aHM6msFcpo4qGB4/kEQcLccxmmbHJ9bhz6Dunqpw4Ul8PDcS
icgXdiYmE09viqzhIxuq/gV5bR7qQSL+eA6Bf5IaLAKQeQ/pTwH6S37VpP43zKvdh9hUlnQaC/g3
sztsCBF9Lp2SlMdHB2gefb42bnxJhmRw8KwXVE/4ZnIahttlKQRSqZhLIY3zIzzBdcotMARd4kpQ
c38l0282OYtEEGfSfzxFwYxBO5WiUta1/zoHPp5mFNV8ZMaDcJIoXvyoYg/DYJ89pvtSOZ+MdUSb
AWSHz5h9xDT6DFSN1v2AAYXeS3DZNGsB63L7+F0X6DhoaVhOCFoSfbrYu2Sbn/p5LfDrcsvpcUK/
UY6N/9obhqMQGmia1hyxF6u9lzbyy/JnN4hft46w02MPaRznhgcgekImnoOtBHmdmpTZJMIQz1Vk
AnXkkynjVsOsFV3Z2sUCW6Ut5a6fvAlG9cCBdugI0fLOCImUoPgfoKkzOb37am92KQD/9uv7NK4r
ZzDocGM6cTu8Ti5mgWA5MD/vAGQ424LWNc/G3vDlJIBx1wLL3yJt3VoiMVg7thxSXBqWWtLgJ9jX
mWp1HdFgfpBrYJqOBk90lSkCMX0ekBAz69x4WyL5grbgGe6Sdj6b0o2vu3U5CHZMZ96gRsrsFNfr
M/a3B3r0IogSWoBx2f7xdLBWFAJ5097Gk5JPnvKDtl6Of+KAhN9FpTQoJHZXC3DT5gm8scqnJVfN
RROuhpMWDIBpzjiPY0TS6Q1FeCrQyU/P24vN4PK4yMFBhePsh78vFXz4bmoHGfd6+Qr08gXNXA8w
nNChwdjrXm0BH0r/Gk7SIaCP+CAv57FzmcMLkyqM8GEOGuptnsn+6ndYe9m5Tw+Awn8vKvvRrlJx
o4HF48GKQ2H7MXaBz1Sp4dMzu9rQAlFZpxk/8/7JM/EPkrYyqtiE0arJl+4i22P6VL52S/T6+wD2
agm4qTR7DyiYtsuebZUZwyXAKBLCz/41xd4IPONbjj3yTF9dIy0v2b2zs/rU2PTeHhoUlkA1MPpo
8Lh9SdjC1xsRF2qduOq8KRgUbsNlemAG83rlEA5ycwPuJgbt0bexotMrYe1W5J4zp3KmoTdE4jXD
3Y9SvJrbihmZALZt03Lo34l8cxVwse25tU5JLm6+KT0MJhcKrDcweugUwo8G2sVGF2IK4iSO1nPm
gXJ4qKHFkTvrVqf/QiA9XuLHQ5MDjtwBPET1lo/1xd9Z2Yu/UcXEwcFPFZWL+cPCP3A3bfT0h2in
EJHY+BgAl0M/5SQOxDVIMk/fibibrXmO2aD7e2sPSlG0vddKfNEG+303Nl7y6+X58oDI+QBi8IhA
6eQxY77Z98/F74zRU7zN+kaKPCImqsSd5bgqlhiidmWx9afFBxB47pcQWfKcmCdDagmfG/9bxQcL
iR5DZg2ROu/2qPkqJE3eIsrP2EhvoIqagJFVk+jrraBverwwyIOeKy3b6PenQo6+ASpEaS7LFYa6
Zibyh3/g5Vpa1hsIQzbgJ4oG+4OmzA2Q2he1UUR3YHjEshKuqbt3YETpGqkg0Vjz9ppGEzcgJ1cu
WbPiV82nSeSvO0dvDnWfgLxVS2R1Jkb2W9fASC0GjVaCmNEihPpOk9rB04nOD/ctmJeQm8ptfg1z
bSUlKDRUnK3hbkvhXfkB40DZipK+OWx5a9P+NH6CpMdnJi0QQdgrI51PTG8GgosYCECB8Fe8xuX+
FfMWXO2O3MvWCFMnq2EAgZ5a04YkJMdpHa609kQfP/8IGaG2jlb6neBSzLNXhHYW+Zf0I4FKxHBv
Xt75xzUBi8mAoq4vvEfPWK/Wqk/RVJpp3i+1AWdOFQuYjyE2frGcyJKYcHxfzDtg4WLbaGGJ7bhI
e8zBJ3HXqNjfWgLYw6TurD7l8wrPyCt7M0tZqQcK5a59pIhatHfawoX+vmgLQKoKwPIgCnOPVhDE
rixsArQ8ZxUhX9FupT4rkMjMm6xGeBjLLnkFFZemQO+atmOZSp1SKJX0y7fqWjrDK5FmDZ/xejtx
1Ls64bgN/hoDaF4yHOPalStHpmNojUzk0H2d7bVXXz91EdqG7rYotStqCpWCNqck6jZiqZ1+riHV
JpxTM5bemgUpjlWmJclY5XLL1HiSefKjl8U7lp17JetikNOsotEJgLKBBAlEs4mwvvc1oVOmMVNJ
zzh86nkD/rIlVf4AS/miTqacxw6oqXPt6zdpX6CxLGm3KYaFNheEmGqLZVe1FH5n1In+/lEQ1UBs
pT7kRjS9ot9IlxSPl5udYrh4lUnfpKzwUizQyw7YJzYrSCK1ulQWCprBqc+J4LZmv1NyXp+0T6FF
/fT8AJ1te9bjYr5D/PTir+yhwejHekyRB1ldvIcjq6lUd6jJ/Dz5Es29QrLhwh3gaSMySaMly6+E
pHY15MS7D6e8gyUEiPRkOPKso1qYyQD4U+98kzi2QNv1AdsjAAFz4WgcJXl4YEUYMlCnz2S4TUy+
ldjaWAmyPJ/Ve11+m6pQaoSUTscxK1dAWG6cj0eS8O2wj3NWb3EFqhyzzTYTKKfIKGJbsBdEI997
5yLwg3zOspaMAqtfR7iQcEr4jH9P0L5NclwzJLsnyy7G8avOOCXuy6GS8v88y4LG0RuKMBRC+YpR
PnJbDMggW0OhrIIsMXGto+YqPc3R6tj+folWLARjfL7dgoeMKuzr3G38wynbVZp+n1Ng7/bOUaE1
+vQPacP4M5Q6/NoStNPL0ck24aflcpB4EPYF/mwecfODiIi2jnOWYBO5rm6gl7AWSKylyyEF5Gu8
9LZYwmw/pH2tTVz0FzTzkEg6qjwqyCBcfXqBahi/DjKx9s9Y5PQ+5hkmmECG8gG9d8u3RwFpgx+a
2BJ8ShSROPfyLA2/v2LENkxaLMeLVJk67hD5DoRbHMmzxoIrXflKf1+ZCbveIB87iiIpqlAAEIIw
wrlGtIwMzyb95qX4JAePlX8d4mOcuudcDKEUaLFoiOOZapubljETFIm1sXdhnsfWBFTFGHP0sb1w
xIzuOoE8au1/dCeLNfA1joGQ/OCy33dCaX3dvaHsR0JoZqi495r82ozRACeoLpwOrXTUazyAtZX+
5ld9tIxXGDTgAeMFt7z3M/7WtVkxKiny+tmFJYvQDVleI7kwSF39NXdIp2J9wQA61AQmw6vm/vsb
KN6xv5EWlRTxr1Jf1J77uGlkiAzv7iEiKjjz+On6JeTDS241Giqb57t6l4M0j7LZYdqQqUN5eQnz
28vdEQoGhJg4zLp9T/566l4RvFttP1MtJQmkVGqVKB5Nr8cmMQ2Mq7Hjl2v5iK/StHoXImblFzN1
Yo4wNA5/yqrqae1ngzBvu9TeTTgtTuMRDoFsbSfFWNWgnPn/tDyqW5a4WudkQXkd7taz6JdNIvTv
ecaeIvJp3a3THYv9u0i6NuE6nEBlqF3flxOmPqHFzIYgD8I1G50pE7fUpSxJMOS8gdq/rUeOrQzO
xfbAtYyWBd/bho0zuU8sGULVKjw/9hzQq5/2f0aMsg/rOLEj/2xe//SMBGncZllAsgOO20Q3EXeM
suxq02dhj+MBX2iJSb3l1ZMag1/EiNJPNqlSkywp50I396eRdiMrSqVm7Pt5vcbJQPJsvaqyvI0I
QOF6t1rUbdeLal7v7TpMIWVyZA0PsBVWBg5dZYoJoN04CV2C/iFd1g5s9vYcAHxm5bwoBTQn/Afe
pg/ga/bJP5B5/JhLVYxe5X5M4sAuhAYSy3eGGbcPDVrz/m6j639Ak3m5Z8wTz7Ok43O7SuLJ4AXM
7QrjUeIOz1gBHEonB1c1WocpfnbXbQe8FvSdiX9JJS7l8rkWFwOV/uDgCRZtJcOv8ePtlMpK3wyF
fHD4EBAVJGaWukGRUxCTSlrE8UAcboHSIGyOmB0o7+W8lXNVf/DJpeP93GJplIsH2bWmIDjk47Hq
SzKDL5PmOuqCWIwvm+ufbz/IXGssLcqmjmeHlDsiPROwqXx0vWx/7DfLtVmJ03KzfSx8R9EiT9qD
Ak6hDYs3iH6IJrpJilvJyyBq3qP2VjRpodNORT1pnRIwLdfheNF5Bro+Ph5aamrERulYl4s6XLQj
YhG9/yhvhmG4lg2/sjpeMwFd9wIHgnm8MH4FLZ+cP5eOtRQRaUKAmeb1BeGpg2dx4egfvytNX9du
auryn6TsqTHOsX6X7DJgLzMwDrGK+PwbU5NN7SxDqnO2O54bBD8Ec8fAkO21Nz5IUWgqKi8GW1aw
LaA4JvThvcfMdxGAlY9GEoQksD2LOsGoajIdAsXUvBZh9eoMUgP0Z8S/X7li2yxZRCsG1ZJJv2uQ
QfvJ2kyiBN8gw/XKTPStRcy3W2POX+hnR0wA+CjZKOEq6HHgKseZTog+mDFLbBILQKzqO8I72zbC
4zc3IpQlA+TvxSF6FNHFOaFcWnpcJADDghX73roGifzh55T9mB7szvjMrMsMTLI3GM8qBgzQQLDE
M+7qUuSSrbleXZo90sBqJZ3No4yay8db2eUAcJ5ONBfEAJrv82PvHcQ3jDeYG6LBJ5cfvb3wEcO/
F+p05pvLllrmDVGXrLc340d2cMZnDYxo9/uTHoVv1tN3odVZ1baDguzKTz+mybeYnhIr0B9Ljknv
dP75sw678QtC7MP1jDZ2XCtfcmoRM/BV0V5t1QrI3HOxB5eMA6+n9kkUCazLlt8fsXs6NS3JLvQO
sBXYqd1HeURi8/bO9W0r1HZQjD/LCleE676xgOm3HjUaYxu4Gz0s9KJ4DWryyIi7zLFVdUpglfiS
tX0J7qAvNE2ts6T3QSfUTZu9HKzWWVLK8xXbH7ANKJgGEFGkvO5ccL5he/Lx/UyGLu9HafjVzDed
xsDhQ6TlrRZDnj5djnD46waVAE7XRB0HbqBAt+e+UrskhpMDhAeavyQSH5fjbiWBqMEtBw27QT4z
x8T/kxJf/9O8k60zX97uESsIpmnmwzoQWUlzhC5h27794C3LaYEvrNd1m/cS2AnmIwV7zRNCZo3A
pMeEgwM8utR6ui/5pBRwCcvIjWDyAai0rDN/y3sOnln6WBCi1+NXDCpMZwyZYS6UpYyO8LoAUJl9
g2mq01dlS3lJ8gvzkccxEG/T/gzOMwJwYzHVl2FhPz9d7Svgt2v6p4aTfE1WnScGbYvRfMpIiyjd
g4oDC2Bj1nZdH9QN6coMJ01YSU2spoV2BEaTSQ1XKmjTsxPQtQO9rEXT6MSgBbzqMJPkXL3XIEUg
UeFYTvvCFu4gzwu+FeG0NiDuKkuMAZ/qlXaXsVc5VzdGIdvAt90bC0WtxCfgjxEk9QiaSpKu1zdv
qKjzrb5Wj9YgASl96kKLbk8E3HhGdHfyCar/t7hBgBJYiAKyK611DHbGLs+sNsNDZp/CTqJRPzeB
lGaakJ20quwSlO8RvWJjcBFsErzzHaY2pv2Mlz0IuQxgCAp6CgIgcheXVFwEj3xzOqb2cVuTPGpa
TjzpD4dS9KjSODQsWMhnJGmC+1DuJL+b/z9Rox1iLgcX4bRATDEos6r+RueL80NnjznASB3YJTd1
DIRgZ2sooFxRJLmQXl5DgMqnqPpCrxeYxRA4HWQ8g/8RttzKFNQFE9Ohijp38/UoJzslZ9uMAZLB
vJjVoqhq2ukWRQ8PbH2K+YOKMyOKr7V9jilqIJYAVgON8HLKXtMtcyxrquwaJVyZaojTjcmaMDDk
ap3M1NvPF2uFwQUlTRhHttqtAzokJfcrWxFzbX1pkgTs/e16jBbGGq/o3V7W4B8LOpzcuR6/x0Qg
UTYPu8NgIS9iknm3xyY9yVapAzVx0IHuzcA0CQq7axe4YOfUpDhqO/xkyGfMd65PmJfHPbLUTGxO
wKxOqwSX9Alw0ttMjn8rTSxaxiyy7O7yui0iNs1D7XZ9M7OnWRngZx1vhbdnEBoAMuXxdXLxgJ39
ZoMP1xenXgmrFPN4JZtj7Krhh5jWaOvzlPC2vj4WHAWxEr5G5uymYXgStO3EnghXhkNQp3wZHmdC
hHMdyGU1gVVB4ESQEveL00H9UuVrXL8XIRjnX49GtNrY0rl25qgk9F+LG3TURHLjhPVwko5ZD7zD
MZusHvIjLMWG2nch0V0HRLpjlwAQeu0gwOzMKSHaEzT6SVD1O4AJerqlfYlDujj4Qnk3CS+PFEEc
1rgWWM3/83cGBKDl/Va1fxAztYuuL2o8YTeeWaqd7ZTysbxbYUBh8KjDg5lR0oROTLw8cSg6C7tI
dARH8OyoZ3EftVt3W8UV3YqYDCUCEmQyjCGsNlYZviZ7HTqse/U46T+VYs10OBnkvHXEKBe7WaFo
fkqxL/dD5H9gOVg7yK0yFltnfU/yOnp81Rfu5wLChiDSxOS9bKWsN4B0U2FvDE1gJ4DUx1FTzjNN
F4OuWf8v22w1YmY0t26ue2C3oz60jHdnHqUr6uHSpRm00zLlvb3lFKJzkbXEOQVRCe2SNRfQTZpt
60KVYT1CKPPwBDVUKjChh8MzyqEeoKpsg5RQ/M9AdGuVqO5wUjUwXqiYEnNHA1gJbjWauYqIcRgw
ug2I0GetP2nvlnUCeK8un8T9VVlaiwiQGSMIUNAsMLGkOzfnDxdgHrsgD7zCzCaLR2iH8oJKDjC9
IVck0vK1lpY42xZWhLHvqE6I9kOHY2wQIC9x/Tbjc/VnwB9OJTez9OqbnK+TkIBm7lMKGBYzbaOv
P8UaAoUZAHXrRpvlfH10xIU03mkdKduWtJtYYZLdDWfOFV3P9SNj8q9ZRk+KcRaAYIdtYwOFpITc
Q5LLDIOw0yAPdo3D6FYaNGKMJPRIkvMb6MKtbJDiI7XxkVmLus4aDqlK3nbB5DeaQarL0PnOkgJ3
DsI1uBj5aIdbbqPaJhTxD3GUwAeBOJOq/0CI3OSnBPKWY39z4G4T0R949P6q9zFzapCSFRbwS02j
gbCXboA5NhA6bce848C46hSitrmW3JJVeehFkHfp7rmvovvIO4u7mWTnFEqbWd8oMT5Zsm7mo0HV
mna4fH0djYF2vSgxXHU9ztBz9wRlhR/MT3vr+r9U6AkwNA9HCZcSB38aSpuCFfTkUyg7y2stA6EM
h7ob2Jj+NpB2XUvOaZuSGV0kXUbQumJ1wIS7FiPed7ETTxFJ+w+dDJK/94AR+iGWUI2/82WYsvQn
O9A3tOfVuuVoZfy3jxhXuXZeyBSYBOdU7IqDADjI7g3wBb+2fuhLA1CBy2RoxRMEOmbNCH+iqF/9
957966ldqR0qmmmsNeRsjiEVNPhTHwhP8Rh3jgvqPECka8qqA76UfwItDo8VE86E/J+I4A8v1ICl
uMKzR4O1BDCiZHpEUJgQpUt5FvQ4n2M+ofGkAMF790GDa9JWwa4HkaUAfgAFtVkrSvP3j2Re7gAE
dk0dtqkFmo7iD2oRiLMQ6Po24wIGfA0r2722455/kIwfgnN9xjEP6Up3WtYBRdgBvu9wQh8OGyjl
j2ec12HoGglp2IhylA/j0ZZLrHZMb/HRgTXn/viJFAJ6ApkzSAc3asSj4xmqi7MPJ/I1zRgHgOu6
UluW85qZDyjvq8pCFns9U6m38JaSrs91Y69C9A9QonbRVyrlHfHnxBKvHQR6AJ3i7I7SNon01gEM
1rPWntzEoMnlf1JLuj3rj/QSezHFLxdsfPBlsQ9e+XYXVgig3JXE7QXnp1ETfytIp1UR5MUOL3CB
BwBZm5VkM2oYBkzuKLgh6fexIo4l0LXy3YthNeRpV9UvIAXnFvrEyG2FLnXF7ISIY3UDLrhR4zW1
BfG89f9RYlOsB+sgY9wt2s/w+KV3/Yum7q3rc1B0gMOUMXM0PdE5exuKTVMrgrNJR//rIlGAE0yq
dp1bp5a5DAQvSNtzHgMsIj+kzl/xGHR4yeBU+BiCxZ/0a8sM2ulI2bZyTqA+HHQJ2BBcJcO7fmWu
4cOyWW4I+Y7AVuGREpDTkRLwZHmBvojBEL3RrfNApbzL/a5sHsQjFI6zM3g36G8ka0QDLGdPvXvd
cT3fCk/8Rarw4Z0nb/K7HCejX7Z0X2wyKay7sOAIiwnPaKhYKnBDq47sXzvFhIhqDmCqg7/FMXQS
iOewPQGnX/MDRJqqhxklK8AHkw5txXsxlb3txK1dF/77UyCF4TYsnTUuasG/RATzwzV1mILQlF0g
l26T+BtXayOS2JewrVI4b0qurJu+Y09++ew3yA1W7g+DFF4kI0yYOPGEZSxNtFZhe8FsI0zblspi
PQBO2nd6Q3qzNC1vavojqzzjPK5ocT62u9hItiEYslrIT0f/PMmdbflPdG3Uu+XJiLwgo6N7M1H4
RQW4sDgvhNlAnISoS8e4Al5mEVwiWkP5Nr5s1sAM0FmX8EuwZ35E1M3bQqhZ6BS8Hg8h880CZgTT
45YYRx1fNc2o9bzwtwvkrmCEmbv4DxRaT7YeBbSAO7tnxU0fMQGhdrS2keT98VxFrio0FYxsoNiK
EoL3NXRINPxWV3Y/fEswuNdPz2S11ZNnAvPDUuJ7XyetW4fzbAoTtrcovO0SmoAJ9QotFOC2ZbHc
eRc8P5+XWVE3mnUkcWphWKxHQEvNeWzrtlFPOBed8rbWOGCL+tJd9xtD9JSBa/sqW2zIFj9VAZL2
9slFrAQ6f/1IRDN9qjeE7+3f+99BVZBrMeji0l0yZJ+OwGYyMYwi7kH4B8A2JUGvhc+VBKs1Zw4f
cdoRFPGpFMNMzhlVeh5jtQXSAVFKhJGVV+4Xfr/rgvqD1M/ouqkbsC/AehQC/uJeYq+zn0DTd5Ih
jjOkKadzlZJXENvh9lOP5VNl5hg9HXNh8if0yjxF5SJQsjnTVFNPImsjI4ZfysqJzP4LPV7UikEd
8z+RNeRywup+A9osjM5k8rR7dZe5ek9uNxH0H37DXxSaMgyzVJURqcnyrsl3sehtIBh9cNZGijAo
gU3OZb+djQZDJbkZi1l4a6wyDq8nQ/bLivG/hX7XBPg1672NpUz9A+42CiHNCND2XWsrU5dAJGVZ
s4m2idv8z/N2gMbAN6qvy/ymYdXlUq2WDGy5ytRucJe0kLrky9oaVkGTKlrrS9FgttwddGspZmPD
xBhBXNeVo7Gz7mjPyDvAbTMgFtxhb05N7msG3tinCJSLVLeYRo/NdNeUX2uLU0gBHO52/R1BLBwI
Z70FE7qnjkD6ZhF1dAX9yDEfSviSqjSSYZGYCAXF2AgfjadtAuS9homn7ZUtgkMdDC7P41wypV4u
ipQY3J+SmPmJqFwcjdSRqkQ/pi3EhZZj3AnLZ4JZw0qxH+IWlVNgBOJ4TL2KB55CSfLccs8wUW74
eG887BQx4DJ7Yhkp3D5IoedG9qshGyX4xeUWylEMZg3zXLvPFOtT9JrprZ0xmDAlzDCimP9+U6n6
VUNl4XR3+6I3yZN/jkUfXy5bEjdiqEbraUkC2hhVJRE5LTjUHv+pUyW4tOvU26wqA8XEFx0qcRvH
BGX3j/ogHe2md+CnWB60nZu2P8eo1NV3mDrfj3tcQNppG6CVbfkTWyZP9XWbwCmb6ywev1S8uulr
lkibnb1FXv3BADmcWuerBddscaaFxguS9ogM6IWC88yQmSQRC239YyOxiW458kyRW05Ga8ldDFpj
faAFqbfsQWIng1TmRnMZOsxw9LmMidoN7Rw9x+FYrtZmshB9QxqcCa55WT5nD4qSnqopGsivOMDT
TyfP3wfpbX/WDrUWc480ijZZsPfDavMiSOiLc0DklTbDEJnj5WumBjFbmfEZP0+xUGTn3CO1EXiq
Hxgy7oezdZPZfS9K3kAUVCwF1cJX1WfqoNQes9DMI+QFV+p3bfD5KaZSWBXrE9PShEFBT5p3Unba
lZm39GENLXZkFxpcRLhv0UKB7vzaxImPk5nr/lTDROwZwtwlamXZqIWxG5a8nzKh47gw+5CkJ+37
0YsU5wWqDBddh6pBpeaLsY/fhhaFrm2B50CchAiEPX1C1amsB2bya8rh13IYL3kWk4oPLt3W3hlO
UChEWu4Duq0P/wAZLCgLEfy8qtsJ3yxOJJP6dw28M7hCD3/I9+n79cwZL3CMhvqjAPVkl1owYZQm
nuNeZzewBHzsff10glvKrp0dnsVnMTA00MKHw11h/ZE9MocoqQgKatnWYwUqPqSafaVK0oI/GsTk
6eX/o7ql7QWPsebCpL81zM5M0p4fN5ZjX6rLOfRr+Q8eh2d7ic/+nTTPhhEVwDOLULx4lCUgipDC
wYHbwaaA19RFtk5IyuVByBH8M2R7aIgHw3++nMPaS+776YSPDDoy3jN80MD0PXxkQ1BqI1GvrRky
Li4AN4nwqcI3brWL+gX2XnCSKKMC23C8lzpFFj0uuaN2XR8BlMeOjJQw0vaGrYw98GvcgNudR1cK
LyD9cAHfHHBI4tMzTWbpXfZGjSdAkv+ltCG3X18LuJ2F8UGUi8SQ4jXc1JjGoBZFFZm6cd+3+Owa
F0lfOrCNmrVUzkCndDCd0jFvQ4JVnALu1saDwzbn/MSUP+OlOhocCE0AUV3DyE/jLlo5G5t5slIO
4swV+fFNqmBjY28QJHx2fprFsd3qJywsNzGmWPSKtZrnwf+WmxnsKGbcNGrKcjaiMaHchrmdpQpu
pI9jzn3O+5z3emK8oE71W0/5+lAn+v26KXTih6USMbQGIKBMYzGfWL5Xj3kffIyFx6MW4dxmS+vy
JUOq4UYHvxrmWVjO9Tl2BNDKnfW95iucDSy9WU+oUvdpQaTyXkqAh2lJ0iaJkNT7hLxta9ATmgyZ
l/aSVxxhWGq6CJT8lljyOJeR0HmN0hnhRYoNHwrxrWUWdUYwq/2cPUH8yEgwyHNoDNLEdkx1828K
d7kAdxEumqFH+FZrgmnikgD5e/R4YoKg1RYmgH9ljD2DVAV8WJ2uPql1L2G3Gv+wUg9ybv3Enx7L
/Kj0zlMs+FdOTytGpaYklNcjLhE2XQnnqtoZaK1tKy3+Yvx4luTWjFSR2OKgjVoTedMYkHg7GWV1
94+yABt3Ah+KjH/3IaB+oRMCGKC4+lLnuAzhiN+eZdJjID4PYON7jUfw9ND22w68VGUFKmtvjmFH
8BDzWK6ogVcbllLsvRLiQk6MbLNt7Wql7Q2iIDumT/zfRmnr9KIiwWfxNdSbWi4Ny6343weheO1h
nDw3QKkYWv5oyjrZHAfq5PKqNjXI+A9NaZRsi9KdKqlVkBAQirzLUNCzTiaT9zlhyxChwlIalaP6
6SLyn52bB+EYn56uWXGXOcfDzxaVcdRjEp2zarixGuBegAVVkNHY5UdgWFQ5BWEcsw9zufThNzof
7Ri7KEoABBD4qYJ1aOEJvDItQU/qu5Awu+Xsyy0tm8Ce5thsjF+2W20jtaCL9nPznQ2oO91eM/w6
4qr6LoBdQXGIqZrF7D0kPYHfcliWV5fvrakQ7tHD8PHhtGHSDIWCmjrLWAFeu3jCTfEld+bHl0gt
rVKjX4A48AUO43y34mJyKSrROs52E4+HxHpJCbzSkcXefyOoE5cWS1Oo4b0RhJ8wCXcTd/PGXFNn
PFzb5eP0rOglQjQiAUSijOT/WUnCvr1Bc4gebtl7KfKVSFTaaqDAOXUy3X41tw5rkdbT8FqXiSpG
+994HG7iPsrymUzqHwE4dzoeo53ihoTUtlmZc8bQG4ULDDSFS1exrdxznoowupeBhHuyrikFedQx
VS0/5+w4/UiuJK0a/3l6FmGUctccEKJ6p9I8WDwlVLznymp/rwsvQeYYo0YEcWR6Hgubw+uPgRUS
7v1nYrryPLdAwSp7blbrWTPUnq4T8dyV361TU+05iTJfx799edptnHvUdyOAeXJR8NnqEE6IrUCp
umHC5j5zqfCAWuFypze7Yrx0fN8Ra85XUG3Q0aThE4KzARtgG0oa1YjpIE7WilzmMWaGWYtm9cky
l2bRQ1Z15kpxD+5pd4shasWuV3I5Ryuo7HOEDgvXpYzv7FBVkAEJWt3xn+HUb1adu5DL67Dxb0Qf
gc2Vs/h83ShL9f2OcdWubvBcR9+/tPP5cdfL2VRfVPtg2VhBP3QBrCmnXkopW/NLQQ/cgmpaPHIO
P94SImEKNubhIl4rmjhnAcR7vY0Lh4adRtOPv7dwB7zHLbp4h9KMIkzY3uVJohlBohrb81/XVLiI
sxmXU34w7Sf19Bnc1F4FwyTsiqKj/Jf/aP06KY3VNU0Nw+UTI1+5yXIMMwbJMR0HGIQI2sYfBj8r
UHH7Z2+vm8t8iqsqu70B7dR47s5h//cz6lAd+yRNeqmsLN+0Hp/9CeImrRalllHeQ6FNqTa8QfzR
Uv86mMYVr8yhdDmEMyaNf5ILPHpJc/41EyGfH+k3/9ldtviU3CvvoA0V2qBKyZIdrj31kcPqUJAV
tCs87mKI8wnm7eYiu00I3hCvCgqL+D8rhMifu6vjlRdH6kXnm1KYZ/MQIcL7ogbmrwyGLDLI6UOg
Dw65yPZk7x4djM5fDjUZS8OkWkKICZR0wX49Bm7sF0gAxHhbWlGRHJiQ4YOLsIAKUiTCpJLPnqJk
8am7K8XPv/HhzvLBZP1Edxua81DeoZG4St0snOGzXUXMuaG5NfjvWefhLf26VXgLzs2loY2E5qsH
F8CLFu6QWQpgvXcjMzuLdkuSHMCoXAYCmtf4BJ1+JzkbX1t7SbnW/yE3laI32j4Y48uSd5wjz/V8
AHbcr+GQIOYxGzf/KTJ8iOWG0Fn73HEGQQFtQNrUroAZoQ/hWVctrp42ni/uu8WanlxPcYWEcxIS
N+gtZ9mRJ+68Jah9Fza79Q207qUzRbTno0QqlzRGfsVlL+nbPORlLzV5lMgQdHWUglQVSJEuk8Pd
u3mvqs6cz0UpLigwg7p2cv501D1Y7ZlU4hvqsMiLy616eYODiKBJfkYfU1slZ+2ahCETpw1Ygi4G
2meAQvqgOfXGFgWa3kXMKV9rDvG6QAKiKDwyR0PPx+gy8iTXGqb+Fzzyp5phHgQfz8QeaQEy/909
yaJn0c71o2cOBXWLu9Qymdbnq7h6MxVJv92uTRwoKUByFelnytLuwoM6DO3GhpONw/smVp/KQXU3
JAeXPuVTQ9ayc+JSXdsnmuyx35S2A27LbRXgtGwHOXe/19+pCKqzhop3UveZUTfaUGUmNlQImofi
G/rIokjn1aCRBuZANnE0qniGrQFB71Xl47YxH4IPUtaeg2gtMAra+vINd+P4nb/mzo9qmDQAyvHS
0t1H0FheQThUaRC80mLdCsfOnstVAxo78gLjK94SMu5yew5P7YVSh9cl+YdZU0ByxypCXAAV8DvN
Ze2Fzq7i+JyAHB7AWiyHUhNV7YtQ+f31xRXjJ4l7mKHX/W0n1VFkf01EGaaxMvwn3sz2d7FFNFlS
uvDZ1x79khzPe6EptJOJJjk4hihb1NWidrJeNvZeNluZYiyFPVGkqdWG65V9yMbVIcvCPSlMEx99
ehkcGbYRAgKhEmbJU79lXs+9Fdb6U7IJUkK1IEEpN8odfEbnAwNMb4rxj6thFWwfPFR7cDdjeiS0
cisxriMFiCs0DgEZadSk6Yp0oyHK4lOhlfEE1nYKxYiKJ01HI//3kKm6NSMMaLy1xdGWsPv7Iy2h
RpQvSBpdGpE5/Iwtg9ue5HvbhY3vfOJI5lrWSxWSrQihpmgql5ostWA2y4yafNkMlsea7NVkA0z6
D61sEr06c6dPzXjXm5gj9dPDeXEMuuJ6PKD+JCbU304h7sE5pc8o3eC6tp+AQxR71327kJg46xp9
ZQ1J8D6sBE9gSDhp4T/VoG1gdK9gKXc7gQgoP5BEPB3UuNRvcxmsIrWUA/Z+M6zKYqld+z/2gg8/
t7cdHK5pZszCMPsO9ZrVaSbIVZ77G3tRBohsTNGYwM+6E7Lf5xMt4WkU8GSevD1trSaSV5U40FD6
z3CIg7q7l3FZLP+VGZDkbdKY+2zR0S7EOR5ZRYoj4KWEg5FDZrHOAPLXuB6Br275600HDw85fQz/
9Fdgs4Zw9wxKI93i484XLj/bLKvik70X2nZFEhWVeC+2/+RWZ2ag0Z4xB4SOxplBgnmFK0Glblrd
PIr+Asx5IGjybn15fWUt8+Z12QPbLnSjea8Yj7mKkyqolU0PuxbKuKB3gQkv6MgVwItndi+SwQo8
o1oH8zWibQtWn4hFbvVRrP13m1mG9CVSCKIgHd6hOwpm3XB8ulemhsPQHZOW0gFig22+6RBrbbkm
gnkFci0wX+bEGDdX/8xXQWAUrfNZ0Ktk1vNyLJKfM0hmZAjba1uHk0ywPQZ6HwYM3VYxF5UQypIs
WL+39K091+cTOz2GoXTpUqfmKniCtQDMdXTkYfdAukNA91zRGFDBYVkaHMtaCbBA5EjxLY5qTFDO
JVtvQh67PDY1Q2Q/ax6ln406WW7XzLQSX4XhMHZkXxtpM/WZqPTpqwW4imV3PuZR4LLUgDZH/Lnv
8/eV3mmp+cRHnO/g5FWcKx8s4SS0fmlJ6r4yV7cWi9RLHPRZR+O2Au+3Fqq0flUGh4WVqS2wFX0W
EdtAO0f7mIELEDRPgK5b6G6BegkO9G7q3jIRr7ZUg9nb43fdvu8TqAuhWc3U1VIuC0kJe6cG657A
JMM62m68GLd43LkboU1h40hUReSyq38i4lXJXydqlGJxz0HEp2QZeVmCQhnJELoDVzE+rZGWzm9c
Sw+cFRvnyN0nHu+VY+d5Pnc1z7nIhKvZlQcZASLT6ZU2M3mFAZtgz4ip8e1H5mCrmzqODh/chnNA
9vd7GadIQDTWpJA2kchTORmVdY8rtC65a42K0eJK4Jdj70epnPTvflEAjtcs3apJ1walz2bVNNNt
aOUfM0co8C4UZVdrtkgKGAjdoi5hmhw/2xZEnp0ODwM/gl59po+giif9rO+jE/bOPTv41CD2zVTN
5ov8O7WZc1Dw3zDUu3nWG5g0WJF/YiFCX3Zc79uMYS9p8DjFSWLDB0WmJICRBG8zkWXmgjKFqXXq
mUWUD2P+5aTP70SYKKUfNO8UrhRVySFwtizFYNMZ5Tk/0yGqOobziNkgaknJg1IU2uv1cO2kACj7
x+cMuf2UH9YJVrtxVUogWv2ZwWbfjjFnG5c9zFw59gVXoxL4Xyq1E0R1byDArXAi1rT/QYqYAVUe
xiF4viEeWStRj4BObpHvLg9hZn+lUFVmkKJ1VU/F7qLbIyjtst2naMvyjm3/3j4tVFarCdDqPdct
LYAz39dZmT9XFMvavK0zCoOdPu+yFWGJabYwC8vmU2Ue9MDLak5xB3S8J7GDv+tYrDarpoNPXenx
KlfgGHTPJZqDHrb/MZm286Cxpslx19c0qcX1Y6VStXIYE3yoXma+QiPyeVzrhtsMglmIFiso32wF
lb3ZNhqx4gL73Zvb5oujuAJlJeUJ18nTlVz6dsoC8G4Fpr2zla3C+cC5snls3nM9Xe79wLEEgmCe
G8P0p/7UlvrIIXBfc5fcKEAcQTzVf/a+S+ObfduVH1pdvu1byuh4FjaBKngqTsaumKz77avMbSk4
uiZXkkJz0en5+5sQ3XGKsUqUSx+QI2xcTbAAdyB3sXIrMghTIwVvbWYS7flyy4UnYKtAYb7UQvE7
JP2FavSePfSvCJn3HbBoFnIHP97F8qVK+dCuZSjEA6ClfQREuEB3NWxr5b/eMFgU5ILBwvTmI1gi
FdJGiKXwEiovISHLOXqn5zxIwFkS/8bkirwRPIwpNTI35Z4JbhD/s2bZrCEPc5uXPowPlnBX8adF
+TsxB2HvPDskkjL7ScAmuM+fxmWmbMv8ZIxS3uyxIFJXqwuRy5fPnHBswi3RRAUNVFuiLNqOfuXY
M/nsPXXRWE5JsWhKTQED2LgeOCz/jqA9UVIBPWZbZ6E452DCPNlKetYHss6zbDDrQJmHF/NFQytf
iNsXXbjc5vj0qpXg9ErGZ0AUgu2tiwPkiEb/QjG8ptayLNROS9q4piCyOyikzhn0u2raKBRpFCUS
n27NXSSiD+V8edC3xzCKTxDwhMFKxLJtAFUbGLtZ5tBG6Q9DDfpPHo2tiRMO4cwMJrXwpmZz5mAd
pPWWkfMfmGPMz/JICI1hr3mqXH3KWNKZuc8jivESXea37NeA/GohmX4WUXA0XHvlIKv8B/yX87oq
yKiF6LXkITMHBmduJwC5dm/9up21eAVwjNgWQyrH+r7vLhFrdZiPqekC3vE+pRTDfgsnCD4fEGZF
O4mY0n+XJRvq0D3x2RrcFQdOcan49Gbpy/z4UN2Avvkbvb/0dW12TRcOx8UJWrNJViR01iWRmahd
iJjK5BFsU83OT+9Oz7O5zG1nDboSabQaFJogRyRKptHQ6nlWSGx1wE/7o6nqJXrS6WDudkDaXRQx
zOUqZyZdO1FutuaApf0k4Etxe+MjaHWKPiJI9vRyujv7vuLgPGSlgcfHN3u7d/Ke1vFbutba+1kH
ZLqIsFTBerNfNaljU+yqILs3xdrXwFYHk0ZqK+aYn8G6h5KCnodalzzsEuXmEVyGPaOVDUosYeY2
hLf9HlMg4cva/MQdkZVfhULM1XlY8QVcvxv5ppWG/7ao14mAbwYBHJItd09+YJ8I+SsM3T3xRDu6
84ehG+L9eohMSuPFlqVYNYX0aZJurdlsc5NzGb45lJX+JlHDJwfj1mVPx2wfCnBbj13AAcVQhGPl
1VMRAFMOLe3oqd3VHlJh9InrJsJjE2eD/5cwRB0xNCjmHzMgd4FK/8Mi/wkYdJEAK33cEjgpHNEa
+OeO+kiPWTvsGudJ0ovc7tYqzCbap/DfomZy/Z1+j6MsMHuqLvp94jy8CX9DsoBmcMxRZO3nLRyH
E8VEzK/icnyrbvFKjEGmedm0tJjCJlXjnB7sz/UzqmAJDW1lffhANZUtHw4+rjNrceg3nLbeUkaz
WHN6RGCXURw5L4kcI+k1Hh9mKFtfMlI0ZBUyN37MUj7aKTdV16u5N/FTqQ8VMG9ZTZM0jITugaOK
/B3zqfpDXxDM7cPXHQESOL3443EN4E7OekKp2zv7/Gp6ACHR/h9SfWTD5wUR+7eBZnhJRcf9ZarU
lc8Gqky626iSxlBSPsJwsiXxywbVScz0L5IKHZHY1bjILM06tMYzDjWLyERL9++odmgbn+j7HXgI
Zpj9xZcAC8E91O/N+xHfm3TYyWoheoo38dtEG45O3aeMqR9/7vKWuHU7ife8D9tbkZT3vJ5Cqk63
SyGhRtwMaIZ7Ui0m5cNm6Y3XYMCqZqqIrKZj9tx5zkpsVrjCX7Pb02tKqcu37mUEM30m2L/W9mOd
eo2R0hHMpnwrmyG+G24Ub2DSakyVOEzoG80ms6fDBrx2PGTRg3zxx4Ue+DhE7As1JkA+Z2i1L78y
ydQrcIA42InYoWmRhlwhpkdXhb54HaYLuEfX/7r7zo3tSGL6yObHtoEXrDNoe87GZnWLjIICUw/s
UeIoBmydTD0czCkVkraa66jhwQqw82Yt1W+BHqz9/pg7MUQwgcHO7EydNUedSmp34vogZOnOScKh
kDDJ4aa/sIFifdofMElI9kL7/qZRS6XPvtVTt3pqeP4v3xErLoRO/yaSgCwlhekO9J/zf2CkTUYm
cHCsiMboVmHYgZp9XcbHuO2TmttN7zmSelBO4XPP7GETc4rSeaQNh5j32brZW6A9Qsr7pBX09x4N
fqvd4WIDg8kK/XmZ7ZvJF+n8DZae25G1iUVMrXP+CjBUaJADLjs4T95dD6SvGoKyYZJ1tbz+zPkP
dJkY2jNJQN5iJra0SAc2sog7QuPh9frRr0iMU7UqeHvkHoBmV1giDCNyK9LKDQePI/Oj62zRklay
onUThGWaKLG2iUDGSU7VPGF9Y+fKsKP1MZOpUsn6DYKuQA+5vF6KraWneAbi48JLEv76FGrG2mNu
iYL0bJ+OGDv/woHKHWV80cr7aecBVox3GJrbMeAFIkH3E3SbC12dGIAIS4qHdzjCZ6cr8erJ0b71
erXyRr8m8NqHmwlwqiN7lTaAbeCwp2UkdMv/apZn2u7254Nssv0bFKJvt92OQocwg8SHewWqDd2T
n8AUIVjRCB5qmY4zmrkMPcGkYPkoVhcmOaxZJI04EzqJqD4251ujZQvAiuTcJ/s/w5VUN9RCv3GW
r+nXUKh/BrftaE1HXlMZwPerb2wN1HyOhYYQoiJsEAKT88mlCrscmIA4nd+iRlCCuTQAghADzJul
H9ZlVDWXzEfheMjhm3RpCHCmElaoX9H/VvR9OsWuSj9NRlbCR8r6rVdjYK6qEm3rydJm4XTWjnT5
LwDzCT6VOYH/h8CibIvnn/ZB7oTl4L9s20inEbsdTXC2+GZ801//RXCFnvNSY4latDMcDywM2PGS
3xt4xE6QBe3cCdsXbxxAB3U07cJ5L0/TBlKAfiDbNwGo3ter582t12b+NSnmQsYGhmX5moNrTwqn
vNUgWlfJ438a9o/HQQH/u/M3Uga1sSgztgMmyC7vSBPggBQYrU+XV3iYpQiX9fCWccqaYDPSB+mS
JkjAZEfx1xs9xp/QxSZoOC9ojWCv9PqaY/CXXDJBWi6nyMkgXJfOG4vYHB46g04MyO71FbaylCO3
uUTr9TumP662+xw+4TktYKJq66fUXI+v3SH/mpoAPIAO3TyiOm90lY7duwJ44VBDW4hY28HGZES1
5VdWn9oHUdZgCRzqCaAYeHtae1g5KSlaMwDBdOcePFkeckWZ61zIboRQUwAyi7v1U04U+B8LnzuK
loFojTEYcYJ5pLnKyDsQcWIJpT/AiqNgvOZrXqWirfU6GVCk9J5XZ0FzeTJ9EqL1gV/JTvrb/uIf
ZgRs2vBOjfn7HKKkpQ2yIlvGphPRqrAAiR30gXcooxSLELWUuLAYgL9eBU+/XI5taa2+90YK4h6w
1vuCAqvdOQbcBNh30z51gLHeV0EettaSLK9ZgYLSLv3loy1+OZgNUB67n47ELRIq/5H/Ixj96USt
9e9CWhMNIOfTZH4SXNapAdXBOcDKPEO9p/5zQJezhDbKUjxOEScioRe2BM+nazfq4NiTb/Aoner7
Be/mV01n0xSevNldJSvIkAGx7EYcV1wpA1zQOYh/fGJL4XToZOghLg2VcSGLxNzhyEhFUfV39uRX
tl+g3y288EnG4hscj0s1lVNuHuxklEQffkQir2Jhru6Sxl2bo5f6EetjUvta/dHL/qJ+DkDtbMbf
Tbon5Edzhc/2RfbFSA+P3CQ126mLKDN8/gR4Y4UWNRjR7IGGAA/QGLwEvc7px95kZ+f9MHTyR/hm
9SvHIhJsXh5za+ZpCfV3cNGiMClhuhh/gSpXdc5HNg44+/u6hixZrxGYOZdHnoHwF89ow8+HHFKg
lnWewz2HCDrwNb3ydG7Rc8ZJnogNSSEKky242GxY/zMFUfUPsv5exNoMioElA4C+fYGu2pDcR0/u
gS8vNFLTryy3Cgo+6LWpShLS3sMNyRZbhf5ox87+E3aqsU69WPNW/kfTKSt4ZDvA4ywIrSGPNim8
8UMaE+5uPDkzLo4EVBkA7xyqYfd7nGK6RzuantKxFt29e53DnoAIYHwNqJbN8FqFHPGNrbWUrtTm
/Aw8toX+0NuHCud3Oesb7IQcjmUSI15BkbkrOiFnga0yk8MjSl4YoDq3eErcbUUxHpljo5HZI5X/
o9D8rkKF8bpV1L2FyvEX2foLUv7nqzcZCxItVwThFpdVIVmcKViOxygEpyA6EH69BRNGz7MQdRF7
QXrZRsodVZr3ukMcumui8PMXShDT3H57Ppf/XYscXUrghqwJhGDMAbvNX2JnYCbrAAbJNLnn4Bjs
Rr67q0qJqkBIR+ydqoGXe8vSH7sqy1l1pR1ztRGzg8jmHH+TCsPCd01QV+kuN6VF81rPYXtVF54G
lbX9S8f3ct9J6dn5zb+oWmTavt6H140ngEqS0mDtDEseCcjPwuaeKlDhlAvyxcRmIpowxiBx2azJ
ZJTyIFAN8dsupJxud/2FU6tTW4fVwefPOjeuqmYK5DMQLUDD+DNBfABPVIqKyphBGXFZpmiaMFip
x9KF9U4/4UWrUaUEacuNzMqBF/3v3TIJ0QV6wAhmfvBa/WlFeYo9Jkknuqafp55Gp0Yjk76HjVti
Qpp2g/qz2eJW9APAPgT7WmWipXMxNHCu6Os92WoZxnvXXDaGYij+L9TF/qAhXfTIYRzdt805L5s6
/iCTbPrXL4BPZA4Kyw1ZV8BR8KVZ4zsbNXN1N9IZCVzpqOWKTyyn62mqz/RRN1zz0ijhZn5P+OOv
J0LQ6gBowqbCJf5c94jfuGgsUOkgJkoCMKCef3C6nwSXOAyzfF9PQGDZxI9t/Eqyw3u/s0C9BOkA
846pf5csUtw7yeGlcc350BcWdxaowKkgtrH5Eb/HBTfU3Xm3rDWsLvZY73+iiNaK8qV2Z/aEaULs
Hap6cVSINfc5Jn8dssnBD2ldEVNx3Kwic2KPNepWl4uXohpBRgB5pK3/x+U8o42y08QCaCrhrlKT
66iHsa3ZWIH7XWk/tkG+soXNowXmQd36Phko1PpZnfP3AXVkz+4OJ9BvIe8y/mSdaXx4QRfeM/VU
Y4vL6ReIpGwrP1/A6Y00Qz++qBx2C0dS0KKvHsvO+aLnPI8fQAzMHlZUod7YpB/VKuuUi/z+ktM5
Bposp9d5c1B8YUZTWzsV4A5i4DR4BF4UqgJjb+CFJB4D3eLBFy3LqgbV/JCvuILV/NSmEv8StXzP
YEH6GwYMiupgBkLqR32NRSmVgLDijhHbg8t/a90prUUzreAw8A5+ecIV1SGnUm3Ramo+iXKgYWZa
BnxxvmPEonfdbrj5E+rPIv0u5+kZHTKVpaIZ52oecyPtogWqJlFG7ma6S/UUVXuVd9n0pn4cw49p
ldeMD9q9Azc0SdrLgYJNy40imm/+xyrEJK7EwwWVgDqXB1kSuqRBMggfjFNNQTgVdSBmIVL4Qe7W
+RjVAtoZ1NZMZzk7ikhSGrcwes8B7KMc4k1TajqlM7XnJR0prTBGxChz2iakx2r6kb9ZHn4a7L7m
DfJoMI2KMkaRir1fQ8Y8Oo37Q3l1hFOfTlxvQy00mAtDlQyENhnojfVubL8iizgkgRhr1/z74oBF
yCx5C4NPbBMQTsLn072Kyz4YDwd60KVl63TF9COvoax9+p32+4JL1ZjnEmhEmZQH131EXVrHeUyK
mtRgv1Yc+nSsl4O2nSkboLxDA8jXQpQOqcp2tu6G7x/pfXlIYjzEPmVqKdXT0D8vPl4ZbHX8pk8j
AZbVi3uKqjEZwDMSg3n18Mrj88hcQa5Q9NIqql2wm5i90rTZIV/TxE3OxCWcXxgaeADy8IpVXlhZ
ZWSBBxT85uwjgV2xm8mZwDqUCHd46/z6pbfcIAYkmdxthM81ahCVbz8hPnSr1o5MrKCvh84pKxYL
Biiq165YCrjDt9kShCglVO+6yKueMVAfNyJWGDK2vISIT1BuAQcby6h1eP9LYP1wKKk1UqVShEpZ
ThWWqsiR/9pDCqEHSwEW/XdNHQGUSyNKcBzT9FHhndcM70KcWdncktIcj5BnpS5N5d7arb9WtRGV
2D5BVEizSyOnPXbAwyR4SSHxgIEyLAXDQPkq0VpNSKFCygv1pQIgWdanJVxIAw8VTz/cxUuAKIaq
xfzGaHaBqIoul/CKWENb2r4w/+tPqb5OCTcX8K2NcMXiLf7PBOc8vPy9xLpHXVJRPPiMXQWGPBPH
QU2/BCo8RWyJjvPDkG/esgq0yl5Yk9eV8y3mqP706/BmX2on3SAD77p938CJSA+LMIdXpBuBxHGn
ph3nbgb4KjEDOGT8Dje4nZiJ40TGcj/8DKLLZGy5tJ4cRovJHtGUEcafU5m/7gK3Vp/bFibCyxLa
Sp7/OmWkcexAMBWxpLgAUnTw+2P7MNcgXlDAuwmUYHwKViel/1NdQ0jYhsUkz5VxvPdAdNXNdNMl
yVFy7IUlM+8Yi80OF39RK1mzhrIlcF0szbcngrlKkgL1vv3JoPeW8Fhoi03/s2ipXDRGSsbc9Wbq
FxRn5rc8Ka8kW8sHxYegEp7JJpiIV5p+Lo6PruGvl/l2tJjqoC3hc71hXDIAU1aPWDH0IR4qlgIR
2hskXCpxUrydYGwAuDf7lNSDkLBDp1rE3lt+9yde2mko6iwtB062VHPc5Nl6XCbaH05+xaA3ySMn
zJDGxhHwZKXr7uTcAlN6LWBUv2K6F/oqBQ3uFO/3wf5bqxXGmLH49PI7s1Z7lm9xikJRq0uR1dr6
skY6LQTFTD1NzzkY556TOgJ456WulVDx739KCgrnFobDOcxXQtd7VT7BKSESFGkQoJA6QeqlZmEQ
SjERJeQF3C6FlQ11RR9X+KU3aYU8g8I/AKbyf8uaL1LUDyYw+X/ll/oq76m7YFX3Vb6t8xwMvVXR
JYh0t38Dt1nDeff1FwZr5dCBVjAqcnjuLqQRt+LZk84l6HA2iQB862hw3cmEhyPejfO5eqJJ/uVq
oXUwEe/TK5Fr1OFzvHYVP/aXNR8bKhJ3G7Ap9i6m/zEu/HOmQcdLK5n4jnG0MiTLuof5gBWiXvVx
muAAWEHwIlKqxYCBTb6dezu8Rpiau1UJz02pKjbmbEcVSj1k4jwNklnQelO2TB9n5FX5amZeH8XS
/+C93lU1k5T/urODHGzCfNOr7daCB013GJwM24ir4JqyEySUY6/AEP9sivz1wr6dgU4yPspTjw3+
p2F7WFHb1o2uFjSb8/Wu0O6ufOyINHFvj7StfY0dzjcmKB8iB6qBTQtWn6SCcUXOyx5nHyukiobM
YAr1AV87WZrgqetpblGg9J+Plc5UQv/fLfhxlYgnqKtKtYltrIR5vkdYQyMUAOGF4szpFpxVcX4n
6uTcMBuaJznH3F1g/buubg9OJ3QOufNIYcAuoXh31CtHrWS3SVhiSh3qcHixk7uhXkt8zjaP1xBc
Mc0UJ+A6pF0sKvc9m0+VmmgJV9psETHI5yilPXJEytZ1dVd+OatSdCyiu/cQfyfVobYMDla7uuPk
Z71u4kh4Xk2miRUaHtZZgPRax20k/klwF/5X7EPByMoUaCHqTuTZ0vaF4YoBV9maerEnTQ4y2Wle
WO0sHPKj+y6AwHrbTa/oXpwptlLTwIJkXtmpnH4ZurVAZMp5Uul9TO3VMCpJEmdkOj0sTMPTeU/O
eMmf3Pc2kmsMCYmEPRpTyoNDe5GopLu0lJDyVY/dFgs+OI0fMcrQx5vf7J3HEcf2MyurOaFn+RCX
rCVzzQMrkpifBr3mmSn5aHaHyWrrJ+UDpoOlggWab8JPmszLllvzjl9i4tZhaANztK2A2p39n0yK
+kZZLUzM67HJ03cmF2gJ9CleUHebF6SXGniz6QliMgl3+Z0DAFFndH+PDxYP+px2hm49haQoOUJ8
6BLYRfw8hKVIFmaZxqx93P7v7Ya3XRgzjDWu9/lD9CfRejAcTQ9bZl/78wVeuNwlZ13dSXGDg0ll
gw9GQ2wgpZIV3x1jbr7UpBPTTm0j24aRsJEFX8Bc8V3PkiDas1czvVtamT+kWm9i+k/oy57RyDVi
3RdeUEXNJ1GaJeehSYS0MBLb0632DpY/ywzkO6OytCsL+mOxKKY+XV0myKqzaq9T6YcPKWY9MvqO
Twqx/jguCGxDhZ7Le9ZQ5GUuaGF004CjIjYLwWakL/tBhXopifht8UyZJn/cJcPPa3nUKiPzdUg6
h3GXrisdrgzsw8tqTRbMN78R+N132MLGVXjVFy7tBUAdKdLBex1IUOldn36pKkuuKH2vx2a6pAz8
8O2KSB4CW2cCgfDLyNj/meTxWzMB9wCLtr/iOO8lGuxlmDTaz8zSd7hDJfQDQgVjZJjnHTQTCQL4
2+gcfXHICTC7lNn+ClEbAef7kjwxEBHPV5rRbT0mnJWy5ka9YCpPDnWyqHYLvX1L1Sp72RuK4thY
OU2tI1eIpbpKrLlMnXeIdoK2AD8O2+51/+7eGONPq9ojC6LbZDJKqSzg3Qqzi5B0El+6ndH450Mi
NgVmXVIK44SGN85rAwsm8bM3xq7ZXO+wkHGygAgng0GZ5I5W3Gq7674onw/zH0RP75SAkFFXn5AF
iaeFRIob/niNXeyrd+dY1np2ZwO0Z2xZUHy5XPM6q2EiNOrwvfzjnj/bRev2bROaYqPozisqRFgv
7DtfvL54XtjYUxbDKoTb5DTihGEU58R1LL3g6TpSk4XL21qwbrO0VWy07/ulbmWWif845LXokh6P
dLIk/MinP8yU4RNxgLXHOIsCKUEK/A44e0JN11cH++xa2aDWrD1HMM1xCSCab1cNqA0hPoN13oAj
LmV4L7ivXTa8DoZY6L5LNcLSTp8+1uA9Ec2DSqSqEL/o5zVUHnT/syH8Kk4i5EaeolKYK5pA0VV4
xPxD7sykFPh1bctiIBiUo77IfET1c1xRnSsSi2tphljLDHJpxEECh7oNySSM36643v4I34IJgrel
/fEbklM7knAEeIEz0jJAtbEp/WrlKVl/8PZTHCsJogSVMBI633bJAnua4RCdrPvXH2yMNFCylARL
9CDZNEEqg/+hVILBpwP1sZBALDvBeK+WKhaNB4JD8/j71JTxaEkvmhvRk/QkHIV9sqQIEHn+p0oy
7Xb/Ah3p2PlsOwasHQ1y7pJoxnA6PhbEeiUNl54/q8i492FQeH5tuD7OFjjzuavKmZCuwu8fZL+N
1XEENmGADQA2Dx6SGtr5/9kzuEHLAFFmLdC+azAh8mhmFyQykralLmXg2h23jHszvEFCT9YGK54S
C1wIUIhA99uRHP7NDjyLGqLSyIDK2/BGvBoU+FtYXbCkWonv8t3TSo3jOpJ2DTg0uOijqrwx9Ndq
CoObOLEu2XLJpuDq3NUzoaMZn35AGmGwPyr57agdFlw0BovP6vbjHOit15emtDQjAyRHGRmBZH1O
XWAAt0a7GKfKY+f3GqNp+X9D2dWib1TPyxLwMet8tXpXSrLU/OFyiWj54tb+oHApGF09vZfsV6Np
K4N57McjWnf4wXUEIdOiB1hBxbn8vkio/N1xYd2vCYbmiCglBuQjCu2l3R/7d/Ly/qOBbwl4EJXw
OKdbMv+erTXa4PznbiUsT1IfMHxosqCwlPxSj+780X5DAL5okpZtRvmak2KJD7/fpGWHySgD7crC
aEt8C8DdauRYLsYO9w+su/+Eo52+sRATXzlOnIw1PpmD5DxGLjKeyOk0aojX9bQpRvGMBWux+rJs
cn5gH3yNIGPUzWU919gCakmQKG3y1rdcs/GnHoaO6lj8oSrkspU6X2H7rggQG9TfbI33SyTuGJzX
1hUPNItOPvurP8UwNlPW5UWu0htKL9mRwbZWDSdxLZIOsB+jnIbEuyqMSBjyLu57jkqh2nd4KvLn
dA0lAmqmnvVefc8aAkqSb+sRX1h2mm4sYD3y6NobsD6eKPLO0fe4GNiOic+35PkKrTdJB6hGdjKE
D6BBVSHqdjpFp3OKhyECqsh8Z93RNtPundOuo8gXCzxKMHS/BuXj1/Kcsutuso23QGhLxYeVByil
nfnz0ZHFLdDoq5k1kSi24uD6X2LnnwDrD2JX4pXgxy3cQiKJn3g4iS4SRLznnXEy3pnatyQ08jiF
NNClktKaUWyMhvi71Utjg7VxkBf1Ou5SbmhRIoDHWI25DeEIY7BelOunUcXTyRm6jF7HA/JW6A8w
QabyMCANr+muDdMVVdzhhJ6RzNcdUjnHO9swguh6JdMizkyj5y+tBoh4lmu/t6Kqo8FZ4FjALlLI
OPY+ho2bGRX1C48ZlsXX1c4fcantAFJG7qTm7LnQuuOeygUQLhPrITDH+Gfk4qdfrlDBergZUFWJ
BYMJfJ9I7TNaz3pLMjcH0NicMWzKILeFYQJp3+i0B+yA7t169WT28p9LtYg17pqRAZoxrA3pUnHY
NC6v/XBFO+d3OyMS1IWPok4l/Zixl3u+S8PpqGtNuQKQrlrJbTcyrQN33v+2tON/jZwz2ejKBILS
/tYk+ytoPiIBNMZdHPvPlKSR8OumWRf3AzXdh3sXEMKQ0RDTrRfCqjISINAGqM4esz5GbGsOfiKq
UT8DdwbkoZsVdr53dv+uVmz0WuIHsgDMCj1gKN3fTzJwoIxPEJ59q+vL7czVptau3CRq/fu0354L
J+e2Jh6niz+Dhc62yb6VDcOQIFm0Czult77guIcX4L1LlIvEfb2OigIH78Qq4kNz2+lbdpFh43Ih
sxf9D2lNxVwwpK19eGG6+VmPPIzGYGd3s8NvO9xLGXoQQ0q3dYHMGyv955kdWA6dLJ3fI2r+17AV
N/3Pkm/sRQp05gIlJ9nOJFA6LsC3uQXolglJbTJWZYPSLh8yZVLAbhLKbjdS87LbXZ1OK5K8y6L+
eTS30f0TdwTMAqkUgU166c5WLEMRtK9S5xEvvl8dnWdS9MigHWzreyzt+bf0HcUFJS7UtJSh9G2U
VYxVAdymO6pYo+8U5j4Uqnvc3GBvmONb9yVFTEEYwbyzE79/Itqq33VWPxKRNgEHwn3RaYKPgHwn
DTCg3ROpFFmCVk8EvSYkbd37iN7AlBbQmhiviMJt58Uz0Mog2TjbQMFtXulb8jtZd1dibN5U8K/9
DBnFA6HRDMVV1avEqc9+1it003pkheHQpk5jKAq3aFzE5blkonTJJw7NH4gKcFYDPlLNLT1zxXar
MQAD058N4YTtdwifQ+cYNZppVWmysHyYrPyp6+s5Jk/oZUzRalcycLjzHvryZe0V8J3Fm0qbsokq
uRvO2GeL2LHeMvNvkgvrpF0gwLwpeyEe/+HCF4Nv//plK1NYidpZZaoeGNGZKdz0FCeL8W9386LX
bHjJEXqy/5yQqjXJZT5ktN1Dc/2dfBzo1VCus0wYG5ej09DGI/0164a2tumP9OGvdMPWjr7B4m/y
GYhiC+GcUfAErKipIoKTptJyuP1FtTgErTdD5MroR2t31W6UZsf3VtsG80q6D4q6KpbURCRtru4s
tGIoOLR6FnuINuJAtV7HLvz8jzZAVcvDhEk5I8tbET6ca38rmETXLmTtfYzT6d1iSSDYr+jAodLj
tv6aMbMLqB4xraTEP6AwPjCUqChrmGpjK4jFJ4m8lhH8ltigcB27cJvTBOq1wkU1hHuWl/g+eg4b
UAr7KcaXC9mZgouyVt+1Pz1ZCJiwHnKVcvnkegfMlZlKmTtNuCfHbdrpr50ZrL7Iuoi9HB4rQw9c
XRRu9gChpO26krd9jV6DhlB3gkn3fB1abcaC1NI/OWFZHzHu6q6Jvl26RSJmHAoyc6KZYJohFsOP
6ZVQXhYZKvz+lFymduYtrJbbSKB0nrYkDWYBWZQDSW/3BPKAxWnpSgP0du6qydIXTnMieKUOTJto
ZLGkt7fu8i0aB1B6bTgL76H8ojp9ZTr1f3vEm+IJMNrMuRsWh2jj7BXNAyFORkQ4twxEMekd6Zn+
JSBccDrAwGw7V4UaAHZX77BNwg8IyTWV0OzTmVQoYO8gOf6N1dIyuSYLhBGm9kQNHqUMfCHRepBZ
QWoh5V2HhiqhwXKVD22NLCDyGvsZetsW0iYWPe6XsYDbL4N6FfAOwzareMRUPZTg8Au5USI/UYj5
OmKO01ZxphIihD+S3MMF2hDrZhR8w4rsjkGyLrUTVhOCjgP6KsIBxheEXqfp7MXtQUFBMWzaAcsv
10aOGneTfziwzkHPJDhenduujWcX9SRFK6wPwzZsO29oqv5a/lxT5zP7blN53YmWado7bVLaP3dJ
i5ef+P9Za95yQntOHr1gFJupnzngoyn7QjE/sGGzpRKrLTOIE+Gky3gLw31lxXM0OADPHP9cHm3U
V0rp0lAyIjw9eu4wr4mloNlBUDSzDPQ4g9VmNGt0CIhGa0hivRaYnKe+4EAcO63++waRJERcLeK2
ABhjAUF2C4jDFj1xmhhb8eiPjPq8vvHG9S8yiuSTnmEagOm2x4E4XSVOW0QgzaDg3HPzcNCW3fny
jm5fT/ZoPNTYTsSSd9YbMi87F+1IwisPWKhQJe3riw2B6srseg4s01eObY2gY7vM9btrX/Twe/qH
Qzvn+XxiPoYoWKQceVKcHbhFhVVJnt4scVMIdNcpXucyK/YdPEoBR1PhdrPzuzjLoZeeS5TI0YRU
E/NJcYkg8tMpDrINcobTrqzq8CHAh6utJi3cJjFHFqBLZrFnnOUWTIJoByHQZooVhKa7/1MiDXWg
h5qaoIpXDHkUQlbY/xZ2F6Rglu8qoatjYS7AkZGEhBEOHhpPvKjMmHTBKFAXiInFhzy430vSTP/8
epBzqjWx6YIRwxSI+hI7czplIfIiovlo1XbBsACwG4RVaeHmBJ3mHwZVSlIekNNXKkNl2IFLduE/
sCH4Wty3pmo0f8GjsnxXaB3jPLa+qIjyaSSOUsg6d8WnwAVPKuhTRhDWO5sNywsFE+zVg7lYPLzm
2GoSt6iK0TFHxbSNWKkv5H5WBiH9WGhL3HuMB3WBaM+lvP+bmAnEZoeUX0MZwfWMTBwlk1pCOohp
2SSDqDUUrOA50ki1XQWyBi6Q4QpOOtTTkhnF7KlPKddUfu6onYMvm2jBqfU/SM4M+EoVwR1ItRvW
/SxzVtH7VOV06kPidNerRAACMPpiyJvgF8kOeRYB2/O6Vl1GBF6sY5o0eiY/TVHyCNRD3kwbPI74
1Au0O4i3aIS4N9GcCLviZc7lDZVhieSn8ITE627K31njuRGi3KoHb/C24YPTpd0UzNOLt98j5DVi
Bnyc8+KLOCy55lkw2MdK1USay70Y7KijeeLI3T2zpMG2ZtJs+h64CJnf5UeCObqiLpKnDoiY9Z84
k+TKCg+boRTPoPGYKs17+x+ryQbNo9+SoUjb2OaLDEYYsuV/ucftrNjxpN241aX0CnBQqxBfW2if
kqvg0KKRBGADbipezINFSA060uaYa8ptgoOZJ4t401vs25AGYisLgpDZnilOP0+30ajSZr5vv2pB
aqp/K59s5buiFUZjNQFziRWwM/gfP1VgDh7Bgm+mcR8XE8DgOp5AvmOgyjj4DXqeNmO+iKIYWbRn
Y+xfd1ir4+cmDcJC/FNtZj3v0b3so+uVc9KtSV9L3C9h+iVC6UZlfZMmMzXnIhLyAXqK+YNPcjgR
7vAz64f54v/seTOGR+g6Bgi201Nop3Yq4/IwEmJnpRG40d0RYJmF/D0TT/md9Qv/Xvdk/KqqT9tE
T9uzqwx/3+xDSFlUXmeBReFbwWcGkIUD0p7gEFh5Z4t8vjF8yLuwOKoJvNyJqE8NBJ0x39XuVWWI
1PE0zURk0Ru9M6S3AoJsOs2Lzm0Q3Qq04CfqiFLFezQhNjP3bc78GCn3LmSVTwOj6W/SItqgCNMI
m6+wdPFxBWJtg7OfERBc3U0/CG02Dy4vh3h99AG8UtSWnhgWu61TyXjpshFyqb4s+nEvaTy/lnrR
9h9ysdvIDL+FNJxDq6uZynPLRfxjFY+5egdoKnfF2nye2LnDfZrFzXA9Lsc71Tbv3a+VxiAmm3ng
iO5M0Uy/LXV98+Vt+VNFRLRe25czyYTErUhRnXOy6UDhvEGqymk3DB2q5aOxLJOqdlEYzIgkhgQf
Ys32AOwyYvwWkEJMRO0ms90LGGCiYtUwQczYclWE4WUbIrpn+WD53uOUR0cBUCY3cJHBNT+DFRvA
e9PpWnX5A/q08pQHXYn2z0y15vmX2OWBf+VHaxFleM8fqpok/K7s0W/qE5kix0IVhIuONlShuMQJ
aUT94CeXgrm0jb0jlQGA4b9xAfJsFUu7lyUSWqqF+LnyuCyF+5Zkw17eK+rKM9FevFg3GTwKm4qX
iVIg8UzXKgk+k1ckXcBvRbk9nGpUQ73vj22w2VMbi4EAguLQW4zhl79FCn1hnFX/jC8RmZNvDwcp
oMnCGflfxz7GkjjS9ZU1faOzHqsqxPKblYFqQ2UB3To65l8LYk6qp1WbmQ8/NMXBrsUKunaURTD7
hDVRiH7RIjI2Mj4IMGRHFMfffMwnwmxeLJmK/3tNYHe4Fyl6sLWs4YM1sux4x62pgACEz7PrSnCJ
3PssUiv96mNLLjNMe/026YAMr1E+r0lay6hHCfes6gVcBo2ak6uMDL8oxrcHfXTdQ5KS0W7kvFsA
fQC6x7OVDgDCoqNJDSF01wVJwYQ9LzeWPUqeDO/L0jee6LBR41AcuGkySk6ASWUn7O+Vh7DrPnsX
vNN4rbcuE9O+uGamRWcBtao/oC/wncq532JkQlbqDEfFnCzwazfgEp0BFQjAkKU5vgOVDr9pEzJ2
+i5MgPC/4d0EHOgI7/wTFDX0U8vQFKFWkHolO2yYIsx5Q6FTcfyKiH6Zk7OqNBtMnaNYXvIwghcY
1v7CR+o4gwfY3R//d9WBza2kbaEr5+sK/pii0h4mrnF1bSt9pQ2ArJ71wKGn3B4TQSaFzU1VmQf2
jagR+P4bYAiWh0JfnwmTttHWwckzaG4eoCGiY4iEkXES5iT6hL755V/oyIPGNkMvuPOlt/Q8tQcY
78zv/BOmGRxXduVtdtvcDd+8QJowvEjNzcE88SC0PRM2ow9qGLRTja/bHZPPZQeCZBhUUAJ/2kSS
e9VndECIvgIqK2CRBZ9HX7mt/dostg+oyHzEwk36VIcPQp660ayG+nalDdiJiXGxisvyJTqv7yaO
D7m6MAGckVkHVp/9TGDpTI1pw1aIzj5BqMULsM/uEkAxEIMCatLCnd/j/s0/Sx5NshmLH+K5unIM
Ru53aa3D5plO4aKETwHXinrvzMcdXEbt3S9V5iP3Sn7L0QGQwWrMrKdP0KvMIeNUVyJicFEL94Le
mCjvCZKH8IoOrWM1rMtiMIDvwneVqju7/bP5vePAt7SuKDceH0q+iLHWmkQ/SZsHOIrVKHyEcXZk
ne0mfqCyQoTSf3iZgV9I5UYeqVowIdHIS//9jJ2pBSKOP/ilhvtwBHzhrQEPxSJrcmeXn6ztg7j6
1FMOaL0cZ0s6fSTNRMY/H4Dm1gp/rWdSe6DhpvPRWFajwI86SwgTM/5tI5YVv+6YFPd7dJcsFKGM
lUhO62uIIVDennGeLkw50HfCNHkaNb+GIcg8CT9IxkvLlBWMsvrbvPcZWA7wWKvjiFokT/TLzcEK
W/dMXFSL/0DcFgkZvbTWvdkBau3mpimMk5n633+R28I0jmafIIYtumVzAq6uitCcszj6yjoi4cJi
NfXbpn0DRbIA3c2ciEcxvtCXlp6TnsxOlklAoU9Y8q310vFViAErQkDRYWL4KKoxVLDxH7TZ+HSc
i5dBw/BevIcTRkwAeJ1lHtGeUEkQt19GbZuuurCJw6/qu3jzRbNS7p0hubAW8VaI5XL0cU6JwdEP
GRJrFbHBwJuNRKly43ieIZK9Z5QhmE8nkhdvMEGeY4T0DfFw+S/uje4AxDZ3xSORDX4OJKrv75mJ
RR4T3kw0Z5vdWhjnsu1cUSkyNxU61kwK8YG0ZaS5Q44sU08SdIZg0R3UQpPhboeG+T216CqoId0D
j4YBKqohtWAWAmedjEcceoCNaZ6vEVmhFBEGhg+89v+hAKjdBipx8WVaQuPOHY65r0bEbopMwNb1
qSUbo3x4Uxt89jbXrGdZhEbBBV0dv/bz8krBydSq+REDHgGsk7DXJKL6FNUMlAoGUDIHzqhBg4pN
6JmKY1Vp75Oot/A6AMAC3WQXLRLVvvxImu5Pm2CWHgICOjXqY1FYg3z3TDXQ8ViS3fK6MxyvOVbf
oHtLQqsgJYd8qBUFCLkWjOrtG7FMmwoPM1flwQjw0I0A2d2o1xfb8KaBVz1rL/DR1gz5VPEa2qat
uAS8qm40HX4IBDQtkmGdv4PHsLhFKOMHVY1UINosMr8mWaNHDT+SMgMOO3G+DFaRi1KZGZ5iChnA
pLqTcH1DYWFKi4MRnBVU9xK7/9I35JxNLfM+TGXqykEetgoLL+u8wnhtCdAofzey5cp00LUarHgC
9dJIkY86GgvFj5QCYCU3wVqVHD3rBVJeEQ2/d83tSileq/WEnmQQFdPPhHQD/OBHdpWC1oeUw43V
07PVEIUkmTTXOw50e2CGOUFNX4/EUI++DhWd6uqEeZESTfJBxNj7OjmaziQZuheFbG8Gg3CiaYqn
szQfo9Cmb2mWt1NpcqjdwVKV/NzeOo/NSQfo3mjTgEDv5pXT94uSR1GB9qO1L710dUgU52wEox0S
hq1T8zZnwni8Im7BF/8jM2SF+tFn/Td6a/ffkFh4cBjfeAmUVfsVnTfwuuyK5hvOmdWiDtwnJ/x8
viCdT9749Kuzpg2Kiu/BYV1DdF/YS+P4ybm9N0bYhTev17W75xyiAY9+kD2AbkKVx1LaogiBhTwY
Eu9itQ8U9/V7cu7vspVXUyfc4y0DRX+5nOOvxjOoyRGA3Po3yw3MzEmF7GnSJVkCjHF4rkBPPgdv
V4rLeQHWy52/Enj30a3MvE3u436smFzvN/2XRLZpra++ztLPK8UzSomBCPolFW+HtOturMJM5uV1
dp44djmj6yUlt+yEHnYR5s4Urm/+hWDhI3K8n4HDhCCfK7VW95t6F5TsRgHuFHUNCA5cGsqoNJ72
Nxkn31RGs2k8bXj0hAUa8Yum2bsiOyokwxasKufGCruXp7KRvdiFCGS6XUd1KnG4C/gKPm4mcSjy
W2cX0B2ywpN+fiRNzihSNLIOL7oWZZMcQOfv0ZntyWzPUXQWENw2iO6pXV9TlMoD15iM5nXiBxtl
mzwBDmeeR6DeCEiXBOlN0W6BDigER76RFs+bCjKYvgZ2ZgXB79yMdxv0I4onlQvTyEAfV1Y6VNqm
9XvXo+zBqR8v44H+v/Uw5kBS5vfmcT8Fyez9LVu/A2C5/wyPvJ8WMVTxVjL1edM7G9iKUCO1vnpK
AgWYwK/30F/LHaFD4Jc5gkbkz7j4x4t8HOlqPZD0bT8ABZvQ5zQCcj+kkaMYSSoG9XMAS4OHZ8Ld
tc6Z+mBckQdkutxL/YBZgEAsQCmgsWepjwfnCnBgJOJn3qo8cQVSKmoCoNzSedmM+5tKzEXuNCTQ
iwQwEi8A0JAGdOJ9U8F0ytipqbrRcEvpfqcmKFXXvPKmIplwY0FN3cVMz4BaMILNODLycBi1/Hf1
mUnhaM7cOcNgYy/3d3qfjYqGg/luxt7Fj6WWiJZln97hzCGIwzTF32T83jNkgDdJ88+Y/FoCcpSO
WXPHY/5YMUkqn5Fv5z0f0oZUyYEcY93Q1eP8Dsk654xWNu4dhRNUYE2LlC0mL7HKfM/kmi0UHSNx
fWsNu7IE22TBAxr8KAo9VLgCye8+WBxZGijH98yJpunLxQ7neyio6Nje9qkLBuq0q2tZz6i6hSB7
/2UjDPezbN9U7dnqKorAAnoM3ME2ONqfdSk0+rbKhR5ezBmSc/4y0RZrKX/XhLO82cnV0zcb465T
f3rtO10gWwXmwEhkEARjK1zaavkL+9xNWhG1PGzztmOJvTW4IxlRvcc5iGfo5keCfoB2LnksyyFE
DTP3hi9YljjIyFQx39TEN3OZ28QgTcj6HXbd8KrIFdUjAZoHe8zOLquew5I5PecYZrlW9nH3lzfs
doVxFSH9NiRInZrznewaqq7e9iTH0AifsjpzpBLa/hj9oGTZGYv5J/Sl+4hZR/JNanB12euV3acj
6plnH/4d03gEGsPlUMjkzjYUt8416nJQ/IFqBokBUfMvRq4WgUhmIALoxROWjRpR4yVKJC48aYKd
O8jqJLNFy3OH5axTYPJfnJprLMC3ewKbcBcZTYVJYsf51m5uFRJCj4z3Nb0w/8CHhN/yYSu0IWkp
h/+nUSptQ8UgKCVOO/Z2QCC2Z/CberBTQF90WYrtfUZ8ZhKP9EJWdsFwi5lxwcG1oSywlLv/kVGn
WJK7jX1X+ytyvEq6NVGtadBTs6eLtiaR1TT8jwAvpz9dvNGfOUeAmAN3eBZ7n32ULgU/xAJCPbyf
EGo7BLY/bP7ToNRavWa8/R18aqttfMQmdG2sxwLbP6Do7GGOmYm7WV1lGkhRkZRzcHTiffKKpTuq
bZjgtqOBS5RXIbgVlpU2btV5TEp/Hjg4cH2IRyasRwAWit3Hvh3guC9XjA9+v3A6oY23jDgXrT8X
zMblEtFtmG+ul3SZv6gF515jvzGZqqU627CyjvKWzPrCVc9Er//XSkYSJb5ehlhh6ZMDtROztmBP
CcVVtD6EoaAXJLvl8fi46HzEPctey4eLpvwx1kD+3JtCD4l4nWrd8gQbg1+QMkvo0k+5nKJcNrI6
MzProL386gYg5pJlrmdpC1QtZ0tV5G0CSSLZLJaaexL/9wk3jttgJhwGZdaU04xpbg3pTCCtadKL
RKZCpo0p9Zy0C7J3v8Wvz7poHmzabgdWPHAScHjq+fnxPnDnG+xGB2USyp7doIPs7X/aQR79MP8R
VV63e19/HBw2qNuT7oUvncisk7nxQamz9XFoi6Kl3W8hD4bwTZFgmF0Z8gGkIdbzZ+vJR2u+sHzo
V0hNZsfwaJaBH8HAE8Krx1XKiFqbWaw3VFx1Nc0v/u52Opxnz9QlRez9XXDfxp1oRj4CnnPpQnhl
tw3JF1jgCSpfoGj/2TnYCvfkLX1121YWmQ11uAm2agYupPsVlQ5ECkWm29VmczWw2gqhCppMoO9q
0yx4nnaoMm3vzIuV0fp1XASC+EPWfMYshMxEdcRp7xZEQfZ8CheDALjqB780c7Oul6iA/R5iwJ/2
nHhHMiO/kWSnTR2HipdkQZZrqoccDq6Kp67XmDSmmoR86GyuKN1WKbW2NQNaeDzLFSO0Wp7uSW4c
uoYMaWg1XrAWUosYiPuDCMkL25E9+CR+Os9WNfkezwymkrh0bQYe13DSaHe2ca6Eo47IS+M8lITL
gS5AfXc1bjP0+dj5a6DE98i+WBGWfEJQN7ZyXwkE0XcTzSXzsJNQ0gkSJfaM2NG7ZgOwI5aaNjMq
mtHS6tcVeojCMOxMZyyZwX3oshFwFFgmyxuat46uBjHpelogggGwFvj3LO729kKydI0qoGG44feb
J5/KMvA4JAyt/Xguq13THpcc2d+15uY+7JjjT/dC926zb3ExnceHvsXpWTYJR8QANy93x46kaDsH
JOyK8xKfqV71IeHi3Oa735CK6qusYjVe0lW3R6qo6vNMpKrV84usdivqQFpgtphEfPfL79yBaSDE
mOkyuxepi7yAyWnWs2ET40zcEOs/vVAfpLMxQk9fCmSYUggtBr8L7HTTw8099EUcEbOxjyjzBkUf
ZMj/ltiz1E6/No7qJv+Me25jssC7HsYCnHt1K51i6V97c/rORnCsDXSkNpY1cgyHn+ue0ZC9btfB
HioGMzxSVtXwW5NH4aNhLHBM0o0YR7IAcn32w8O+anNHVqS9hoojOpOyt5DVV28aH3XFGB+47iA0
Jsb6oQE7ApgiKBr43u61mBGZXB4joqRB/loc8Bo2AmprpFZnSnfGlYjlZNQFbZzYzCs8tVFMHkDl
kBFCgx97ZEWsl2nzslqix93Z4D+5Zs0mFrvNHqFuxgxEpC6/lES/8r708+eXdg2J/Y/ivjpAghbu
QuAe5xqN+N+ynaUGC1LayZkTzvlBqPaWOE4rQnPyVgugryldcHHIkr0q6MDW21uf5GK1IE2pEjqY
pUMi0x6sUOs4LuFHh8yKwv8VsrPfWuBRHAfNZ08JO7rm+6sGtCvoL2lj739g37ND82xPzk62NgIx
vYoSQUGmkyOqDzk69ccZ+e9jWMmJvrpKuOk2sxzE1xvJ5YOVdMyQrg2F72vouJZ0ulJtel30Bgf4
2ajHMnX6nf1/I0e7FmL3swSt653bXGByCcVLWWwMTibiIPd92RHZAWUJD1mGdlKy2N0Nmj6MuB0M
EUeUUD3v15/UKGBRi21WpsNsAeQ1+xh8zkAgMJcJPALMoJ7BMweb0P0zVHPCHHe1xy33LPAo8y/X
kJZd8SEPglStQzg2q1WiJ92l9TAoVFUuHxg0m4l6CydZcTNDPRgq8yxYKf0NFw1+rtzzJWyDO9Xh
JWqTOcuVgeSTLrSqAo6f6fkJbssDWTkMZU6dnUKXLnhRBAZpIoGyzqZbGrgheOPyP2+omas53y/9
i6/o+8lLReGqAmTx99mBKDxp1BEaQ9InLx6M3b1J4uNV8zauPxP7YrnlMrURf8U3/BXnqbiw3s/7
/2ETL5kh8NTHJWU27qpTsE5sastN95xo/ScSHWuwZPQF5zJvHa2TfGgGkLWxTvL68j/wtdfFzUEU
jqezlO3eg5/B+e/tLkkB3cjDQBmNRwYPnbubpfeHSsNgFLlO1VVAgMKRYKCC12N405daZ5/ezOM2
REZPkHTk/e4gUxcrvQxdbCZiv+Gdqrv+2mi6/lMHSV3kG0dAe2Y2ou0YaqFuAQfP7yNNonCPNyvX
z7pGC0E0aLl5cXVwkz6NYhIiggF6V0j2LiQR/eg3FfuNclnf4i27+/BYzAZZPh1PLSAc6cOTgfwy
Ltvdk6YwdJaP/8aHDfaVUA+BPidrQedjXwTxh2ffj38P921cQ0uaJUGy+Pd+YKQU+lOIYiadAzgF
301QnOcdvItGXYcVinKqPmCgk90r3uc9rp5C4osi2foHX37qg2LALxXSSxxefyX8KEBoyouoczZS
hrZv8cKg7cbR8q51UUhaImqShMQ0LX0bSkUR5Mpc8GASdqCo+VpiT+RfxadpziNbwP1QeVQhUQvU
/NoRB/ujZswA+OaL70u5V/CrSPmVACQRHeO9VsOCL8lvQz3Edg9cWUrncjaPB7TaHJKZ7f/pZ1FG
dh7g0lv25neB+yZAv5WGySPYjMMAKfkgOLtJz5qEr7wKSiKysKO39WAL+wpSuTT9IbG+k0kpaAqg
CSaeOsaPsNWjME+aSGDK8JfykCltrRvBszkrV/oD29A2aMagDFRiu4doFgt2fDjDqfAK420+kFaw
5zaMZ0lFlUoTOgwOunt1CMl3kE57fOAFf8+QeGX688pW0x/ACTe+1cgbLQVnGladjwNRiYeerA96
92OkvLeBiPgt47sLAeRqURv3INd608KguJjzdxFR8ev++9d532SKnHRBQJ320aUhnIIOhgwMoTrC
y7F1ptZLpHVTwcjyfHpHm/iGrvGKw1M8XzIeAo/Et7Mtb1leIJTTwW0Uw0VIIw31OJUC5MW2DmTi
lNKy7XX4glyPZgRWl8biLtQaJ09BCc2BKk7+NR2UiwoSr7REpbO+7DeZ8arnU3eDiNblaKwLO42t
QEtvS817V6PLR1rKWcc0MveKc2GgGvp4cQ492eh7m3nj4WAudh8P/wAk7qE5VLjNfjZ69stTqRkd
AFr2HLrPhaC3TIt/O2+Gr/iBtoESPjE5WRZ4YiF414L4IdmD9BPPVqAZtHPAQwlThJRSlZOUvCyV
N4Relg0K4uURKI0cXySsX8jYpyO5slKVG9Knppm5ynz9E6PWjfqT9XLCq5n7hM8kYRr+1g2km9cW
qXBahRYIiyUskxWsXzPJ2NgLx7yeBWd/Cvy0/4k67/PFsm/iNC0RKqLcemM0PVe2IiiwKVgGbSi9
xp5DwVvakey6SV/rMCe7F1c1dfLSkQ40jBAJT6m2M0CGh/h3aeGJPr89TD+u3i4tIXHS5yHZUwMd
TxkB2GvAtErk+BR7rLH5OmzYEvHP9CaVWRz0+TRjKG9MfcprtGIkg/Eo3pxr7p/b248PSrhzJz6L
JSbDzRuYNCYVEk7jarA/hsRwg4kOZhEkjwikM9jB8f9YGY6Xf/F089VUyNEDCikU138NmomseJVh
QMBodB+tvNWmF/mj3NM3JG2yZEtzsj26LAUclQYAIQC+PBYiI14JDsPWuOTXaHQmzg0sq4WZBZUZ
amXjj8ukkyEMKyoVTw8mIj6RMSPLAGUSlhiLImRlv0EUp7qKNoRssVfIDG3+fDIUwHPpljGJQW1O
LmxrdLmIcSttEzCE1BVjvphaNfIh6WX1OJqmtGhePQvx0iDWq7ITCNnD3/abE/PCdQR57UfgvGiX
Gik54+r2wBIWYG7RR6DwlvbnVvF/4qJW0DAwughxgmNKV7QzCTcTtTztRqD9Y/w0j7gwUFADSaKs
SAE1igkVZt3LkpomSCmMeM9Rk8DXDcBj6d59YPdqDCDbAxYlYESVwCd1NE8ySwq4CZcir5C3VjOm
mjgT+qHuWt/Tt1vQiSvAnfXYhwFD6JsqVt2YOtqUAb4dFXoFTbporpv7aymEvtEzGQ/9qAAdbEJD
mzmpLBWoLlScyLBvSbDU/pYpDGUXe/cXWlazfQ5w7ZvoK2yFDImB/gejJLXmOogGx6wob0aFwrpS
aQalGKS14NyqcziTt6lZFe7au8oLt3l4RBSV0kK0A+VS7DMmLEV58CNZ5RHYar2BsEedeoL7ZNNd
tTiJZ0kiZxmc+07eL5ANXOwRzss3hIKoaLvOQB0olGEIC46Uhu5xW72N2+epBG2NsW5SYyjcvDcJ
9h7R+b9kYKHKq3HEgr09y3SkVmUhGmN8k9uwyEY5nYm4pWynKo+XmbVHlLrFSNgfY9eSQDW96ULj
pfwfz0Yev6ZoF/HjxtZ6M6YMmDIVrxSfb/zarTAKhzRdhUU5Oe5a17VsN8hgAA9/jkEuYVdCDytl
slJNhk1UOgDIWMNIsim9BOh36xOlxrPn68uC6rguDwD7VpJ8vR9i/zOvJ8z1ef/s0ZVGq5zQr2aQ
hilacLVxaVYxxJ4HXl+q+pZLuWFjkXLOrV5+ZHiw0ACofHre7Ied1IsRUEKue9gbqEg15sGMCv0y
jSspaAgG9+2aWkoxcE4bMJADaf9Uenvwlnp6iY1WuCiiSJ+4MB7U8ILQNjIChQj6kDOYPTvH8Zg0
QKkm/7wahv9/o5MZ9VhgXMonTc1caobSrWhfR3UPu5qsr/cI5R2ySXBMoOEiUndoigijfxUJ1fKs
wYN4jQs3SGhjJTAAS8K8slt6Hv8NaIKYitTw+HsRc8FdRnoGj3P7mwGlX4IPReQXGhazH0vPcluD
a44Ayq8Bkqjuvya2uiktflA3FH+lLlcS/DGWhbcqeYJWW0L4Y2MaIsJ8QZ4Elgdxh3ZnYSk81vE1
bVPLXXnOsmbPe8tdTaZVDKYn1YhgPQIE73KauZXNv4FYhZ1OwVj9jWLK27WzBJktjis5VpPVJh5F
NajRvTQ+v8rYvM8els7ygPF5U7rzWsGumWM2tWCim8Se/push8ud3IAOsRpUr8Xu+eu3nHOCEAsB
xFXx5NXaQ97ty9pwmtNPMpU87rG53onrD7X7Zo4oAHbyc6SkauXwH/0M5145+1YRy58S2cdsLxkQ
64Jo97Z1hlcSvVhC1Qf2cLeW2VwqgoByLgKjlp1mLp7OobFId2Wf5MWjm6wTW4dPW+XqFaN4V9N7
skfNqBWCwMZu6N3XBvrWmQM1sILZLTegq+ZUep1OXyOMSEXy3NHuiKkhOGe1CB5djyKrkw/z6z4X
cgpPMK5AEDGddCR7nNLjBr/rYtnVU0HPwUnKaZy2ETqij8mfcDJkvxSh62V2FQxsCjDVoo16Bt8b
578K0NbqSlTolZ27qIINRdyco4OBi6QKU1DT1iFruwy6bQUOE7VERZmRo00viAdAkU6/O6Dx99vj
7PDd+eti9UvuwZB5OWxvuilwKByNVNg18jiInJlg75dXxOwpIfIY4LLEpMUsdmInrgfqyZSo3bYD
Ltrz7D+AmgONla1nqX6z+QKugkmJTHviNxOVl/3Pu+JoTuVTmle01RpAtEAYZWtneiIxqsjqgb93
bjaEObRQo9IqYHYc5PUjx+/rJxk6nVNlmMbbaCzn/vUTq4IJF3qScpVQXuSqGe0c3UT/9qo7B8oS
CCGZ2r0CH1oXPuanjmtWulbzL8OSJGbioAYCT1jwI0MhXezl+NOrKPn7OFYqm6xGhtvNz8DcKmXy
3urDCjqdcNzoiVUYzZIyAsh26eju/zSXTIH45PcKrReNGS4yMUqADZU3kSYk8N4LEgkZqTNbGXhU
xiZSXS0G8tb3xQ9/lojThnTmRxXoT4TMhsnO0favhnHd5LHIsUMmQRASOe7k/Usx/uA40Utg4HCt
SL+AdikFcb4iQ9QOlC6r0syXtyZOd6Anr/qSmQAWOPGtrd+OAoogPtuAfuc8FMHWsPmZ119svWrF
Nvm7MfoUm7mkNZjGD6MLKh5BQ/DA1O1cBb9W45L4THzm1/km4Jo6sP4oHRlrH0+sqvl3QikU58cR
PSYIfIaZPQOgm7XIOtiwnypc97IvGk8ppAv7r3jsI6OCk4yZa6uhTWCOiVLHa6LnnMmX+kiGPhaG
8Se1WgfdFfgIJ8zqBvZCZZQR4vlvi5SL2SxgrhtMS307kDCP6N5RUqC2OugIePA2CTBCN4nF6MCd
KCtf0hj3ZTgCWjCqYsveyjV804wmW+iq+QjUc0unchh8nVW5RF0InIXqemNrSgwpImb3xGuB8eH3
xb3iO9CU6e0BslPX8aMa/hIZ8J0xbd4zKiYBs2BwMkhpEU5EjO77/e8T+vnXqMt2dxCY9P1phUDl
NCvJnAq1ZjYmSepvjOVbHuj/m/G3SZAV8xSrVUgVpIFsMNN4fcL794PTzIuG1waj9VSm4r5jBYSE
RfsMHtkstuGoSMEp8XCnXFmqAS3hPdtYGxpPHxfqrcZXBQqUYK1by38nWcI58XpXCl52+0FTtxGh
cxfmU6Rpp3b2uhJvAMjjSd9zUBNWvbvznYKIiqJmvIATTVfoPnj2iSQNIeE6rtGKOHxhn22cpJnX
pVe43N7/9NapabX2ubbD3vq4Yhue4ifeySP0az6XYZEgvS1xRd1z20gHwWLfTBKvllDqUD2rvauY
wUqgvD8pKpS0M5unNMn+4adHlKmgTOzRJJws0mGbjhROkhVdWMPWNd4q+HVqCVnDh0l6TTFmL9/H
r0uwEYBS7YMB0IUebxyGcUi+VQAOLW4/Pj7MXHTV70CWu9mAEhcGglh7NAM0JgleXEOZmsK6+gPt
jtwX3x41GimRzFJDsdClGeo8viLxjUqusRRJN/mLydH7HkYFdPk1oloHo9Q30nJNE95/xfY2WyFx
iF9jp1kt44zWwQTvOaE4apWQN4s8jNkycpGFwimEi2PnMslxRjNg0tvHioFCUF+deUronkOzpjU/
ekTAkigJdbnzEyn/87XTfmoP+30o64s+yluDz2M6dHLgN15OIEbpZn9HoqR8snj/5LZSTUk6D+T6
eCscu0Ms4aNS0Vos2EaCi8TZy50iBn0ZtHwAUTL2FLNlsUPeYKDRsjp4hgZ+rlPDSnB3DPScuDPb
vEHn6blWRL3Ezb39DTFBkry5r8FNqOg0RKxwhChFwgMI+xpPTxRk8Huc+xdEpUp0f7KQlBI4gBm/
t4Ezdca4cSXfq5L5Maa/5p8z2FQfjEItCth6khyCpi8xoHGKb0QIptMY2uC0xQiDqdhZzpSvE8EB
0aO3ljowUewDnpNEuTlz9LE7bKLB0NXyPQZ9Pvu9Gi93L4q2ZgW1OFvbxtiyvd5ItrKgDcsnU63l
5vSY9RKaDHCo+yBBr/dTNneu1W7D0C6QDpOTzoCsU5ZRi2iwv3q9c0CcTtNIJcB7QUMfu6p9l8ws
7j3WcOWPOU2oGcqf8q0Qn0ie6pVOCDODXKINP0F2ELOnwoigufiTWpR/lUqOdtcC6je6IN4rqp2A
wuqyJQdIOcEFoYwkB7eUduTfjkwH7sWF28pk9GE/9OiO8/lyzrx5kG+MpmWsnG8c8JX3Ler0OhR2
oCpMPACwvxLcoNVU/DRwPIcIhwHaeuqLMgPhPhgpuIsms1SqQEN4lhjdqDtREHPr/UXsjFTt7IWQ
QX1WTGc5fB+LEAVKm0NGz9GoDUz+pF6cs6F8MnPbjcpF1+icA+2212wEla0IA+ymTE3EVCeFnpz2
2PT4hkJqng4vfwYr7KoQ5ad5m1DdueBuE/+CVzVj8+BvApryc2Oz8Fq1lvtxcky38OdlpbE01R4d
5l/EtWN5/PKn4tZcV/2zeiDWpwmgDc2TwT+Yj9BRtVzk+0svGqE0tMQKT8eN340nPTawyNjg9H9r
0TRPGRk+7ZYyBEbXVrsYdnSiDEicUjuGkmMKgVPEQT51b8w8H8GV208o2GVHx40ZtIKZxg/1N9YV
wSu4R9v/8ktJ/pQdow0arbn5oXrcGAo492qGCsCLD21tT40vFljx2dStNmvUw0xxmq5B843eiKzZ
My13IRe/KJDtTiY3KQLuU0bLpuLnUtks3T/VDjiEx3UR6qMonjRFUVzRQKqLI8uiB9MejF5TU6t8
zQkThT6EThnWDoaYo57wpvxb2k5zEpr1+18l28vvqd8rNb12F4Io0LfZACKQFPDjgIFfN8Vpb25Z
Zm6neRf5sAoN8yfEpIm90JzxA2MqYIq7tW52LmEnK3NLOlFO3LtQ9tmg5nmUdBnBN8UEZj2annHQ
gKow0N4PzbRU+s6wQdVkJ5gqpPRptARTu0mX5qoTJGgPGIWKVzGi6oC9AO53AgHK9JWgK/P+NfmV
7VBxsnD9uODu3mlx6tBzozfKFwvaNpQipKMEQ3MXLMa663OJTw1FLGXVp33sO/su8f2aXamRaYOH
CdnBriEPS4JdnSxdIt50TLe/+I1voobkB7H4mCcT8vodW5zm37iPOi1UgfiVYTl8V6+VHp1OLLxQ
ysaDLrOOH/vNmF9m52rC5mN7v12wHHtv8blM6jiLGp/He504Lr/Orf0+uyUlt9Fjahhj/mlgNbs/
7xqFI4D67uQ553B2WBjQfoaJSxMl1JVdPdTyNehq3BahEERhkIytoIaAqkgZxdcAmKE5H3DXOc2l
d5JQyxYg8jDNX9f+bgMrautaISh8gCVhlXljGvwtjRA12uthjRBRulEg9blz1WO5hNhvjdExcass
iYnY6jywJrW/bho8woVOfqpY7/ibOGRppWXBXNs3WK3tyz8ERX7nlQy+Dxerz/+DOuHsQbbCsoju
4Q84/nxj732yRKhJ4fbQWmpaBkYeXDZZnoOMnh+fTxSSj6dSZhrFFuHh9n9aFnOd7nc2Das7HDml
TCd3PVrV7K44m+KDxrqJQ4SPVtE6RjZlQTmPAQ+U6/bYJ8+DuDN9m8jCak2BskGugpJFx7AkZ+Aa
4A+EkIG+yvDLxuuGFDHIVVuooLiXYuW6LPI49wTZiMMI83Dk6EW1SFn0D+EaurutQko9XuxKEfdM
g22nRt62XVGHF6Gim4LhspU5EcT8QTet6VrjY3jHPjl9rNMmgHGty+x5pa/BjuS34ngnQlzSeA0e
P8k0PNvkDNI/HSfHVhnfkaxe5O+xVaMQEgGxBW1+II9JrnMqbXfW3VQLIGTGvDtmHKJ74Usvl7BS
6tYTiSCGtAX1Cvh2uLQ/I7t6DChBZK9UeztiH/pwqeJp7X6zWCrGr3G+JDFIcagGcinvpxcpyHt9
icFuuRDH83vPMuGwTC+VBZtqrwWmD7rh5RV3XQsxu6THkVj+FKujNJYL6l/znLm0eSnB89q1cUln
lKVHUzo0Ujr07aTyOnUb7YFEp7Y3mKa6PvX8HS0vSLDr6fXNZ8cuMyKZJN6J9a6ZDlor3zBjUyMA
IblAiQI4XouHXdFHf3Cjxb8jEtovBWOu3WKACA2pUfBsbub9Hm9UTV/pcVCAb0mnWQf2hbpnNTpS
oCkBfzp1hzV6tCOzRY+KQoywN/QL5h3iJgWY/AfaUjzIClk8KRdqAiURkDr1EPXZ6gUJSgWtBOkZ
twF1wmHW7F4Gt+9AkX3OWrei/oyDbMarYBAcQnp8S/WOBxXJ6eU/iRXTPzpU7TiupqVgTNSoKttv
P+gjsOAtXWXy+QIlmQO1YDl08X2fNjcqEG+O/tiIWx4LSGOxarSm9DDL3pseRn9CF5LTGPRshCSP
BIhdOIAzD2h3/gkMv5zHGPm/20uFBWCeCA4R6h6tFd6RP8aZreIGsWqXXFDw1O5c6y7n2Gjkg7/s
n8Zk/uB8RL1pVXpxJq05hhryuUQeFrDDKfi2+3X2UX/m8M6vclwnJ3TIXTiAjhFxBO8WjHj4C6C6
DuOpQ/2tLhYDLVUwk4rHW5onK+88ssXxOxhMxR+A1QVSzT/BVhPnON49GwBpjGCh7VvUM2o9GKQD
Y8WF9d0SdQefr7nr4buSYHKY0Tj5chtZmpuLetnMhXa8JCdWeIn3c3uNT8UmLpBTFAMURy9sc6t+
r7C3T1/TCZbv/zOnoWylr40pgdQeFi9WSqjGAJ1CM1PseMIqdxhb8lVIKkkC/vu8t+frDOIZG46t
ru1nxgXpB3OEXWN8uilh+Z5oraknXSbMLAN9IU6Fe7iEjOFcl4VhsZpbZn7X7cQrVwCKD3p53DCD
sNUbANuBIxntAq5376EUnjXxzUg6zN0J0Mq12ODJneDo38pvG1ryzVNsFZQk6tlbxvt1y/q75KFG
HnBy5UDhjflsAvepZbCC8rScFLiseY6fRFlYc27cdvU8TkbuyzTX/IjwYwcq1a1yY4doL4eObhvc
1ssGFutU10lGBjYqtem4NFX03oZmj59wEhv7XcILatiJq88ytMyvITml9/+wQaigYCngmxSfLc4V
Pyxz/13I68cnNrYXFXCYMhZcuxdJ+894FYcj7lzDcK5yuYmYYNE1HFx3S9uvQchd/wvWwgazB4OY
Tw557lff7GtMgLAPu+VPRgl6tgFF0C56MtFloEzaR9Intl+fdPGxtlgPVt6l37t2HaA0IYQ6Jc0a
BlLm6KRqcTNVlG+JsdXVbGmTWoRLVsqCleGpa10f3mNWaXo6bPkhQb4yZI0uWH4czoTuLz+h+5wp
NkXkIVbFvENcUAoQbFrfQBui2LFv/qkf1Zfg64POjfcM76yeNtEQUJzv+UVw8Zb1xxCDVkxoLFdB
A0sk7BXVDfi0YBRe3ug2UZvI/HRp6wh7XPdDQX1f6cuvOZclYsc7PjgiTqsa3aorvbcC6VhTGNNE
zZFyjFOVZam+Kequy2yxV5DfMFAxraN3xw8qwVCfZFCQP/PawXywhMCnDf/3ia8PPez2OngJyQTs
mKiMulKIQnunLWdb0FXQhyMfUqYc/Xqaep48ZRVfNaGmNJF+CGUc7jk74H1KS/g0A9HwZRrQp0zr
7bKY4vo+/9P+dLpatrxy+L5qtjtygeljuzHQSzmfB5Y2fVywMnhthfp/OhKQFAlCXp3nO19KFNCy
3Frrju1U4fVPoUc6ANYt9BvR7x1/aVnHWBGOY5FnlgMdBB5qkzhfVAlsyEJfywa8kSQm3Jh6+irh
cqrvlhQjGmo3PmnsbDvkiWCKCyfIn4YrHm5cuoy68s5KAQYgtu7ppGZahRxImnMbR7YUVlW7J1K5
kkbNowUmcLel9M5OPuWGG9YWQL3t2z3jl+HaFddSzblBX+HDBg4H0m4e8q1OXZEsHnsTnJgCAqKC
Y20Ap81W+39zsliptRalt4LFq82fr0xSw5l08sdICyMapFLE2UepBTV4Z57PiQOg9/64FjGttp2y
hK/p65Q6nbDqrO6AhndrH19FGO5UdHtjWYxRm8tw/oB+CJ5/S1XfgcMj9mMe5Gl9ATBkrOrsu0B4
nMmTbXl1+jQPdFDog6Q0sD3ZBR9IxOoOCmIyVEjU0lP1QDZOSrpNPqpyaLDid1eeXcQl1+h4USsK
b/zH0SMVzAGTbYjR1PLr6tx6pB4cO6bW6j/Ys+Au1gpz2y+EZ40elcOvtJgiuwlaaSfwZUC4RChw
CE1GcxlvcfS5jqjqYeqbE0xjfg0Xs0J063ZTv6z+JBbI1xS6J8Lbu4dTykLy8Gn17qTm9eM5W1JW
JujHjy/YheqCxJAM5HBMaJK2SHXDsLIyfutH9w0Ybc0tVJahKBGQDYda8TNjUID+21HF91L/AOfS
hAfym+WEEyij6O9sKsbeGeAR6f3kCYBfyt2OIayVYc3mVSQtNZT0kFYtXcey1sKd5qkPVg6pqHJ5
IY+st5ysDSQKurNeA4xixyfatT+q5xc6EKZRBOagSHvPKmtPPOgTuB+KjjFdfyYum1TiUKsgXjSi
iDIuF3+dcXHiYdWyhZzrHdIB+9ZOujR30hPYY1dvQI9MnTFhabiWhN76c34BKxOHyhhr04eo3KOV
Ww45H+49CoTOMWvjAxpapZmPSqLpp0FcmYl6J6gSlUStcfwWLgR4Zt+8gq8tkhDuNcJAXbJ5Va7k
7tEQ3mysNdF0PTD9mY5/vf3i3P43QUt/MovxFaddfDHikxuNS2+S17vFZF0qWcSi3x6qoAR7JgCa
bHt5cr6fwuehLx4DRXID9fTCDyeeZbsoPPaV0d4/jFq+zJSa+ZcoFeQfQu+hZ3hD/iZU3bVWG7yo
lMJNdmzuI7ZT2gwBVsS4S3mqL3VMI5DyEhzZdiWqiEVWjQoM8xvLpXzQCY1guZXPwpa9DLwfd0Vs
jqTaQYlasKJHRqYRh2OTiNYMX9dWecqtBc4IagKHQVq14bAzM/Vico/7xuNuUPjwQRU0Dh6R9aux
olAKtErOhg5gGu+DgcdnMzy4zJgLna7HimhXvvoTN+P7t/s0y6qHLxy7KuhixYtNGzY2Ie0sujCv
4stfvYbcofKkX8Rnh+Pe6djw43zMT1wkuZ/nS/FC2w6TS3cWzn/ZNrhEnvSl/fi1PMKloTYLqIUw
uJp03uuB5yUEsCIC08DmtGJjNH64CQmE4UVWypSriW6vGziE03yYnDsulXGb9Db2i2w8KeZwjVMT
xVHV8DSZqy1Hp6mAbeOPSVQKGU/hVYlVIfmVdYFFiivaTSd59OiHFvXXFjWo+lYVvzElh4PtmTHA
xjLoRu7IINPr0OSgRv0DobBgXSx+px5m+4QE5vlMPdwJ2MgELb0MkfnSGrDCsal9cDvpmX0+6VrB
Wqq089fa39Rzk2/Q2PfMHCOm4zKcklcvrMQq35pmLpDCHf+8JwNCN0u23MTbaFRlBO6A+8YkwLz6
9FFsCfswcYYQx3aYL7lEkdlNsF/i31AmXtce+OtFdTdqn+hi+n9x4+nffBjDue6hgevqcLBLrCIs
556OWwhXtHrbqiZ2/l9VLtivFZ9bnRrvd4BMzT6umVSF4Jgis8Hd0+G3q69S70Z1gngv+RYaNOfP
jKfDWtuoRqUXRPSCjX65b7obF7txVrzWVj8ZAdtQ1dnq3zNDL5+Zwdsn1f6qqfQVrcoASaFaySh4
JkFBUs0uth5FRV27gwn6BLTjI6vD3fuBB9CHwjGvBZPy86kLuhbsCExNzFUTQ3ezuJbhQir7rXTo
h+U2XVxckvFvIuSU9n6xg1d4kEhJO8gUuUYehc+f3pvtY7fs26IwpigfG9AdNJx5GJNy9DnaS/cm
0dTVnTZrEV0mNEpkFrDgV4Vi3g98GyFaTWthx3xbldaV0aFi4gSYfHu9Bj8GDwV8KykdSdfOAs0l
ysSCDefr8G7Fr/n2JuWqi6RbvuOkmaN94yryUlsBCIOaNKJ/ydZA3PGyCgxLCidOqNHGxnj7Uwbf
5L9Q4V/9sgqPqpr2J/fyfk7oXzOqbij+7iG9vWDhWu70vn9IjOMZGSu98LdNiu/4qBTSd2cBIs5z
0vFhkI5LNc8AL9/BY+EUTZrIk9b/aN74nwCc4YxJ2NwfLbTaCZ51EKbqvi8smv/piEuqmAfV+eD/
j909iUF1RgpkKxq6MmKB/8qulZtGw9OxfQJpH6gKjQq1PYxbzOhC1bmIDohsQaJxES7DBCQjsnJW
GiYHA12UpayWBW7SuTkVclRLF8+i77SONWsMplp75NOWZwZgEFVoIqAuhD/5JTQKZ3xFiQnpIGaC
8EdHo4rsEnI9sb7mOt+hKPiBOD7KS8IqSASYakKDnY8bw675QtkfFFI0SxF8eE41CZN0fSfVrF3s
zvQq3hKjBjsWG+Yt20J7F7Ho8CoK8tDrvYYCwCU6KZHYhfnOTpkPD7S6CcCXHIt2RwkGr7esqVt7
h0tEo5KV1oq/sI3soaekuNB4wzzegFFvPpJM8dPcC3Ycl8lMDBPCtC55rBOLa1kYUNi7oAzQ5KOw
g9eoSlSzn8bkvhkxVzvz619BwQUonjCb7rKy7ZOhzRwrMxK0OWv9PA+41cafkQ5nQgXp+N5IRd1C
YqSyKRY1XUwk8DQSJeFHVozw1uFov/n5eDoZvMoEe3eZ7kSFURb/YCwOv2F/hlIzrKRn3ZwyP+mC
p3lHSOP6WhV/Fym83Kg6EYRMJLThMEmoNGb9JFGpH9puyPzw9ZnM1oX4KWZchGdHuGGmBYV8BE50
8Tu+2Y5F3yPw51Q1HiQt12tzOg/UzEbsXF7RE66TTl7FkVCL0szO2jMJgXT9N9ueVpxV6RP27T9j
iEnIUQ4EHcSM2kGCX+yWVh4kodb7YUHdzV6Vp046mmd6BQUEOhkgb9My0UYLCHd1otgh/nQXPXPh
b2paqSt/0HbrqUs4KJTcsF/m1K4Sws/fhfJ8JiqclQR+XioZpD9aN/Y8R+plLPTxZUhUsZTUvcbS
9fZXcZbWYQjFWJJOqXqoo6bPhiP+UdEvtxzbaPjcGtWdKNsoH2qgbHr+iznFSwsnsKE6bz9wfU8o
Gr1G9TRlbh8QyvrUsrRyWvBuINwFDhh1xjgivnCVkWOf8pAhU0bDXqzTCtRlIAdwSsqf+p7LpCwf
qTuWC/mSoYKazMllE7HoJxFYgGxzWb5Uvsv6qNLHrQa1yQT7I6Kr40Mi1RStc3oHH1EfvACClTtS
RK4OzSn0o4QusmcPPsFsKjNNbSIDVUbK+IZTCdsnhAlN06ATQTPYky3CuxsBoVKM/CCDR9ldyLo9
7iC+X4SsuwSACc+luwzyo/kfUO+MBQNeZ8axm7D7ifeX5zJBp70jaAMZB4jJ0fDcm42Nw87BDkC9
fSW3Oph6f36tp23MZ1WYOGPhDbeiFSdljwJFf9bdhe0svHKUQe7/269MwjURc9PhWS4O4wD4fywK
awDaiKdX1n079fdET29LeF2/HBW1Boo5jzrZdKFAsC40hcwVHJOxk4c+HcY1JYBLTWOON9nP6DOP
UXe7TZhqheMmeIl6L6b7CnmMKxZDdDrNaKRRPipgShwhmqEtuJ3Ts6FVvjjGCII5BKRfjNhT5Oi7
tXnONx+uuZnnIqZi414FJiGPnoL7YtXZSeu6kxENkDI7fhkeATLwO2R4S3QNGrrgdVTtpyqnaMbb
rBvmPn3atOCNYOe9WtDdewNgaq21p4/YnFxHz02VvQMxu9Lrbe25zKGIpEFt+ITyz38hAOqu5j7c
VwcOrn1eQk9de93jPCKNlQ8SYoE1dFyR25bHuARUXCWWHTgozjzVPXycnKMNntQFV+Q5w/wDxbBV
syIeKrxIKxe/15YMdmYKB3Um/dVY4ExZq1gZsK1i8jGpvNZHiSSWayhxqJfLdhmgyGiJR8/FkObL
T/6MqaLipT2CJCiHocmiRdK00+whwdFodSUCSlRx2SXGBwQrte8RUlP8Pz5rVvSa8J3Gk/1b0UvY
LF9we9V5fQeMUP25dqVioAQwzoNPpIKc7+JLkeoUdBJ4ny/s3srHnQKh7m/+VTGW1GiWch4VEyie
e3cNKfzr9/3xGGCCzYbA9BbQpAiETF+MY0oirrX/lsMOaDLSVuF5SJtGeHRuTiIwpPQfelerZ/3Z
FGlmPTOn1tJ7oZN06Yjo0Fi/tgiN11+MzkgIUWRqWQn9rzOej1IzimSkqKUHvMUZnabI5FgRCgA8
0smR6vEBgE06qjH0Fmn8xEhaNEEr5Iox1GHadIKks4gMKHT1EI1h45nLhgf5tsB3gO1wNgx3ZdwB
2xcbOplOLlte4JiWzX6AyfSCYwTQPXCbryLuj3JnPzHUipBUf89iBWmij0y7oSHrLsdOKYZ2zPzp
OpGeCBZweLS9co6PBiSKGQTXNZUoBGwvRZ6WzMIkqY5mFpQqtKaNwXd/riaJQ4s4pvoNwm3QS5yV
SCiZQXebcN8z2trb/hCB8MSiM/5EdnKeKFpRqkCxQcaojpK6LqVz68s/QkEWFOD/Wq9L6eVwEwA2
JYVDnGFIPavicTDev7os7ZaJNyuw6dIzJ5DMcSpU+3vWKRxiuYofCX1noHWX96CgeJJAGnr8ONzu
vNoxz5pbNU7wkfiE4FZwMft+MzrCuapCNfhGn7rN4Gj3AmYs7A+UNyk/UEriQ26wzRUVeIwi/OoO
YEHUv7iJO+7aKDAfc4g7bOeh/1TMZmgjCWgT2xYJzaHz9Ujhx3UynlhCYuM/xSXr4KVW6cUxY6IK
5WiC0pN+zJnxgE6uHa9uWWzldRIWfKbUkKmpIesf3f47nvvpS2La2xtAAs7MybB61RxEaW4ZmyV1
5gZ6Bcw6g06MvMFFH4ABPunaxT2o3CN/YCpWC0tlEhuLFI4ZRAgVZEfJmPv8pGP6RqqEFvoaQyfh
L2XlCB6cooq0y+QID+WMk0LOICmiu3aO7PJ24FlJ6kgAMhHnv+HbG/JeHwIMy19KkZkCwuDaBinp
JTuqum9AAssaGzUG1Ag4+cDXL5SiGWIRrLai76A2Yj+qjWBw9+1gDzwZ+5zBfPdzY9k+W71qfakS
qoOYl/zitpYdYzbEjJxpg8lrPS09ttSzEXnPd7yJqVbwavcNjaRUTbj9BxL4rFZMW0oFHpzRxcQ7
vKZw+L4lgRpibc3HbYNo6Dz1YpYKlhxlsswmTdpcJxNPzEjdthzYYY5xd5VRwhFoZJymxsrSzUzp
LkOjBtG04mUbzcJWcLlMOipn1kpNMZQ26tArhwVAKHcc32v94lOqdjw0LseWZD5sdxpdJ32j91I1
J/hrKGYBc//NWOrq1IfsgnQ8mNCx/437Yb5wqPqhJwzgQcGztEZVFqTKT3mX2ahIheoz9IzyGvSi
5nSksXHoPmQiTsPZFDyiTKRT/MYkf+igchNIfxegGc0BJ3Zs2DNm192Vskay6RRFfdIipdFAX8Bl
80bHfjZPwPzdHF4DDDwgSUR8DuhRcb2Qxvpx2Qp+boedcHn1RsqVUdGth8Eg9Ah9WH8VsAPRTNUY
2ErkESYvVxVTKD3duaG+KQ2j7j8/kjuZKqAP00Y8MOaMMNmZmBSdBxKggWbY7+IrUCdwaWzdaUrw
+yeFtN7rSSkBGt6ITK32P8CoqPbZEWDrqOji/2O/kmIYn5cVrnh5Aifi1v+D1nincTinpKl3UScW
OMF4vM+VYUFcFcduc8G/TmfA9QXaK1X2+UvzzuXAMEWD5gb7JgLMl+DxMaOFGILrDivq+bcXr4dR
8j4gN1KYMo+6jZmAfybowRJDVlJbks0G0kXg5GUT9Ww1OGosKIPCFZ/afWHUA56vWMJv7Gjxg70f
QThwvGc8BFN3XR5J/YwIyfP4Dd6OYMs80sXmcp00XGdC5ftVktvQ3Mw7TKR+cdagNrAcVQWkeu1U
uYcHXdwpuBYsDRFElONXYTekr9iqQnFJwDdyodA7nNWh3H7KsvaDUzNSEHnbW2Vg5FpySZmqjuVF
3hdsIzT56ZAi0AmWnTHI2kreqWvqlbc2xSCduCApJNEES+hOBZkdI9nse5SEc/CLjUmveoUEgudh
jKIHgRsLWoV4b8iUZy2qFM7Ia3irdz/RJJkIhsi4rVCOYmJ7KpFeYjthymDu9lPFXtOO5K3Z92R5
16J1MNHKzByVDDLo6Yi05LzPknC1BA4IYVUwgYicAJej0pp2aqX2WJuvCVgGIPhsuvMVf7sY5NRL
Z67vkO8AG0XrpWy+2AI3Mg86+s7rOgk4njkOZbUq3VCxKhMxOeS88sLe9dn++toQJ96qjclr4q4k
0z7txYw18xB9DbkvwBq4Q+7V01iczVu1X2qxmsyRYPxfmRwi6eMWzZwWrBbLu1VDIeKUVeh0u4wp
deii+UXgIYXA4GuJf0Y/orwXIeCK9n5MbXw+ZxHDDH+icgkIfCjK71Et5F6wSmgiteun6e5tyllf
LpLGi2+lkF+QAkunGZ57IbUx/mSFRhhGNlvHt7rXOdTAYzQAPvQOxnql5TXnJDotBmeFWyCXNa10
Lkoe8avLnpXi/bVBWj8pPzw9SYU1ttnS3j//nYIMP2ts9qXqM9DxStnVahTkgOuVhuGIrDN93tgV
EwCjB/txv0VPASjaxSQ2OIWU2VEJmkcjfN6wYgS6ye0d1Jc17kSww+svQ2xt4GwRIYrrl4HgNvPj
tRMqi3gLLIk9mv/mwA8vVK8D/Tg44y2ON/o0nrKsQKc/QQ85pJvYLjC65viSyJhKIccnyynSWXb/
Vqy71KcU7uKKUXMqy1EttUv0ZUbmHzpURJuzJOdZBpqNEfIBP4VWoAfCfoJxfiCAxhMg28zWiX7L
Afcs4a3j92UFpqOtCVs1wPfkecfq8rE3tB0R/tzxeNdb1pe6s0DFTQlShuxJU5IFUwzIRm/c0kxB
uIUv3zwtiwhyRpfE5zYe7sOK7vCPiGx/lIKDcaOY394tSrOsrOLoYgLA+6zSunwSA5rXotmHAfvw
KJ9tWpo9t29/xK35hPS/PTRAOHWXb9RNZ2lK5OUBxpLNvBIMKXBu0jmjK1VkFGgoXPmxTiZQ0eLc
XoYATGKrJwUqaBBJ0PeWSGuV2zF9TOMiL38ofRbgzfKP63Q8EVSQpa74eorQkBSvsVQnZ7//9yAB
Zb0E8Gdh4X1eHE+sReZqkoWbHnl7rm8zzZzr0fqcfDbp2SklhYZdD//XIfXkpoAkdDZxj4sCcXXL
ej5s1iJ532wbWAnADwl8uv7k629QXEZXN8QjybSf5LdN//ens47MHkA3txxOpfkps4azPOhpeJPi
orMKCd6E4AhhSjrlXjXI4OnXdnmUoBQjONqbiWq/Ii+ny7vdN66/zA/1HpPB77TNSwk6F9V1XPCT
rEmEFUmrzqJPN7TL2rS7qfv21MX3rhEnTAT8tQw+aS5KPqWJHBPBM+MFetc+CyrO7EAAdEhkkTQN
bxefSmJS59ysRtSiNRxIgUxQsJk/B4i8As98wob+gSUIKYEiE+tlddVWYRzpMeXOKFojG4QScJAR
7gLYjV+lTSpbs3P6vwvsAQTYiGVQVDod3zsi8mB7CxXYjIEzldKIoq45ieO0XLAaWvbbSW8ev4eW
efY5RNY9SHLhOz1MwxIWcA8NiBnDWoUdGeqmf4O8IU8xvwbgsZIXtK3sXuygkGiH2TbhfhIBdzHT
aBSdWK4JffFjUlgO9VqJ2L60POfOM4jzWLq4i/awc4u1nbxYf6LWZYAQom8+ouUGZpPK2/7y4zXv
fuNGpu6JHcrR8f6i3xnGGCqXhPXQmY/yvzLnnKrnAw/VQaQ/mHCBVSL89268k6R3n0Q6lcumP0VW
AdwjFhNwkbfOzgAFjMa9LsegqziiNQ9bi1MMi7EN3DKFtKIBL6PukEPZOky3N5vIodAVgE3VQcsn
ETHvksZDtquN3iLpX1tqNOLPDbZ0CFDHFLYdcMvU6eNk7OMwAVI+iin3OfJsy5Yff7btEWRSUdXw
16ofxCodOD/kDApTuQiX/N6Rh6r7cNHfChXYY+fS5Ojc+cB0iZS7dq+9QIN2N9V5y8f7zrz3QPIG
PeVKEq8VBeBc9ArlUaT8db/twemiKVgqFFqfrb+UFgkhOJ33C749hGWTnWwt79PxzIs5I+RD6o3I
pwo7g3RQMFZLYHDmX7OoZxEXX3z+DwEEe+ob0xZ0aoNo9iAiTu1alSHUDJzZX5r1ccZ3/89RW1D/
YB5KTaIH4ZAxtuf7rG8DeYDE5nP8NkFJyKnwRIE7j+5Lq8D5QsQ8IoNHa+FT4Bd4M71wWD39t/+d
5gD9wPC2/6cRL73fhy0P2zFsxcIrFi0UjnEoQED4TOX8Qp6ZaJiCO+OuBDCL87UgZT0GLAZ4E/I2
XFPs5NAC9i7DkZTPBnC4ElPRV5Cq21ldKb0jzWIZe1nDB8AivgeAkI/fNa47lNrQru/n8FICqtgC
m1YfAuXVs/Dp8JusheSJj2pvCzkF+kknxao44z6ndQdW6sj8Lczfes6Z+mWoeYEveIKt20E5IOdo
QQd0Kwd7pdRTVJT95Kvk7Kq5XDGdyC5sTcHfcEWlOUJeIkHfqAAjwZPMRBZ5LtqOLhbnBC8FrHZs
XISN41NDcIEVV7ZPTzDANRVjNjTjJNoRpzoNXvhPBg9tiZ6WxE9q3mOi2N5rTAz+rr8ax20LIyUa
EdtoswVrKFJfNN/qJbvrIY1c/DJfwv4DW29keOS5EPMLXHbT+ISCu4ZfGaERSEYzEG/EAQzkQ1hP
jTi5eBYL85q/kZgTimtaXJGt7XRZVEWGWhtoJbJBtz74GLE1+nCCc6JBVL2thpE8J5mCv54RiKRl
GLWdGLgpi7qJxnnTZCiM32xOWaAwNdrUGQDsBYp7F1ekRX9BBn6NsIjVVzwP8PmW/uC8toiVCvMr
J87jNzAIjdpLcpgJRXTzPlReJI7qTJJdgyx7dllwJ/UyTSWG4geWD/4u9BZPBwJvVJkKRb1yN0g3
UVZCGUgNz5WtdFtWAnxgCdBWXVUCgoJxZdah1K/5ed5Fv8SG2yrHsX/yOfRplAsRfZ2KFgd7eQM0
AxJcPzm2qrRYy6YhJLXkWLQ618c0Hysq+TnhIOMUaXvC1YlemgBgd/jElpsd/qzlmGr7HvyQmSPs
XePZLavUl8NL/gZh1mvM230UwCcDK7dpjI+kpAPhgA+Ig+qJ1SDw4HbRwO5QqdQ6sZy99x5XwkZo
iNOgwD34Il9UypfgzDO2TSPomhuWhKiE4V5gszuWT04BrkRaNzk4aoQHpexwDLhCHkZ/E4WSqjZB
O2FAo1pDuev/yHWHFOqReUpOfrMM2W8s8Yn8A4wkvHZ1k2SYBNf+sN7fvwfwjx7Qq8YIi0fSDXRU
yzd4rxN5sfh0DOZxcTpiM3mBFF4zbab6TUzDcIwMnD0N4XYPFkNGXcsJUM6ix46gDtKd6SMGKOnI
Nd+ay0V1O6VvfDhpa5mDxX+vKHWZZcHUImknhcqwGx8bQSo+Y327vintQIOKNKCWUQ2tzTzZwDBu
3I5fNrsP4V7GH4HgC9K8YDXo8wDGxaBkEvDF/+hlqc4xEIOo3LoVezpNYqbsMCXcOaMqnTD/QSff
FitlrpH6FAKHTTepNqhtA/r0twC5wpKeff2J0/SI7kU5rlDHXG4u8ugtejLVrY1Lps2ptBCcmcer
oGcRVdA77fz/LMeybFb1W3MxS9Qc0lGLBBiYcOJyt59ZwbLoqLMw3193GPZZ6a31R6ESv5uQppRr
rsnEMj+VNnHlr3xelPpOQUjWhhmRCq9RP2fsZmFHonVIYfkxHFjvbp51s9weJfIBU3OiCkx2gFj9
czQdryRrGfHuJkq/id7irxRLzRMbRi7EQyhjmegPQUtWuKP0m5vx12XioyYCUZdVh/fTpuYA+jkJ
ppxzYOsv6zG39VoXplHfhpvnd2z4RQSOaSK+WzOWDEIw3yEH+VDox8apv2L05piqnxTBWI+TzqMt
4fBz4gxr2L2JkHz+z+DUdpCTw7QTr6qxcc97uZc4MgzVuzrfodZ8fqXEwwcmN5YJCsiV0dXDKxZ6
YLlfFOp0M07LzT4dsxih1UeqaVL7smm7g1Eqx4p1YkQVyXoMGWNbYL2b8n61NIf438Eg9bNmhCAR
7WoPJ/cZ1BkoNCqcmY5Rk5zawDdLWlcxkCFJ8JyIM+NzMbunS6DDLurP39nRcVnETXBJQdZS+v2w
vk6Cf1v5GR6jrCNUDv9TyVkyH0x7YG5tAVFZy1eexGZcUdPYmGuNBYPCAZKie11zPIzFVsOBX9ws
cck+GgcAVviGpL83e0A/zJDgo/95FvJLtVTK1f2aMzZ44efI6LlkUi1xAXuLuiSbu+Vx7yzlqP1K
xfx/rPGOxmvtnAlIkOtCRp2EY2s3fXlFyaopTCMH5NIO1MH6Rdz6Y7vbLoXZtcSLlpU58DS5vlqg
Yjnahh2v/xrqY/AC+jDPOq+QQCuP2xMgUNa0pJwxg8U1rQzwYk15zmljA4wo9MXJLflkGXra86+9
qGo0tJYia72aCW2njDRfUnz0OaNymhBGSiLRC2/70MekTbnglv07u3BTF03XcuEcxX4fync1S1jE
jAKfm0b7RAj11ha8t0nzQQty6Zfx1e4QYY6sRMNwMd5leRiqYOiM84ZqVd9p7qeXIkzrwxcWW8vC
z1jNbGuBGcTweAM4NyzmG9V4yFkwEw3fv4b/xt2vlXNwJmFi8/gSnT3LjZdjesBe9ycH3BbL7Xoy
LTbPQJVMYSw+bYbMsxCWsAAJMEnWslAid37sIP9fdJuBozwhIv5EcOd4wpHfTogmjsgvSfaoI6+C
uy7h0F7ZNCg0MlA0ZZPt4pRDowV/iK/SQPabI/qprY26iE/np8e/E+aFZ12xNmrYNOU1nVLPRRCn
a79Mux+xNhN2vfTQAhbkL7pnO6dkzfg+RO6Nz2h33t83JsWvsZmT85yc6sCvTwd5m/+c6BBt8myT
F6F/2TVQc38NdrtC4Y008UWUF17imDyZLGVN9FMn/wRmmIsA2eSK1KAIIAHLH42WJQJ1Texkl2td
ypfThnJNh/QcHCXBPVBqIbf/jXnIeVIBo+WpNArzVg4eoBgIzFFxcbT0oePA753O7dDiOXPk7hBk
bZdbqDvH7KIgy7jPpzqe0oqbngKfPTh3da2hTnUKX2OUvkCGKdEEmesSH+QOAmKxVZmakK9UjUMO
Rb5xkUKSz9g5CRpZSBljeleXy4THIcbwHkZCIozTdk9XEmBw5oP18TlozM4OeHvHZr6fSdEy44YB
meQ8USmtiTZUFlNtkoYUMkvEFMZcv8paDcQsWhj/e2FghgqfIaIoexQd0UvlG115lEEQ3wNA+ikm
f7OIcyJsKQyCuEKaoaLXYyMCecVdlnwMzwVXpZLjopazdXQ0XstbBQ1nEwPH9H/qu2U7OOdwarpD
a84f89joMVOeuxcrlTRiMe8GwOxnvn84li6FccytthFbSw2kbfXqJoGZ4E7xe5yriruUT5Klgl/G
Adr/w+AaAUUM67SeWzi08FSIRwj0hVrTS7s3YWYcADdmh6pRBwz42Cqky4nyca9TlBjPmzjoQOXD
jsb4/utDxrOm6A42DTHjHwbmUuRjW1/dPVBkou0J8W9TMpfeG3w6SDNhBFCKzzY3VPRYQPdU0MCY
Mvc/s4ZHN+fuzAHpVCvgdHWNoQ3UYw4g2NjTOYFaH+P1KTvxGxwrT8VPMdRUdT76k1YeKDxgwKAf
+Tz1HdlZm3cwit+mVsO/Mw+7pV/MRVGofERgRxAQYB50wA9YyO2uLOgaNJ4+ZU7Q3/isHvQsEXLd
kFc7VSygr+w01MPxxI29u6Zh+lBAlj+vxKkuWPcUi6VXVts/ZfaYSyo1WvjcV6k3xIzy5yGpXq7e
WzRhPdG0mYr69T++o27ZQny9s3BVfRlnATU6PFhAYQIWYrBuHP+s70ld3ZGSSV0z+BzJiySof9Nz
WOO8V8jZYZ6HRp+HjH13ZPEXzOzZmM+s2J/KZVaScind9NoXPCP3TopMV2DL/RHr7GqiJQgKU4eu
rPDYymcEnOnT2YpEGoeRq7Cnu7seXPLlY/wuCyZZi6XHqJ+NMZsbuF7DogUondbHm0R/YFLBoMdU
QVmzYXghqaeW4G+5InQyLse1nV7ZhNh13ztzMQPcSUI4ktYqRFVUoHqnypkbqpdX62B3c6+/g1vo
DSTQwzJMGQsrZHe1FTyTeNjq7Z2aTtBLHBaH+jEc4wbWczq7MKoHQT4ZgVG+USylKTSB9RlibAx1
d5SPP+cA4+qaWarqgFGQ7R/uzGs9Kn2T5niC1V5OnW6Aukd+ld1K6gTtAWMqObNABsQnoCpbxSdh
JnLnXZdOcl27W/sxVDagd3UGNNuw1bqqdVyv6E9d18ztpMo1ulT+/6L3/Cfmh7F8cmO3qCiS8Q2j
6RUbGI7a08cQQqeMqbEOlB7oXQ3//Qix9dy/gIA7Ek8vLae24T9Ge0SDOLOmjbkcLQdxzQy1wJXs
8BP6DhoW6QdrmFtQefXVRClyasvHCDz0Ic2MczTjr48tpUBhSSAepsIafS1GAJgiVRN9VbkIYFV/
KIm77aQFhBTcRAqpx3KH41h4sa/acP6ElnKdvC5NvK9Zy33tVWQg+/4ggwZLBRVHof6EUUHc6tlu
zDNben0gS+9YMgfvN6nWeO+VjzCNGWezf25YbnD8EFRiPKoH9rsyfdzsjwTXYmg0e6TvVO/9IIbU
tgzCUzEzY1T2uMM7A5dHjxrxIb+jAWRompklTeqyC87SwV9pxHUVXBAmfCo3mKcGPq22Sg9pPjlm
IW2FzrsA9VHK5W+qRcn1hqDQ/rMpbTOd0244FH9SXjd9X5uY+ki3Ezcdg+od+ffGMyBxpfaQf7NO
JlhErDXc3VXFVT9uGgILFmbMk8+PM/b/dz/0wIRyim8pgDQHWc3a3SZNfFY02wwdmypUDjvDFh2A
Lzhwg3OwZ0g+P808kwbmoLV5OejAHIDv6zLTQhigM/tMPQHCIsNLOFq3Hkic4tBJcpNyfj9xNFRx
oWzt3GxycmvK/Y88TEaMiBy0lVLEiqdd2B2jOrDANboaz5wg8JJo1pcoMbbJa7Qbj1scDHiKu/EM
GP9KClmNfN+YW1uRhoxCEcoedMbQXTzIN+sqU2KZRC68F2fsrzcCSp3VQfE5Oa9tWdsH+gfMYO6q
Dx9v8c7qkgU41V4r332LJaBu2Xdgo3zWRF3mylUwmG0Kr2VTfAHN+5QjzSHMJNgdVBweG8Sh5OsQ
tKqhZoMgrypRJdV+E7tHdMHcY/7fo9jP4J4Kkeo6rYHIJ/Lx08q3NLVCwHD85doRCW2gnzY2+F6q
t2n+LvzARIiz+Vp6mX/iFUCveM+n9HPxk0lzl40811ZwpaOuwLenSSSYboFIfIlg1O/cHLgMPXcd
jOhCzXV7rtjBcvzIcJOFxJRLG2+Olp0hdpbS8MJuMhKLpGXRiqHcESBAx3WhVkmCgHvCCAZZu1Dj
+NV6j4dBLO+bk4UmB75ZGNGTIsgwENQJI1o0EiYEveErr3jLdJLJQtbjsnft18hpvkQIZQnFIt6x
8mgZCwUAp/YL1p7z6S8UlqfH63TyOw/G7nydfYhomxi0vLjgCXOZakkknpLDd0hAWVc8NPzVBBFD
Kv/p0cTGrk2Y4eXYgSgCalgV12tnmy3G5KCtIgJtAVofZu7XMbIWBNvila7iwEshjyhWOvQmsZfo
QlpqHgXcHkrE0FKnb+dh2xKY/8ej0vwBVdfKmUgH3ieHJ61qKrI27LkFyuzBw85bkPjp+AJFaibo
eO3Sx1ifNEeywdhZXTAV+rULA1gmiPyWcGh45CZ7tlrKLXBTg6rRZLb8qxkl6UdiMRnLoHAodTcy
sxXnlRHqn/Xqy6ncq/+awSjK4x3qI2mLnuEdasmKMRNkmv/eQnT++ToeHzOk0qPTEd/GnQz4y/Ll
6wVlzJ7s8AZ8weMVy3YvDblv85ZRA3AMdQoVzKIMGilUuCFN5ibmQoONVzBnGvN6vxPiHlWl12vY
lwLFdO4wN0YCpCoJGQ5wPMUfpo1Kn2YeM6RL8PG/RgHhW7bTRXWTplGI/m7lBBkIj3lNZjdppoEA
6D16jyi6zsLgzyITFAXs7RJ1joOlR7sdI9td5oic9fU4LWFnxdPmdJTXtAoMyDSXOzmOljGN6VJX
dGzgjC9p06xnw+GMNpYW3plqhxjFUm+nQtox6DvBPQ8gISbyVO37auQ1XVA2tyNovXSYGSPc8c2v
T249+LfCvRFS3fBl8Antob/JxcOsdcZCI5euNY8LOat9cdtjAMmnBJoAUfzLWkX2eTfVHvWiTkjL
Wr8VbeV9eQaYtbWqpiEzo/wbglmS2TXEdBQpZrk8JTQbyEajD4RiXadoSGxljBszcUi6myo2e4+i
529fgWCLDRukJPavDpeVxsuEvVP4eyr9g4RgATxG4eO2r2S1Kq7IaLPEOZUDwefGDHlDwGlgesKf
I3nSdbMiKG9/OdNWKPM3ReAb5VURA5S9hx3EfwE+BDBLgQepu9G0sSu8sVVjX4JmXFbkP72snFDK
UbMJtamopMC9dbwEVgWSuq0u5KuVomUE1x0osJaGDm2UTeCQdOP1+gL9+ASocur4IRDOZMg04N1q
jqr4qIvyKTDtaf1Nai1SiQ4NJ2MXG0zgqLN3Nh0I97DIyn1Vey/KifN+V//mezw0GGWpxOZRy38g
Z1RN8sK0s9c96oPk62iVC69GXmDhQUj3KIZ+3UanKxtOD9uuOJeTIp6k5oQsnuP6kBn34ZavqMiq
uqtTTy9s3bpdDX6xiGWN6h8VTYlavgMFUZ85jLiyW59eehPNJKB5tgaBYQIETW9mn5khy1V1NQRk
GawDpImmVREVYYl63FI6ySkay8G8jalbhIgSN3JjsG4EMycsMJG1n7vFoqoOIaMTJPv4KZkot01z
gvvUVlsUZq3zTgM9p/tdtcr7BYT1VSkOeEI9ZzAE9gtuEr0kCKb3mGgxXVgKttqfHyS1j7pffSx8
Q7d8x2DhUQmZnOaPCdpBI1eVInum1LuCBJBNFg+JBfMvbjs4iHnkRtNCFK2ELkVCD+1No8O1yVrH
5ubMgQZol7v6ZC6HuvLlHcyErzzCDZypQRnBop7SPTITIMTP01+UWHPJWH3x72/YyE8OgUmP4nbo
nVcmdOSodmyW2JNbZZ0e8Lf/2xxkMuiuBzugpg6h12tIXE6N6bIZVpjBJMB94P1bYIR6Ri1BzKlA
CzM3lXTmjwfwqlMrsNF7o5NjUnbibBmPIAnnX2FBOve/LFxw/wIqXGk692D7zHvGqHMqG22tEaRY
q1oj2ibpkblZpEZaMi46h4Xo1ZE9RaMlm15sZpqXUlhb4m1ZjVQDKkbmbsF9Un1WkmZ2YgjMXyq8
59KnLUNMbPlmvlzOayJR/jtCaVfc/G5MW/piFZJSA4zZxWE1zZa4+kynv8cpQMa7wD/721LZZQAS
Pq4SfBzqaI4Mdx/bmMPwCw4rbzAeGUszVdgmPNqr2+zx2uHNPcR6XlI50Cv6hhNlEZm6G11KzM+Z
a3yiRXUApbWf0WiKnXcm2EdHDokx7zkwnVgOwn1hXnioVw+fapEMPe8hpeAn/kpkAHBfd3zdF0Jb
065peq+BdP4fyNKBRAKYATnsgoCJRRKJo/kyKsQ8paaADcN6zyub9EdEN1xzb+Hm8KS8T+vwHcji
QjlbHNXmTBLW8zMrnR0zm91f+YaMOM24GmTjFA1dmVqik4ZC7bO2gvMoHFBNcyRhtHJIcNdDGwQT
+QfHBvmdv0IWGJcmmixrmHRkvIVNcjwzrem9XDtQwPk0R26Pu5Db7sZuqJiFQ+xwQleJPLmmPEJx
yD08yQKInkPOelZQIkVH+xrhTsFppOTK4E/r9fnEk70JV4SiZX7H//BZ7fKOcyUxva9xloXQFWTY
cziJHi7MVFgRLCkzEI5wUu2X4qseMW9xRGdIbp9CD7RY+YQ80h0BjUMMNUamkFlK1xBpXT5yJfVb
pKeO4gWkUWGVU016nvDfO+ug+TiCw7th2reglrsyOVcjh+mL+vLvtPWS4LMYjR0Xzw3th+r2pJJK
GfJNOUXydWuT9+HH/dNBExbeJYMMarDRbm+fmkVsmE/MqJ8665XYGEuMu2C7UQajcfLc6Dfkrc4B
H+p/8srUigkVXpWLlmAOH6VwreSwG3Y0m54058wBO8g+6JhF1Z+ewloS/HSgy+6bkkhsd6/esUyQ
sPFI85YIkb1k5p1/YE171SP55xojH5qyjStCC3noWX9DeILX8X6gOUTNZMVGsUFjY+YvYMEaQ9E+
N7OXwxXpZNCKkOXSQBr2BB8lajdQSJWTYecQb8NwUrL79ySS61F10wcRNq5i6jFD70l77FwBu1bz
PmyMIt/1m/luEY99fxE9UkJVc0eJkea4bZPIRlsB/KwnB0yM9e8GyQ+LR94M5B6NBO6Cte8UxyvS
+24zaWin6/m7iOFCwSzWthEwtZYqcgzuZ5fBgSU5nyBf0bJTh/OBKqidLA7V4YcghIelbqsS5Q8B
nAzBf8noYxgBaIlH/Z0nhf+nN9HbJXRIHu7S6iTjFGm39u4PFym4saanOE+wIY5TrvaXH7nBJhCp
wC3a6Gc9yyMSVwHt6tWiWAkhMAmOXydVYNAmG0JC70Z87F6u5wcDHiJSaTEmfZ2ga7dqawJrg9lS
UmvAa9sA9r8SgxEGHWgVZjmvRb2phbEG9L1AofDVDgxkde3Jy0gW7sEzocZKbtAe8MRavqF4NZpL
l349l17Jg1X4GRQedsO6TR2R3llU7PnOF30lFzvXAQQgQx4cBwUeoy5xgAf0/qHX0p33mVAo2s8Q
wijRuLuPc1VSt+p0eShiJKfRsvLYYpsV1gO1Wop+WCvIvdSu8itMiTqLZwuVXz7ldSpesqRxaEq6
yedL9+NY/gGjXxtHLWMsJhWEBQTl658aNhgRzuYnfCtG8LzIfoIpHjvbAbrnanGvbB+u6/tkzvXW
SOS/Yl/QFlL8sqhRMO0jXOT89Pze+Yoh3JinS8XIzsAZNC5ryvnqntm5tW9ZxbiTeJyQZ3u7QGI4
ze0PMd8LIJTZQso6kA311Njp41q0M2I+8M1hOqCfN62pyF/97To/kOI1mLDCGdloK9OOTZ8g1me/
/ABlany2jWprObV7wQa/Zms8M7vsfB8lBkpNUxRxEwplbgIh6MseIiemqN2ZZgPgPDbG6Megv10i
frpS+nN1WKrNI9m7IfB7UOLVc5hFMK8hKTmV1ZVowu2Y3rJWmcvINL0xZxvQcpmyD1cvdfMgbPF+
7WsstPbAR6gEombqqhzjJHlXaD+kaKlP/pR+CmNXECjUMssIJxGK1Ykn/Rby3ffxWqSDiHGukZ2r
oLOo394q/Bj+KrxGqiFCSQmOZbjXZ6+C8B4RbwMfFyb7BRAXhTcJs2iymH9zdjU8yfkNcnbwIwNl
n3OstXFnykWffIRbLODa9L3GNwrGVfNgOzzWHTJAHTeDxa7EooGy+uqVWKHyjj5bII9NhF9o4/3L
dovdqE+K3M23EgLghgfAI8V9jOemk5wPPPvCTCXM+AU3zzxa8rWon/3wnq/HFm0k+eypIIjPP7FU
YDSp5q2A529SgkbChcDu3cXwDdJNintdXwqH0r6tC/oxBBkKO9gpQpxUt7ldA+7hRWv2TzUIBtDK
kcdjnSpqgTimPJT04L0MDJV+uB8IXpxL0rFDLvdXBGcRJQcZqHhUe2SjQGZnzBY81J0vpIfugCj+
9fGc9DdowUt/CAJM4Yrmy5+yZJ7TczpcX+oN5jgQRlEwtaP9PwNyc0bkVVnai99h/A60CPJFUIOE
8uWXLy9AhqadqpeLpYhHV/b0MR8mzBwJ0ARaV6RlduS7sle9J4LBxfq7CddzVP0DMy85ebamDu8q
HZVwpOgYjE96HF9o8JD2QgQUmIgYbAl/Zz8rUym4d19gNfv7d610lQp5EqWpmCXOMr6Zn8/0sP88
AULa2trcBVgDI/sr5kqI0nWWui+MsEitUZEQjMah2BkWqsRUjadXzk3mU9934HpduO2VB/82envG
FWSlxo6/t00wjmoi7Stn/WPABP6+OUnNKUE16YFO07FBJ4i5WoCf3dYkIS40Fk8WOkVrqBvt0uHr
+GEQa0xSUB5TOQA6om/EXt/ImaxMlbxyAMy9h1YUzS2BcNF4qLQbZNfhuc7EezZCNwJ+GmZwPyse
TQmshmTkev68t2f3A41wxbg6VxEdi2V1KLY/hmVt+8CWAPCebNT7kebLXyDaDRCsrDKVq71YHAHw
V/S3zCVWlLZv0c4WDvUOIkjB0390HTUahUL3Kd0mAiA+jKZiF4YsZGjJtCQ5RCu+FFFG5Tu/RD/J
p9FRi8xFL5/b7nlNiFmSBjFZAb0i+1aeXppzwsocMYsAFx2wnBO8iJE1K33TWjoL49ToEKDh9HGl
Wx9UTs02BVJTsCmXyDH2gVYOCWp0Cn9cVpmYRYVKCWo5KigNtW4ysE3P4wx8IBW0xgyr2IShoBj1
ubjkgCz4c8uWF12ZYlvyQbNhmnfv78PwN7AJv94EAmyUg4ROM0+EU8RJqZg2J5OvKEUd1Nb6Kcdj
Onj8ooNW0cfggVYO5r3+QNXH+wV5nAofMexAt21vzuMONZXK5xUQ3nxOaZFXPTGwQ+8YanKegXcC
Y3nH4QJio0DBvesC5xedJT7/N1nYc+ngrvsXGqzH9IGPytOzHH496NTyNw5bN3yRZa+XTWFv0I9b
QT5ggbEk3z4yOXnMfTQRnbjULKcAHX0EsqbZdzESptgaXre7gexrIqyQCIruxAjGH4MJ6KsGMgW9
OZZRXJq+nl/By0YQNJ9DFT+WU5T/jqgLJdsK7/CvJVUMSkyVB/ZAwD0C7cod5BNv/sha/yJaO7xJ
Wc1Qj7v48/CBr4uV7rjO/W8drJorM+1ANntODNipFWLkqr5dq4yobrk6fecvP3M4T46SItd2E7XH
iIhcHBdQKPBmj9wilPnZ8DfygAxnPFzdINT6zB5PtOkTDRwMJspXfGbp8g6TOX5nV3vWOpinnjYH
Dmx24vZ5SgTPWUKd3JErVaY20gXDCiWgDRGQ63h86ZVPsWjJ10Ong2xIcp2/+zj1HFDVGsSs4APY
ZIP2vhaWJ4fHDTpnnH1cSARXhaLHV/AOV9AThDghJol8bST9hJ3BF/KjvNzLM08iT1Amk9yp77FK
im0gV+khxDhU3vVlrJReFaSqdAr2FpwBg8Ki9RTBgRvKFK7Db5xDCHISbSD3kK0SINkea6dtcjcM
uOfw60cwNag9P31auI+K2RtnsQZzk6+MB2BGyMu8z6XdPHibnR9XyKKcGq1wiJb7A/He729mexIn
int9+ON19lUHlprJW5Y1++xxrEEi/h/Ta6+xjzHlWJMC0aqvtVZCZJ/An3jx33v1+9SRxEoyv8at
U1RZGZpclf894Ch4haPGuqreiWECbJU4XSx7WpWU2nnWWyLjxpRqUO5tgSG5orua53oSaXey6lVA
IYqPmSFY12wrMCEkakmgR3gBGL3SqCHq06gGnUyDN0A7DK7w04XZ78auuruXulH7/L3fKSMe1EsW
/6K8G4UEJFooDgyZ7zXbncFLJa0oPgcHh78cXRAMjhSgckT0bWCGNpanI6/SBuu1qEwIl73zKYzH
TW6eY8+VDXWpXIXsv2pq2Ttjs3miim8NJ2uXa3PXpPTekwTl6IjlH+PGiPSo8htZbeOkF/+8fDth
txEJbjR0jlX/a4esuP4YrZ/j5OXA3YDBQjR7WejpMR9kkk91QcjdntvXnOw9bqFOeDJfV4wEZt7X
PTcNWQBfpLhuI5WXPhgPk3TP3pSFPiRN/BR0yXx9MfGJ1/llYc1oY62VVZdpJh67pCniWK6WZb/h
MkdbK9doXR5/ZBPmnUvmeuwPnOf/7o+GaiOVsZMExUWq7t1bOTHijSNuqQCUtPY3M1vRT664Un06
D4fIPhz9P2ylZiPAhRDkZ5RdiCscrfWjEA+6EwJWd11b3E0Q1C6I0zxJmjtJscqGomGL4x2nHSsq
hoHmUZatG9bgu72e4FwLtVkTgRy6CNy3Z9fD0ZtT7deb0/+QOT3FIyfQBBgU3AImnJyrpaxxqTS9
h1MvPrUMqGEykb/CL5PzsXE/eNqs6hUWjp4w6t0BJ6aIlheaVI0PzHBzPoo4jVjCa1Y+LH8JtFrt
lZu321No3SAyDSORBSRsKoj88Tj0TheVQQzgm6eFkTO/COuyMdQjOMP+E/lsfGjIce8yK5TPjK8Y
FBoHkG6csihvrv4GzY7nO78yh+KTimXa8P42bv75eLV9hK/66X0vJ9L9t5B7rxgdooFTMU4gdaqT
FJidtz0kKg6mzrpzKpG5+CC/KQyC6na2Taj8D1lRaf4Xc49TZS8KExE0wxiyy86QUjS5w/Q8hyF5
f2STgCpcIuH2qnKGDKwsVB9uV5/19zfP16wP9Ey4MKaYLlyybpKdroZ2xQVyVIB20I14wODsivzq
HEih+FfW+ckoZPJCPMB8IfCbLNGgsUfUqtzWhHEtSsGVlCcaR3UVzoG7ohsYwX6D08RXT1DFjTv7
rOxRXN3M6ANsBmgfSAJw/kLdntjIkdKFYX2jVRky2akJYz7Op99Smcgyf4iw7Rv29mY8Gin/uFcG
8AXhD9JwR5syg3cUo929takcmeh1FNK56CICiiImCNtNB3r4poUZLiAeZXdJPcahbBq/JzSoKWlD
D61NGocQOVPyE1cwH4wM/t6VlFhniSlJgDTFMaf2/cOw7Y2V/IHLGBc2zKz9VXBTn4aBqYBNa/nt
1tJHgxO8arK6mqhhtYhtlgkm51TQWSdFvCjPAYTOBEvwYRLFFGjEdESSRC57GkoQWIuh+4eC7WQ8
ZQ4hCfIYFJLcDnMi3MEX6l3XDBVvsYq7CGE8vBpXnnSAW8MU5ulZfUHFllFCeWolnPAgYSr+cYue
Lj9AlELDjiv+bkVwTQi/jpK0qt8TYg2gSBMb4MuL2Mjmddn9Vlku+Q+MrWcu832MLEbhtYrYB2zo
jqddNN+WcLhFqrGZBDfzEDjjLVQJcIIt/AeqJ+f/kW4eTtEZZAWV6oz/ql7LdCA2quuHY2oj9xBI
iaCilWSqWcKwEt5YphBZ4uJ/BIRG2oPkVqryqrPDKRxupa2mjJaiWmmDNrwOSZPhDo3XISYHcsQe
zPuDzhufKJMLZMHovO+6fRFosnyf7XSeI+lOPFR9lz1YfRTvk1+ysKgeBUR1BjmPh7uPnIFTdkiO
NefVAjANntsMak2fP8yUIi/BUTlRlME2TnFOmEsjmC5jkvbu41nDVnXJm+21mLZ1a074fXsACGa0
HfhGEnWygI4Vh8mzMiu6hw3hD9+rh/RnUf//39fydrNtmKX8PaNqSAtuwp76X+X306e7zZWViNUB
+KoLXxiE4y7hAwJPD1XglKGQhVSPgYVnSi1RxcIIN4XhMOkcNcs/0zXsQtmKUkWH+eZzXTvA+Vwu
Z0SoQes4QSncGj0be5JglsCee6kGyIfonD5pEIRqRn0b0k+8Vp8aKXMxBJusuHiTmlaeLQiuoJ1V
Z9UEIK5fXCO/wcpZuO5wYrx2qR/iRyVNGqUqMNVBPx9DUiIwMSPsYusSkgbXl5HucnbFfM/Cg9Ma
eythAubMKt7IurSyW8oITx3aqDD5qo+Rb9MFpxbEt0RGQrxpN2oVCjuJrAzzXMzyg1p6Fhl3kCpS
vzBr6XjfqbWtjpJUAPVdyG4DAHNzMmhS8NooT8KUbtjig0YWrvcA9LcXDVrwqif7kiiN1NyGu8Qn
ibheu9ra1t0vWxgpLZJOJOIY8rQZ8ctv8VggCHUJF1VglDu3/LvrfP71CrjvQPLtKgtH/DWjLoP1
P+zp4CZRs55GJFUOGg0Z9EJeuIepUhOjMfVYLVm8V02ta7kB3XmibKE+/M6/6VIYCPzXEt+ssQMM
Af9rGzvEX3YGsVWuYUFTNUxjq62obAVHgTD/1jdYbGcUiJqcstRIAS/7RUeq5ZG9QZ1+9R7zZP3Y
Sqbrd1dA/MNBNCinKrk4dk9SjJBQevo/0MYGJinM2czrvrmnTcAx9OfBJwE35nzALN+DLHXxJ5dD
Cu+7M/Tm1wsUrn+2wzaH7rj3pSZUUtlKOBCTx7+6dSlzyhUIzqs8qiP3VnD5dpljIMRPaPvpHUv5
bBdzdR1pdkb1mD+Do/QBvZuKJabwr7aeXl+h3sfzLeg2NSO3Q8Ku+xCllkhqaLuGiiz3qLdVKKFz
oTMMqPgTafv5jElBARTXHJ/uhLMrm83Gb2wwXidCaj4WTE1k5rLZ7jOhbMXsoilTjVhzHrSJ6UbD
3FWQ3YpMNkOgXLGf8toZnuqeLj7GKHPXIug09ezOaPWGD+/z3+WkLJG6i1XB4i4dkXJthFJdWdN6
sZGWYlNWCD94jhjmhc2iIAHrSZOIbmOo87X1BtAP/SaIYCA1z/LYZD1cIULVOq9saTxSZbkYKlkM
2+XpEGrkgLD3TDwj2lBSvbmx9RHxiimSDccRyGK3jtCYJnWnMxdyYZy3uJAw/VqRsCElnteav5Ba
JDrpPw7kb6VZY0tX9CE1G51ll1lTDu7mf7cMpMD+ZazDSPwXUhlkKlyZlJl0w1FhbaTZOU2zAM93
naNZ/f+KPEra0JWcZ1Sgeh/GYj34UrSvVoQ7dYKk3+ZicubfgQNGKhXBmXlHX8Byd0cekmSwPPb1
fauNqI9sY+6yOZYsvpFhMG1JfwJbh0cMLNZp9JAAVGE4TuHKFfHYYOUyFfsdRTfGppx1lp86Bac4
/Xgc2rEq1sIz9ebok2lIXgR9hPPyujv6jPzSVmspR5HPB1qm0vCXZYg/1F2Wq+gh8/1V+NgUtAh7
30XGtODDGLTVBaKvt7h8Ey5RjVC6SiifzApc7fYP3bWjz3SxkQx0VC1Q3M8fNc87dZGbcGADo1DO
iQ90niHnuim7cu/oKRlut8n3aPahqMxgApF6ZBTt3f6wp+si66qbBLozrcKmEUS59ds0/YpuXA43
i0t1Oytv2mu0Ub6nZQDZGnHdh5Cp22qONrsIFk7ggArCJz7iznTowg51YQxWWUOA8/hJENeihD+v
1GDiHIInd3mnDeNExdaDUq6wN0btXNj2l+HoQptgUDhy5RuejXOVSGza396LsZnLCn9SGbnRpDJh
0YLDX0dZNT5Tc4xMPz2nVXhOgGZUtxKzRTsnMU7QVig1NZmWMRPa0BITld5TZpEAC0HMfNNwBbgp
znlIVghxL1XwbApl8aPTxd/BP6YC5ZOMnQ2ryVbPQzsvZaQ2v/nSpUzpLL7N179KQwr6hAdS5Lg1
641hlLigEL16hXypbr2ZU9jPZeBLkTfNkGcJnvcBW5XKaOksm8GnFulrXbrUtw3V+tG0CrT/YdOs
gD2+tMf+ttzg0Xg8nepFaNoGVOx3CqkkcgQEu06s81q0TpDx6eK3rgwBFXta8LdWJU8rvaeHAIf8
txMum8oTtqWTyJFY/G1H8x17EHZ5pSdNMw7270dfAuMazVtWQKFeIcMadaX2cBaUs1ko1u1o7Rzn
3ET+0tQDEkgqSG0SzaOT4/4/d3cCZ+NrJ3eMvWcnxQ1S6xw1OXNr63bbTUynY8Qyxo0/wWG9caKR
69nFApi9bbM2miuyTuXUVV7J6LxtCG3RYgJBmCnx+xUdmg5ufWnr0xkc/qlkgQUJlZOsXgysB9YJ
DeTAumCXASYCfrPd7q85FZQiz45OY69nkR0r4gvdEDzHpZcDcVURu3TThDvwMdF+gFVH27CxnhxF
O8tylF0LEv5aYNTKpzSCQGa2Xxo563qo+TLcXrWXMR4DxNNk/EkPUZaWIrnYYBAtBctN98tCWYaP
vzapK3PV93c3eqnHS1ziRWmIUp+QIXLSgPLdaqdp+JFZi0iKunOY405K8z7fvHKnKbrJsXdWP3GW
ZgXpXV7B0ch3hCnceSt9GtFCXURPceOPx3EgJXT4a2CfN/xheSx8fwiFuSHXqqyrS6nrE8gXUy5Y
ajykcOaDM96dyJxFE7iNr9YORaP3mvr7yKHkLG5HNomjx8LCV2h1QRMH4o73KzbJK4sker86pAje
7LCv6BrCVpihFy7iWoKpDFcfWDiNeX20rAkR4003Lw7zFkhjkMqj5Td5tesc24ZPwUUW5fiunoH7
kCfHxCWcJeif391zNk7Kard/9/RxIYjc2DCbFRpROc0gcuetEATmE3nCu/AwB+03/GZnISOJfDBE
tjH2Wazd0t629ZUgbioMFkONUAXCc+TqDfwQuSijoAAzN9aWGVpxDSUDuruzy0+fXhCYG9C/Qvvv
s1D4pPSJDsCIKWXUHAz1QfLJmDnuHQIKx+fcq64fUf/XXtwJgLWKTxmtfezUnGhcecG5CyVR8lOU
bniJEXvmaWmiGBUskcrVZadtnf0Bk4Ce4f0BgGHiyDNTLoWZCu6Tyr9t++9rlcotFc7Sq9vPDbVs
S/P4ftn72gZNncQB573iwJlHMfX0Y6Ujc9CjkXRncNu5vX3DbLhF6zNpPdlwuxo92C7DUyfoVVyh
gHJkefKNh+/7CvaAhDm8md0U9tyNdoXnECnHAmE98aiqEAnspxSa5EGWOrS5/ki2DIzVxnFxi6ZW
bEzTluGjcRbNLECCZGkmqIfFBToQ1J0FmOvwNVXK0p/YHTiNuvRBsNePpYb/ujY4Y3m396TKgytY
/8cCtwfWGiXr9a21STQ4BjW9eUNovwgYLRlw03QUsw02luBqNoZRbq3AiIMURtnNzbaglEizkEdt
fgmY65eZ+gAyIP71PSJQjkSf38rV6sZmwcui0k4eM2CoiRfXmusOf3p+mFZ65VzfxgsRdzj4ikuR
SaugX/BWVkw9C6VXlwy2JRctQ/8TF5inytwIKMB0Vf1H8oO4qoFVh+hDQqMEpZ3ntgAhCj6uhNaU
zaVYXC3+pQIybC0e9yTNdN/tEB2izzQBr2J/90m4+NdaCVaJE8BDk+545agbgYHW1yXpfV6uyESP
G0R3pR8pvi2pZiTzUaNzsuefIRFm/3h5sdAeGQRNKL8LqYhvfOyvLN4L2aiRpxOyINB25ZZs+LBe
Cn0elSH5l2HeThOkdkGNRYsXepBvWzaxyy324QTi7Dw9I8lB4ozMdG6S2PwbHoddBpaRm+xjJd+g
CUu21VltBOSlTyti0fL2mir5k8GVGyFjmuot/oyUaJ8EQxyGnUBp6VQMwwGl/MU4QZrHi3GdJY0w
9greMj+aPApcUijWAwTBrca7nPAwjCpb1j43YQaL8U3aBrHMZUmc6H33qb6rTOZpwOBkKaQi8BjU
9ekyitz/C+iZtIExy5T0B0two1vTmmYmXpY/ks+4XwtoAJVAexRUA7AnKDSYbjyKzqvIV9mu6qqi
MbO/evjOZ4iv/TVRjcjJcHEpBxk89tK2txqmm9KLGR6WRFY7mx05UTxvb6EhCkSCSHoxNpOo3ynj
Jx+TARsxV0W+yc9Tqy5GE76acUUCenH3TVW/0917mmFJ6U+/mQdW/mD+uayuuoOs3s1DVA8iPaa8
pq/7EmZ2Mk23H8V1J+GsPUxFzKC6nIFbHbppGewGTk0U/bLrhsi9eGuDMd/rLZYu1928OVYYxeCN
xE0WLrTjUVnUvGrm6vnQ648P4SNNHGLuHhSRuVK3vx/yf2wyMeXamDEDqzRL6xsWRz7VQ9PwB/y2
7ZZh4Zstxyv2ezJGI91YsVwDGiMQ7u0vSUuJMrUuJW9o3vErma80CGSXZUsi90HaphV05PYV2xhI
mxXzSq5ZxOXuv4vMijAvVXYv7KUgwqGfCV5i3gaKrzCMiBXRGmrL8nGTXCoiehVfiXqgCspkXgbe
ASDhDjZmsbApiguPaPJ3wUcGjP8pyA5qOwPwv4IoFFzWUWFdQwKXFzaqvGtOWn06kJKkn3ygrV48
Mx2TlmxONJ0mxIbh0a06AZ74hakjPyO4tBe8hEOA6xsoaJJV89f/gRTCdrjSgmjVVPZxdUG90OLr
6IwTn79Cx5AM0vwFzl6Dc2TDD6g64IepRM2wtuLIaXixEFISW1wUQxoB3/CjXE6V5K0DTFUBFqV4
BrlFlJjHVVzjaeaXmtHI7SirGDTuG5OTRHrUXv63oUsHcEAGaTnMJY9kEEho0w+0ZfkJiwi6SAk2
kkPWIQqbKaR/o1dyE/M634RHJHCEBC7FQLJ/t6WuFxTjbiRd+RX30RMV7YD/7j5zPY6a4rk2xnCi
TW5tHPlD8w0EC+sJ2EHwJpjbDtM0F3gY0AeROWQalXEWJaS++Pd+CnVkbn11LSZJoJuV2ZrcBV+i
YrlB45sH8KRjvF+nN6+wKWeTLKk5hYeOt8BVrVUF9FXcvfF2Z0wHLMSehAYioRuRjMUpRV+FhusF
V+2RdxUNOONyHDltk5zwm7C0CFHeg0AYy9AEqiwykYbQzHAZWBpjwAryAj1BvzapfOoMcxRQOGwm
l8AfgNvH3FvMI0hvlydW5GgxM9Go/0wRidPD0XVd8Sjz4zuaDo7faY7YeR1odDeIxghrkqq1OaYj
fBkmGG/uPJ0YeF29K2yB+GeT231/AmXN8E1ZlvNwHDJwQ5uAygchmt0WBMzS7XpN/Of33ubPhjjs
56EWOtRQzr0Bw37tw+fmkswDYAQx8PCuw0FJhRFJCu6Bj9v6YTUspfN37GE4s3EdQ4rp5fscmZyi
YwGc6l0Hix9g2Oo3Psg1zi86frT3/vR9epabxfWiGBaUlUdsdUNFYDD0YOXhyFnPcN3XnoaQW951
6XneZUVyP6DhDE0z0Kwx4htNc+RV5r+7rot6TYEK42B5u1vCtbtdTYbgsiSXa2Nt+zx7a7a1Oz+e
AD5qjGAaA77Un28FsD9DcSCsvR0EO8LZYdDoCKtTA7YOTUpDlbzZ1eVedMOoQBMqTKu/beHGMheW
u04mswHxIdQvv7sYaQS6BYCAD+DY7VN2+teqx2ypPHczq/SmYFTC54iAO5eLEVywy4mOM1rCMUaB
HXscdgLsvSo3p83fREIwZunGHUD7rke10TlOzVwtNAP7d6gLJiPj+x9i4Vm1HxXroi143OI/FyUV
TLukQU7oNn8UI93bdkzTHBOWKZ9b7gr0BNmZzo9Jdrw+7mKvjh4POYv68jxr1JnJmpUotGUhjl1l
+hPtowUYO8Ecis07zGssqkMdSvQ6V4bR98tIyb2Vpl0GgcCwsKVFl97mvde74jDXqeUYklEm+lpo
vnJ7zSlaNTjeGMLQwYfeaKoW77wN/Z9VQnn2ly9VD7VpkjUgG6HLujWImHwv05UkRkvYWU7bkwdh
Atx5lNtszfNGEgWBMJ+qn3JmHbPCAndef1rs3FMLm843Ksp3ZKfWKPC8PT92IJytzf+qbsoCNdKV
+2AZMzbTj2pJwW+a05aH9okIOC0PyfvkBnkOolNNWr3jdot0uII3txaOiDwJ9JPn8e1Cx8l+M2dX
TejCEAJ9bfdzbzb/MdjnkQdzcrxMBl/qpqwFBhu09AicBjcQea4Jbs+WBAe8qrXbg8SYBWbSNnkN
1oyDz7D7wUvL+azxaA0eQas1Ift+7odZ9t1Zwczknybrizns6VlfXhwFpWkm0ZEnuRp/96P/uT0K
safCbKTQD9c4wZtaU1oqBU+cJcNRoTiDG7lr6qIKuCsHUI+FzpAwgNM+337TTwFqueAZdUqtnzcg
G/p1AztQU+SarYx5cSh+ck2WZXAQqIL0strNBURKtj7pVZuG2IIklNxaBH9ezBLKYPWzj+e73Pjs
n96efmEXtmZ7KCo7be/Td6gp2fPt7muYX0M7lbCbegk00VWkUwuqaoyr9+fvu2KSNSigouUkwYft
n4DNMlVZxTxPOxOc0XMn/459VxJ3yReY6m0oZ3nY1vowYM8yJvjBzPsZJEZoJhIJzXq0JDujEgqv
p7wjwFN9zhgV75iAjxCTPm2sDhjtfyBIKAmVy2lGwzmGo2oLzY5bVzGDK9JDUdnDxWjvGcJg7W5H
6vbdDj9mw5GcLWAV7fGBoH1W2ycL297aunpTd3HSEu7qKID8h+nz09G8UHPHZaH7VU00YGhJ5Cq5
mdnpagyM3WBINGgvQm0HxzUrawMiOYypFLuHYSxkvHeNczwyiFmIT/OxaCU91xAabDcVqBu4CDsE
HkNoAVji84cEbp0i8/+p2PWLsHtuzOaZoYCKgoIaR7jY/WsZgSpDamx4UmUDXReG/IG+/qnMFJmQ
154492hF4Yr4z5ky4rGouQaG/j9RlDVfShp3KGSUY4lGWkaaJVWodlKbm4Olt5hFeuOwS0gg+ms6
lI1Uddau4UG5EieKyD37xNoDD/1pCpAygfaHecWrMAITWCxOuVZtsO/+//KyRsMrj3hbr1WhY8cn
L0H5QWhoy4f30cZMgjJ2cUKYilg3of5IGqR3EflMTlsHusSs/imdpXnOCNHxhaOW2SFfoVtohpXP
NV8efWrkxuqZvhB8XDHxVDVM0HIVX2fu/OpsZX0bDlNHYY9znnACVRtG9WzJcGMUqzuWqRj88r3Y
KTnIhLmPfJqx1hA7A2DpCaGOXaa/aBHlwik2H5RYSjwpU/5KZKZV2/zUQYzv+K8uceZMb0JYjauK
ez5yYcmK+jB6Jm5UCjLAzMLCkuU+kfCDDzOwiy11fUrcf84rBBciOubFjgjsUOlPC7Hvd2mTUUDo
wJrKHbFV+CzUHQZcTmRMDDHwsRmQ+UPE6mzc0C1pQ+8Jt2Vft0g5ye4XdcXdUQP2Empq6rZADhRk
TA9JCNfBjHyceXVBne8lHL9epYm47QKU4WWz3M4zJz3RbUuLM/JGOm//ZgqTQy/KzT7rFKYWQqqR
YJ4ex3FxAUTLpT83lh2ANJuaj/yuBndA4WOUiNVQttlRQdH0+oPgPTV1Ly6/TAC+GK1g4WB1C/pw
lidT3koA0xfhx6VSIf+n12OQg1LGfzdwNJzDaByL9A1TlRc0jTIw7XdTKCaOPgaTxnD8T3J/sosd
OVq+gKwYhumWi6lKek2Kk5y5jHEoO6lk7QqYz1v8v9/OvYvvfEkDbgcr9m6NFUYwt/eQbjvUPDm7
ArDEKF+pvR+DpXDv/g+z6qEXZeIreNknUiNGCKcsvhUJNUthxD5xkJ+oM3UJ3v77DP7Mo1+tOew3
OS4a0WaRkenkm6Fp/hcMqCVGdNkd5oXWvrM//4AXtXM9j/vmnC4JmV5wbm1cBY5Po55OD7oSIp48
03VNJ35TnR+LHiclNCgX7BNGbLyioGh1mTEvcHfFfkGfD+QaCFp3SrKHzXSyrLxxucv82z4K8v3Y
2bA4AzPQbx6r1JdhBPEGYZDVd2qnuHemeQXU1U4VwLhLXeFo00wFtmZjJ//lDtWNMqmjAqJ6cB/1
ryJvvRg3CLijIq+KWfN3hrb3huo28OY+nGoaHdFyNCl7dfdMZizHZ5/seS7Bh7j8C/XlYU9RCypj
pRJcVPfbepLPKrRnaqEKYomXw9EQ+AMe34v7l/k4xkTGSnn8kheMcW1OBH3yVLpxMneY+JyGIbP9
Ovx8wAMHau3w4aqlQfQ9ftrVdwmDcY2UJFILFgss5kVTsbg68Uocw3Pla2fXXWYKWsmaKNCiGO9W
KUWN8JlPx0RQ3xU9lCechJ/+xpTEMHCf68OYVQjiM6l1wryxR2G3A+EERb0GZa8vfGCPdJvu53jp
OIu+5JbaegBmAZYPylVQ8/gddSFqColkyKWqsrxo4fDOgEHhtvmOjqEXgwP3TIfvbanDoIK2nACT
HUfqYMCMLmpp5F9s3OJQdTC1sHFR238G5GNMGbJr/ZnTgsNOGh5ScoxN9aTRGFvMKluyeU9inS/d
LHdBdOg1Oby+tchDS7twGqlFnDGkG5/RHd3z9Gd57zQ9eBAtK2nq7++K99dUlIXAQqFXYBG/o9Iv
/L0pOkJGYgVOxi79y1ns1+mU3DkmJRtr7eXFEaqgdSxhMx4nqOv9QWjL1rRUVzHUWabBu1leFZS0
PbGOZWmL+6zS+G7tr7Wu9z1OukIhSeBje6ajDNxmsYTNFQDNDJxjz30+2i2+JclEvGZrVT5NklsT
ZujSS4+y8qW+r4bZaePpJhzpVaMRSBy3RmcryB+DM659FjB8BZ7M5ghOx4UQHFTD9dmn/EQezjhk
iZpIgDc57+8UruVIjrYBKCu4mhoF20us9PzmJ3UR4q9BZnyczXSZ4B5XzkN6xR6eXta3HdPQSEX9
hjFevDeKXVWx3QKFGROla/jfo9yGQqEZRBO9enVPLKfXTEitH6Z+hc5cuYO6M7mWMUqsw5DX/90S
QrrUsVJOJo/05ShX3vGGVgEcZzoc3R068X+7k1ScOlj1jarOv4OOCDn802j/enxZV2rq8LD+iEsC
2TI7bQWk8acgvN4R7QRJphNU9Au2Hu2gNuQb1ASgqOfYoW6pDMN0j18yTM5ksAngH9/J/cLz40iR
5wgjxvvJCokOqybcV9NLhI1h68hLaReFi51GyRVcXVeHFeJZ+G313OkE9L53mjEN0fDKsmPNB4mO
klwrNg3kceQCcglB8UYvW4AFmu4HftXwi3OISzhZHRdiOGb0ROdXsNk9gSUA5dbbdTpC0iwYbsnj
Wu1wFJHwQ3K5XQvMhecSlO8jCIcblDpyUY8wiOMOwlLjaGuTeOgJ+TQMwEazTrkrRtRZ5EtxCCob
DYmRdoF7nqloG1f/JVz0ifdBsuW3Fz6p1BmqC/FjFp2gveCcwZXFR+kyXg21/bHERWvAwYbo1i/k
1Hc2eaFmh/ZzlR53zUSXEWJuQ2N39u2v789iM7dz+SenkOqkis8SWLZUof6OZK+gCwBeHcz4Jsnm
pxwCMQ0KLVLG9uDUy8KxF0CMzXMhxh61i3Hdx1seZlh2+DK93+lFOWJbhFQJ8BNe1X3X/mgP0O9I
N5W6Hj+PQ/JUlPouksWPUORQ52ocdJfXNIvYRYqQ0bE1JBCin3z8/kRNNwZVm1wAWdjn51GwUy1h
v/hSDiVkhAQDrRlMLjoyUcDfCR45uSPTjAyTp3r5HXIGBlj+nBuSkBa4yK9RKp5krxUZXf7K0ESo
0vGSHYFwnZgzUOP2W1t0LOSf34b9keaqgJNKAebgUdsDWo4xzNErZzjjnP0fM/j2YLRusqQuYFon
E8kgDx0QrPCleRBN/zmtErx7XsYop4xeWImgWN829fb+uxtIhn0E58c1p/FSlw+4/MizvBuQujin
g0YlxDcIgzgF7bA40xO0ahcShvoFwxvwknefn0LXV+qY2JsfCxBEW2snuNsX6rLMgx2iFgLH4tuH
b9xuUzxwIXzZMOdLAXuCr+tiCaAPFdtP34WNBhGpNHNvWkl8w6X3UR3beF4qLtKSiO5TYXnH9ppr
2BEWEL3eNvObbrFBA9cjTtfLUoAz5E2Xtvv3Rdw0ENlP+7yWLAyWlbNUIbKRFQW2IlgUy4f43wR5
MTY9KL7jbAxIYPKgDDF3S9PRqoqqU3fZE4+A8iKs35umiX87JNTqTgHYK+T52hIM+gklOj8TC7Wt
2uZeZb5FmFLjBb/+qNTk3RSIb52aP7F++HSeD4gqP1ILdH9L6z2qmatO/W2E1M2IcovUaNkTwPZz
+F8FheXhQYmL3KGhpWtgKko5Nl0XkNhZt18mRb9kl6IO6pcKSP53JCbNy6ni+lHbxbUq4VO5/DMe
8pPw1nDT9u90GSqAh7y8+IkmPRrzYnE2UiM4G8Z/9rxB91FtLCpHb+5v80f8D7vXptpq9ey1mUvk
npVl32TelyPkAldC24dEgxe6Q4LJ3VvF5SFEuZki64Zeml0df++jQoWqBZ4d82k7oOqGlUom0ILb
P7v0Qx9IwgwZZ26Ag/O776GaoiOJmDKgz/9lmIJekhUWU+/+ylI4h4n92mUPCvF3T0H+gfHThE5A
e3Eh6FmLId88PTlVbmyXddPR28+WjuDXkYJRGKk3DnaUHbPa0gY0tjTbze2r08fXsUihQpds+5tO
gSNhcNo7uM3SJ7oEtSVPUl3heFIOBUEYepo1a06IsNag4cgiPG3eGm2v6TMWGhjUpJaTW35u00j5
nIGZM3S5UxnjXsSwgjvboMlUGyc2GaET4c+6Bmoi5SZHXe42N349G2cPQE/b5jUhaMIilyb3IzBD
8eJWX3Zw1JUWgA3SkNH/FZPYgw59AmGPvHqEhSqsMvkxIIJy1b1AdHlUKqF5oDZ+JOvNxVIBvQUm
kAFsapSTb7Baq/PtiecEO8acOXI21pMMzLr7K9dk4dQyfuOBAzebMwKzAQABTDPCLr+UKSFjAPck
/JbFA701Q8kaFc6v4UtUdx40QSnrN4bKrNzdiX/W/aMJO7JE8xaSICvCd8xluOP1vez/AfP98Mpj
P6r11tlWbDyLO4uLDYqW7HvRDVlDBC+Oxt1cedpmZiZp3I+qfenFOQ0w7jVL0xuNotTlWCkrLg1a
66+lnXm9Xz4QeQr63s3e/IvMxJzzJoJPHO9jobFT7YBxuVIvA57b/1Qe9v3IfWTr29WzaM0yYII7
aKHXs+KVu9RnS7dgQLrZyN5+zIVnxXuyED7OJM+4+/Wn73OMjUP6mQ9tIq2yzjpj98WFw0h1wzrY
/Gax9bIUuiVBuu7l3w6btIV0XK4UaHgZWnPjAKOs1IEjITtEQuhFo5M+GmEiNKmWUTWsYIYTCFBj
/Qdyf5g9wcoyo7kwzRW18vBtTIdXwwVZJvXS12/Duo1tOwX7gSg5kKlMU5J0z6mXhI1hniFMjIAH
6W0bLq1i783fZnn4M+rCHTRQ2vAkHzh6AiEZfi7MpLVn+RB+R7CMok4rIDwQie0IOjXFb79Iufjy
UvJ7BOg9QVcxAe46r4C8k3hyusfu7qS9piAFCDEz+BdknhmDWss3gZI6k2gqd9x6++IswPjha66g
4dRuFX2jSbKC/JIxp9hwjjN1imDQ8kpTtkowKcIVRwZHOI0QxD2hwHXAtOnqLgIt/VNZ5HszbIzF
RlKF+lIVOF1PBXTrrhcjPu/ix9a0lsoR1Djoz5groinrxUNwZqlSNXs3gWt0lQ9SH7ki9ox6sbj2
CSdaK7jKeMRRLLKMgdllgVL1z7eI4TF1cgHb/ocPHvzpgX+9XIIRw6xrTjtE4kkgz4qPRxtf7C8C
1Ri49eFEsxkpzusgwmM+WQ5FLI/AcHFnFS8UT6FbrVpkQWHJzjRd646yBVYMETaICGM6rd/zqKxu
js1G6yjpkuSsppLe10bDmrBxv6N7QQjup6ab645q3TjRcfTZCsb+r/zDsxaOzSGzuN2gAi4sUL0J
VGlKBfdcXO7PMw0zxvcGvXyw5gc/8bz1IVxZQMgIgzLevYhk/ZjdtbE9ZmIGmFbq1Vu5gFoM3H11
YVlkh6csM+eDT2IRol5RJu9BYV6ieMaso7dkXi4/qaCt3GQpbjRE+yIHJtXDEDs5guwe03xyD202
Cbr9Lubse/KzvYZc3thrEw+AHLdAnr0+JaYHl1f7JaaPQnXqBFwneSfBJblKs3DNtKMih7MBBO/c
j1aa+2y9WW0H0xjqt41D4omhO8x7rgUR1Fxc/xRFtcNoj79yEthu3QJwV65H0qvLS9CbEmk+sETl
GJHHZCzIfcdpwldBbfhH+SrrZESgcP6IpR2V8InFDGE6SUpdjuxUj0ArGYMx+x7/a/KMK+g2ZF1y
uzgghuQ/UpsI563UrBOntbGsenN5p5yoS9GQ2rkp+YprXN3Ejg4o1LPzHA0+NH0yMmEKs7bL8G1m
bB0WEUu/FoNaxltyLKE06tYlqYwyelXh7VYZm6a6Rtk6xc7UawEnoVL7cC4lqae+FhAP9/gjyk0U
lYm8Q0ZVKOh14tcAEwfqVTjqKfvgoYu+4cbnVj7iSrl/UcEHZaD1VWp97xuPSblG/bipyvHdlUzi
I+OWqi3YLFIm+w7aQwY0FTa7srRHsJDehwNrK17odz/8oGH3BXDfctycDJdJJuSJwNhmFBECivZN
F9w+wCJ54N+hZTDTUARrLoG16oAXp7mhAwKw5N+0fnuZXhyRycKrc5wL5U/75UEiI6LCmfkGL1CW
RkOWBpTpGt7Asr5HMgzFBu/VX8U8cbqCXI7Jle+R5jtyARJwUKbf7SC5HIXovnFLIAzP83zuwHfb
D2s3T1fjhHUtvugJaolrORYxXVQxpMR/QE+38PopqeOwcfvSzTvmUaR22jcK3pdUyoooUQtW4Mh+
sp3B9cglgnBoM8ECvOME1W5D4XDIT+0pXDpgkcJ58uPifg5FBGdr9aTIS2QWdVbkHgWmOXd4hUXO
qudGWiClLy+ecxbFjeZeLCJl19T2lQ6TEwqYqfZ26/oW4qTHQG3fI6FR8TG5VGMQfwy/jiX4cfp1
A5VxcZZlRFJuLwy1R4NTAWm4iDjPNNicFSAhDOGRT8jdevJ8tFmpswB9sEHjdr+wchtHBrXr5/eb
Vj8U7geVd5x4mpRE7PZ5gWOPIJydhZUqfWMwIY+y7pYpbfAplkKKYy2bg5fnv8WFoFIjhuwqH2OD
g/YhkVSmprMP1QX8yubnlC5Vyr903+mqnlQ5auMasBEHClhEEtbBOWVcusIeIDArvFdZUSuzb1SW
ybEXeg16wejfecuiACxzzL1zw9xa4P/QR49IIMb9sOCxjrLvGq1iy0avyAhk/OpQTFENFkt9eG8/
bXgKlDFDmkKr/oeeoA0ye3Ds9aBbSm9XWgdj1p+oy2CNtv8y2g1SpPHvZFxz9m5r23MDzVdMsYb+
1cvqUwSqpiFLLa2QChHf99idQn/cm332iDUNswipIJ9h3MBZhsKSlodDL1LTGThiiEUGDD8dUBFD
qYluks654H+d6GA9yAiTNC5YreSH9r2Y3cr9pO5hNur+T3GF4z9vtMQCTuU1PiH/6tGSPNryZL8Z
Ut+pR+qqOeMT7dK4TzAn9UtgoiOzFmdg64CZw22nrTCxilLZKFYEw1mQczuwTbiC1MGwWO5mxNYj
kS6zZfMmRj5LPcLTbXiOKJuAkHAIywnO4mJEFuUjtmRfLIsJYAaatWaRK/m0Ya3QrLT3i0dT0n4I
FbGe4oi+fwpveijcB+psa+CL3zC/fkJVZSEgIOzof/T0TVCSsuFR9AtpFxUS+jjG73ce/GEENvgf
R+GuXtplTCjN8Qx1En8z6TYs7vRYpvQh97za3TLhj/vR6VHuZkXKWdMgvhTEH9mDmASkWOWg7MbO
jeGl7ZltzlXNF4m6kduTPeUHuBHOV+pViB3Yz/m3dViUKO2GUtQBljKPH0Gx3fPfQTKBnCI4gRic
aDS7ZQWDdKGbmZIBTn0aVnK4WkXbVJA88NkTNukWid43B6bCCe233+V63DI4qbgPPHlc2ClBHYAF
VuhWNyvDVwiblIwsHf3t43y/gctwSbs/w46Q9BkkDq9MAQuhiwlz3r+h+HeXWZuDx0rwGdFe20GF
vLpP0L1SQYYKEeYkvSMUgaxwb89VFEov3wiZx33xeLs6iFSymHOrXO/CaEyXaGhD1gQdrgYLuQyD
y0Yi9se4DaSrc1crT0/w5ohE+gxR8zzcLZdlXe2b50FsQWbNw2uaqV3T7b34jzbqmnnkQCeDXGl/
0isvt6nhg48aNsO5+A5cP5bDM1+5cs2S+pgHj4gwJdlybA+McV32p4kDKfiiBKrvOawG8HvmXY7C
QydqCcxNUeQc/sa8KvFhhlaVszEsI9VuJ37brNacdK/A9ysRePPSBb+E751vtHVwcwCLb18qV6+P
zQIQuOH4XcmD9glirBvLYblGaCeuoK7HEi8Nt0P9bWvQ2/tfWOkdFCjlbpvg4cjTzNUbeMxYsHVF
W25Dz2kqB8ShOYhVqMw/73KUif/ksu6FLdlrjOdg0Nj3Cje00xyl2c6Ix8XDGQxYorI6IqrK9nvs
tX0QzWO62uQnNDd3bn5oP5J7cJjRML/c/SDHCZYUqc67d9q9BRlFbtopbJUhSOsXj7mUgu5yXgOU
LncJiVqk2QH4TfOd/zVxSksq/RGQG5iEoZ/6x/NK1bsWydJ+uZ1aIBbavKr7cgxJI4qRj2Um8r9T
5co79LfDkWH5DuUn1T5O4NirfLbCCWiCTtSQdfIhJuUQedd8tkzaQUR3tKyD3qLjKtoJD4EIQU3T
oPf3qqnQ/CMdnkgRAQpqRGWqfA+kL4xJGPYSf0GnUUFCXQkfoc6V0qyuTNtnN8G4cOgmLhjGdyT/
0kSEUfZn3Zpxf+BwKfo3KUqXAQaOKno2ilizkypMZM9LOJWCZrrIMYO8wHRbsonZVbCK91siaKDq
KOFl2qkask+2Ew1jW1HGlFysBrT75eyy4jRH+Jqe2VBpVbMayBdPmZUApmydsUBSGq3qOG4sfhJf
YjmBJhIUp8VfTQQGEB0QSPnCZIKHTkx6b6dp4J/xElF9r+ZakjE/chxhHuwu3K/Lz40Fs1x/jpgo
8SeijZnlUZWUSPmOSzvom+OWWOE1L0BrUDjYAPYJQe95Cigw4zGhuxjs3vgsdBYhGzlBYwYKCCvX
xq8W9s/X9bZLzjhb9m2U5lLcqWfvs/HDQBsp7eNJPdbfU7L+5z9WWYfKme/bZUPRdadsQRlZhFaq
MdglTbWvERZtcmF1di+vVBbepVJ7BXgQ9gI07TccCUlkd5TMnHW9JFh1woHsKoYnAMJ5vk2+gSgP
1/Co1a1IfymW9iS3e8Zh6eS4/k+HNvBKb2wJup6Knm0qaB8xKkGlsBmeHbtLS+Y9a2DbZIjJ3mdY
ELGernHBfJtCg1O9D9+AOpYsOxBTuS3FUkIu/JVKXpR4dQwEIKAMEXmd7XU4sqxkk+C0zBxqFp9k
Uk5Uwol/dRUoq9tnNJNm2WVdbinin/E9Enz+2USMfmYXcFv+HHKy13iPUyZLbsk1pKEdNCN7RiLV
jKkOkyOxDjXY1eZEHWU9GEwEZHCsFh8ekh2RvZRHKNULjSUIfFQ7bOrj2MeBwiyyCRUtf+liaJss
iVNAs1ONfypqqZ5l7A9m/pEaKQigPIYPmIYafhwsa32dylSBMci1uYUS1HzmjDaUJwZ60w733fFs
v2obZvGB9XE/Z7emLex5EcuJrLBvtQqrfPRfHohTT+zeza9ovENLyHQAXfJxIcnECZ3/Yvco+C0C
WYA74c/RLqBeT4ZxqsU6OJZeJ5OolTxS+cfAtH9Em/m/R0JrB9EK3ECrDYaZQwR2Xgdx6Ux0/6F2
vIsi3frlvRXkf7CSgiw/lelwycvLK6TABaNkRaLTRdHfy8KyK/ryBx+oNj162gEtWzehUFA4ZNF5
HNT4HIAWviVobOYMTAvp5BG+3ttCA8ymGbeYWHTDL20DNFQnbRBfQNXTZwfRgH7qg8X8jd3WztDH
RO+wPbo/weQhQp3E+gVTjyneioZMa39EqHofkJwrY3KjoLTjSi5XCSwCWGsqgHXCyacWh+9trSX6
4ihwzfWpyDBWDjH8JHgngLgSQDYm1lbQdPWFihGoWfijs9PeP3WlBgxWbj4PEI4SofTFUA7g1nNB
tLkbYXauUM79v0i7cKIjbBN++zNY6kj0jMOBVzm5A9PB811ggbr8pn/s0ZYO+vKJXqCkz/vhNZT5
rw8I1nySOPqiYSj8HIjMyT6jvfwWtZ3dGCcVTStGQDlSsviH2fiw6XOGQmFHOCJzeE5ldixBcN3B
E1fliiOiQzQdSyMm11sLgWzXM8crOFaFMltnraZAs9DM1B0PIv+lRUBPZITRFVudhzo7ZbIRY+TM
GVHs4JNmx+/bolankre0Bl1tBaMLkhhCBAwYomgla5G1lzVefR25XLLeF3mipqfS3gjW33bgoH5E
IKuIbACW717XqjiG87IkDfs3c3J1VJXdBwlgKickp/fsiLgYL7egtKm5CbRGidE4QzxBtUOrGfas
SqJ/3UxVe7oGXn4iVgOVdb20DvBvnOKLdDDLiPkjFpK0GS5Su/kO2nTBSVDPAe9tFFzsKyFPFnlM
GO2A/2EyqLtBSj4CvepDvBYFp9iKTgh0AYz75AOECAiVTgjMNzt3qn6yyMxD+DfOmKeX7ODFKl2+
S9SN/E/qR2YoqtqXM0Dv5abl/wuVO9bZSnIeNIgrROp7oCKQ4s80m8PsI18B9IH95f136S8Nh6Xf
sDoopvYLpOTCOo3Va0giU6Sdr4E34hgeOKQHw2Ei/TraVOBSB1ZOb1ipbip8XDA84XFxRhAks6uE
MEzXRz9yoFLD9uq2KVopxZYgZ4iIGG3vEsVqI7f26caGnPGKSS2mvwZPh+VRtLPVM3+So8eo4bfT
M5BfwCbM7sprGXuQS5++zvAUchK8gl8roCvYq7AcqNpBrkfAHzhY4eIdcZc00D0+1LssXl7Z1S3k
0hQ8gsCsLpl8rG6xIWC5HVJm/VvFmnmxOxXFK0KkXcQU6TU+zwdE8c8lvocZc/YaBxHF59DJXAz4
7v3UMRcETyvcm5rF0RGGKjKkfvNpPtslhEK+f5xHnPzINoN9nyxilXHNc5Hm6IA27UFT2m3iXxD1
bR0+j5P8VmtrvYcz4BfTWBoudpMCqjpGQyb/wqcV6x8X7lbdfv/HZvpRNIqtZ817MJFchCxftSAo
+Om1hJtxG0rlWblYPpes4cDQDIHWsbwGph6oA5jeKXtrPUsa7P2A8VUMaMrRKIE2WZTMBb0PwsZS
kDVfQ/w23+dWWRp5lX0Q0FjYwFjwU2NpstBHCyPsdAEkcuQ53lbLGKEaByVm8AUyc4GeNJgzsSd3
vVbqDDepSKWdqfj6BxiQ+xrE90cuQqKhUFupTH3kdVexDZhznN013G7qc/rRMldgWmiT5EK1aLxP
arDPVdwfDoyYvwStsBG5UgMhq2tRtfcohptSmeRImLlQrBfX6fzQky9BDErOcK2gRvDo9uHMK9kF
MTMBzCLsxHz9BGe9Yuyb5zIzttWxCZbLVTpIgDgTZkUnOm+lIQPhRmlgUX+w4cfEP3Z+3VwW4PFV
FEUlWrDZfuI3nWvQPOkLfJyvfJLlSkk0GpRcTxazJtnvZ4Gb4bKIIQxzOJ5mdkuOlRMErGadxoDR
uUx2HcqppWVE0nZXP+MireCQt2WtGP9dP6M1+BHuuHL0knorRyxg2UEpGZYtvwq/+J8OkbluRaGR
AzgY7+3iWr5whzRmXgSZGj1KU79G2ID+EQmLzu74jDb3KHCsJpQcZOCfvXXm+ewzctelQeWpoSET
n2krS3h97XcryDo/+Ph7Kc6r88C2i4rl1mYWJizxuEC8jJeo+9TKXjSIWXnm9UXEKjj1BLvbHTFv
vL77zxqHBpYNhtef0gkCm9ICEeMkLb8TY0dwz8niWM8Aw85pSlo03TVDR/FY3zm4+Z5lrtIkZMr2
PHEL79zc0p7T450ksTqifHF4FTf/W+PhV72yTil6BnCjSOlQODHD2/vG2deGnK1yuHxJLEMocVnV
fmm737UcPuFOQKMtS5IGxo3Hs7hUjCyUsOgPfB22s9IKeNeJBpU20b+wWBLJrffTc0aLGkeddeSf
0HvMnODLP8UyE6GbOM4Ih8eni+UZ6+ppo6KSu8p16FpB4Zw8bobGIzPRJ3gYc5hiPUhiEiw+ZJ4s
tAe7oBxY5FSOoa7KX63ZctietN314gqMQraWVP5TsZG0qfGuO5NgbBo45qvCB9chH9xY5bQOizWV
qFP5nLSHa32pt9uBlIvWV4m197Y7TM1ZpyumnfDdhkWJ+rS/RsMre7vl+Pz8K18BStPwwFetk1sS
9M41owxJX4hoay997sO7lq2tuh+6AtRRRafk7+mH2KwbQ8Y5S0ew0J6tuwwyWpk8l6S7GX8XeG0r
QYqMlKMjjXFQ3iR7bJGPuTBIGLxrkUmX2fCVdhjtRjY6xBBGL9O9Fbw0EcORzteCOKWhoBe4KrW1
qs3o9DVnjf8YYWd9pOai41E3I7mozU3aUXNkWUhIPJ3HZbv2FJolF60aFeGIcScZ58qtREwHjPj7
HBNxXVSgV06Ua/Eau7b2k2Qv6WfhvMVfpiCPotEFDsytl4dk4n7vFiFA+VBm23w2osn+0ycQu2Wv
aXsxy/p/N5K3UMl8V1c5/zBkJ/e3OVTYJDs1laqEworUFdps9vWjO2YE3FuAsJnDWw8S8uZFB5Vz
4MiEDIX5oXdQF+WCGXgtE7IAeUl/77hobw8kzWfqNYlhjNgekn3YgbRgqNaMIVJYEyEUMX5TJ6C9
kb3T1iS7vvw1M1E8e5tP7E+MulBh+m94iO8aWw0bzPJ7ygPv4ShYKnCMoN0XJOLQ27fSv45LzYBj
9Z2Bcj9X2vL+z0NzbI4gNj6msgk4ORpkD/KbwLmuCO/PblQvyGeSFTLxKNybB0ozis3o9GRwoWUg
QzMgrXKreRHDJ9Ni/k2DX7+gWGe4eTF+mUP+45Ef/Z2+WaVWcwPyH8KGu0jhEHASmGm/TQYvGEUS
0gsRr0K1qNgxV3g93cg6mSYpQsT6qTd0LMImlkz+qYX1e9S4yhb4Eq27M4+MD6mBFTiXoSPQKDOX
aVOo5bLLqthrG5IkPORbzL+iwJCEw+yrtQGCbOQoLmuUPytv44e1CU5hUphToxVRxvE7ID/meuX9
RCR0Gnk/JPAy0w0l2j5gB9vCX3wYx/nOd5zJILUEO51n9i3xNT620h4qT/Svi5OOytmGio5KSf6T
+yi71C1XgDUSnubaDZ1oJZ1f2zmNv0AQjnhbtp+t+Vq7Ly+AvKfhJYSkTIrYoWPerBv4bD4nVOAv
nElad3gszt76VBwOytpVV8J/t/98M2G5/Vs7ZST0k0hVNq4IqVTEVc3rPUla7l5+slZprYvDIRsi
IWxr/vvU2XNuedEwiMpBs2NU/u+rUJhLF5m78dIOCi+P+bRA5+mZKTTclYddwR+zRm511aJwr1OG
ekYJW8ODsedoos54ccJ4MZ2OQn3Noz3/mfHXuh0I613FsnRqsSpA+eBAGOMIBA3/EdCIddcDSXJ2
9+vB3KRPy/vOE+/PNfooOmmu1qfzHkT7dypZmQHNyPRHQDocFC36x9pqEdrByMtLkrudsk0G/Ial
OXNZ7/OhX3hQeHi/Ob0v+sM9ln8nCiIfsuc9nSiSJdd6ut5DjMqvsm5DngFVey+sRRGRGX4Oo/Yr
efQtroEMF/umFD4pAt5J4gAvWF2NKYDRbGJE7B2d1EfLZaIFsFPqqxqkWzu6ZDp3OMmKXHsPLQqh
xnPdcl8+DrbbABBLWUZA/rdQ9HVR5S7zaydtMbCBy3KSLNavTn/FZ9u0TIbV2jAKY047aq8ylZLe
duiie6nU/pikrTQZz7ajxmqhUhtJBngvn6QWHg/HwMEynmQAQr/4lOhnYwYavueXDQi/L54+PZ6Q
hZqkldBY42u6yFs0uvAsn8jU3KYIcNCoMDSSujIkZ7FDI6PzURGIvUWcDymrVyN1DqN9oX9Zb89e
fKRfFyJiexie6LxNdN/pGvRQIPcDtoUpaTNlDOX9r8QXgwDdn/3wkHFR74xSz8zLKfm9XDYpxOpD
XktmqDkLXEOQcq8Pgv4w7uH7Hu8K5JrxwQhtHd8JP5B2c6ZXVmDEcssSY0jIujvZ+MobWa2v/5aX
cpTycITl+wIKTlDVMDWeQgicFRrRHTrLqinX2D/NX9j5AfxUvGx1XaWDBNa+IPV7O+3Ywv5TGX2V
1Z88LW4auvn2eAhvLoeEWjoSLB44XRkT1wWPIsuauxk52Ewpmmigs40f7Wb7aqmVIdxkdvoJKREx
vb97YgXT30DxOS4xGgUFMysxCyT9PEwHDql+2JXLxA1HM3F7yHvs6+yYerDEohLEvDSCL8sXqYv2
p258SKdYQqRdu5dOyrPJRg8B4P2/c85ejhVADBEep8xoBkd0PsiEsHXS5nMt5rTC+07FnsMTI8H1
l8r3r3WRxyj9SgPHh6NQ20EoBT73ThvWeAMdmCLJk5zIX3mHWN+kx3tArNHsIcPVG61jrojm5ht3
L3J8OWIGn8vEsch0pMDFJ4AkQzhmTKPvY5O3T3BdBdVGnQZkXwMD29/GsRtAM7s8N5mPS/6skf99
FySYqh57fIenSEU77Nb14rlADh1o64geWCh47uSqL3gjspuO5/qKY2W2BImtFWFue4p09CE02362
Y4E5SR1kCBT9XDxe2YWTttQ1fXbVITxnzvPOMEFDAWChll86vfC0VShkNoes3tdSjKe+fHw4PGfP
XCJ5b3B0X495t3iWFFvUVNv3rtxgqe1/Wb+lhtwuV75K2/dfOR9wIwdXGu4bgG/JdrgalLRhZCYS
Isllmq3NENZh/lGYB9dc5JrkwiFjnYkiDl7B8ruGgH11ko389sx/H7wvxcjNqJ7nf1hkRxKBtzoR
+N5nfA+FGl9GkEMF84aYBAnhCU4eogETnoYaVxpoI6fWyJJeX/JUvDNnsh7DeIPixtp1D2b+FSQX
t/HvMIv1hyXhpmP1mxYBK8RH6f0dGKQ4dyQwn1RYje9jWYpzc6E9SxLovLskTAyEcmNSemtXFJgX
bQZwgMcfK7aZ6bYbfMkCY6NZQ3qzCRN6E41qm0ONuYlQz2ZQnLcpVdtso2na5DQoWzFMGWIQRULf
NxlDZ+2gAnRMIRCnldqytEE6vlcUUzgAfw68pJXSVFjXuFLQ6/7gjSc1EiGZQsVAH+rsfXyWr+Z3
OgEHf0v9hUfd+SP492bhZ2h411tj4ulkiaBvBZIKAEaQFpXDrV78ABgNrAAdtnSHoNCQ/90ipLfj
uzq55kgL+/+kkr82xp5SbG/fs0Bovla8XlvW+LNMbthdAeWo6cGWwWdpogWuz/f4EwMdG+XMLrtN
AscyLLUhEcscSZeP5uf5uoZF9L7LnqTrQ155WKpXwpP2HV+8ojEI4ZxosE6TgEv/TCXsmsURqLmB
YBVgYc7GHO0+mensa4ZIyQjrSjaq5PvCTY2qtlUbHj4aOhZZ9bpkInzVcGqxPaUrWDjhspU86Pm+
sck5oOPmb7mGvdCEIkX4zA8DrSQarn6cg76PgIS6/OkJXxkwFCeVWoFm8mBTGpJj/IG4QeZqUiem
4KNdIltEP5GxrVsak0CeANhiv4UOl6IVH2S6fnKBzBXHibFnHOj22ZJ7+2l2OHcezPeCgsqA9qRQ
dC/HF7sdKI53HSnC+4ukZb9nKezXRKbPheiPLtFt0ejSR1xS9XJ2v3aEpqLpVp4Q8FNdPX0Sh8gs
ggIUgVXJd8QlpWEvvhpNNrwByOtADmG9qCXCyQq5n1YE5j+YpxHAiRcYJwXLNZG3iWS8jLrXB49P
JIbd+/0wks7qOq/aqCVWfcTR/X2m5hEKTHu/V7Rc3icg60cQHeik6O1yB9H8gcJUPt4g6pMxy15p
+e/vrLMpWL2VV1jeL8mfFvq3IFOjfj68sJGGTeFSC2a2SG1CDyIQppFJPs/2sWeYli0E3F3j9q1X
mhw2dmpm6oZgoKgLOYLgvEMK/GnGeiAOISOsPEA5GWxb+oM2AvyWR41PeFCpDE2bhlzbzosTS82M
PhO90tDVhlLKRy41XjWNWGdHHKR85TBbYqHVf69NPhuj3U/VfxKesiVQisrBRXwtFpJnPfI9EyXT
AqPxEb0UxP+54mJY/9B21mflm3smj1YhBs7ZKhvjV90/LlmotrQr5rRLGu7LKcXTEFStL0HzDTx7
bD7mtEz7XX9CUBUezlP7/Qlob3WGe5zmnojWCNZeOqLMO3Bn0KLuJciDP9kgpBnaXxdjBkQ0GZrl
XOpAklW5vtrJTwDzUI6w12LjXalXkFQXxqcvKxpO+3OMVqjAYpNdUQ/lh13jfKV+iKvmhr9+ugr6
chOxZcNEwA7rwAu7yPo06HXIEqfcbYcFmwPQC6IEaoISOeH2SE3IkGEpDiGqibLPTns78CHH+BUT
UOHg5moen+bqXfTJkhpLlkTr3ESEgvyyV8L0PuXFBZL1VCrk2gmBRepO/XLpNYzuiO6iCADLUuiV
Qv7FMn6yqTnYto8OghW+I4wrSS3qX/VZ9R9xsMNdTo4HzUYbsYMn6NoG9vi1gVE31sUgK+aZz7qt
dlOJjA9GsGklvOYjOkVhknfQ2h/ahbhyVxUwhmpf/KOsz40HHnX0SuWv43jMVad+eNeiAFztfP4K
AYPuJie0ixvrXiQuWyTByD5QdCxyen2CZ+uLb6K3yi5YCNAGFTUxE2wS3L8tghsEiWLjhyDMXYbN
JiaC6ACDTAU9jR8AwqNuv6cbyLxSPCMRQ5N4fMXF1qbKlwt/4FVJOR5BpNouQPbG7AAx3PwdkID+
mc98hk7yUWFH+hCWp4Ef5SvHs0lRQtv4BWnQRj3T1mTVr2dcy56kMm0KDELiVcMZXiMlRGM9hPSe
MFYl+/Rw4hzSZv7swzmAVGK9cfcKN9Vt2ejgpNzk6F0DQ3wcPW/7d3CW2WkY1VimlmIFXxIVMnTw
Qp1m9VrV1cTuOCh/QxjPjkhKusbYY/fBti4dtVt4BgnwsEsLdQiVn2kNm3t+Ku1WVOacjjEhC7aG
U1vXxNqr6C12meWn5LwCECoJX2WBekr8ARBr6sX3Twf4s2BQyfahFNUekY80mR4WDpkkXWC9S8nm
DkKCnvR8qsgezI2C+x7alAIJvEEdCd5te0wRlEsc9H3so96LzBVQCb9Wc8GPiViYdhyOVLAOyVDE
Hhm8kXzujlm3HsSFKfa4GTq1gqapmW0nMHIwsHM2iZQoBRUK16ce7jaALTnFipAi40V+e6e49LWD
dgWW/W88P4fGE24wMH0UN+sR1eUqeFZ14QBuiLP32IraZ0fOQIaorjGnFq8OfG1QBLzZbLbAcgw3
teLhPC7lsp9ZPyG4S9d8HPNJqN+0yJPbTtMlSWa7q6WX1JMNvUS8tAna1fCN/bwJKAdZTPPkxiCL
JQwInijqsMhMVvZY2kC8ECtHYBXYG36dURVePUbERnj2bO6bzx/R2fomMix4S27Vd9JwjxPmW9wY
FE5ZNYFjV+PbdWWaAH5/Pr0gDtgAUTxjrOYvVgnSilTz/DcPzfjdKe+i9VdYuMLIc9YaRayRmiGI
FqzDPaaAMang6TF3F63mLyGzaobPYYVOTsX15Qc0bLEIGxdPelFDBaZyDXLdUl4TxntIge5hRACW
OAf2n/hkrGLMQ3uZsxZnnTU3zCURGZDVRpJThrcO+2TsKYaQy0qEGaOzPCMJz7aHDMGyyL3Tgegx
Z297Vghu+xkFt3AkCJyaAFyYDr3geIKDh3KA1TmJOiRrCo/PChKpWay0/rFPcjL/+b+HARjgi+Bd
eNSzzNOr+qhpUjQ5tiqJz+iG4+mzU1xyUJwerM6TGeXvcRNCMx1QND4lvUwK3OdR53DZkXcXILv/
hqaBVFZVn/9/tBTS1xJSfRf16YufhXOaC6nKEr+/ClogDW2GQVFAXwOIAoDDjnKVz/J+V/0p5VMw
n5BxR5gyrPPQzgySDoDSS3fvRYjweSzfDdteclJsUtqDWGmRadeBNvCXKfEye/ACLPiSNOFBRckf
u2cI1QeN6fPqf+itpR6f5MznWKl5JVhkxoRkjLrb7DtYky+ADp2eAk0UPeo3iAfSjXSXbBP1fscm
YJaB5kXbcSEm6/f+XOzwpy2pDMpsdKgfSrspt1aGGd7n6P7LNfrVe1y/BAxaxOcAtUDg++VoLZ3c
Ev3UqScmTaJNQEHw4Nb2pU22zLo/PNHNBo5S8rJS562JUsgPFyDu1+jcMVu1C9MseUAkshUdCDCq
nVgCWkUI0YhgwntwKu9eVZvUM5cL53HRmGcXOLcBljLyQZJZQNZ3qE1CrNxuFi1dZ9bqcmsoGHIf
rEr9tcofETDbRKBnm4PzBAPBDEeYlS2Auf9k4AXJGc4c3zxF6pwPnD2TikJkFDLFUN5WdkFSXYY4
omrZjMLmEqE/26TOXNq+NOusxZOQMkynaAm9188Xm0BtqdXWXvVmPgd8o+VrtMypw5cpyW5/mEFO
WEDhh8xark6DcC5B0uP4HiXhlvdlZ4F4cN1MO2zyPxKpUpMA+0LYhr/gHbCb8PV40GyY6yiOn2Gk
F9IuSWYk77unG0Dxz+b1aiRJ9MLE5p41FTjngMNd/7JruGX6TXmegg19IpLj4JuhHbemGaJd6HFE
Idd85jK3p0XQj0u+ahAUGA7f1dRQapoPvTrxzGKz3878C6ekfiSYLYWbAdC/WsU1s7U6kCWuhTPG
Hbc+eFB9nPML2YgalseMPQ2vifbLPcFPvIIyUsB4kRH7cO98hGj5y2QGWGb9n4j/VK49gYREHICj
AdMBK5Dons4w+8pHe6rv3dXzxInd81aOagsW+0rKH4Hk/UBvTYFmxObbKMSmzuthkTvZeed2FjIX
kflaAi06tsvx4znR7JzfO0b6dDEDy8lVGN9gTAZ0/ys6HTrLAJtELld/Z2HPcXwMHUK+z7DxwLc8
bR4Z3GvFCYKpmCN53OZDfnG/dGqNUMycAlB0CiUKnDDFt1cluye5uK9N1iyW9BIBPrmQjocmFNXj
awv8YZ8nkz4rtxIad5+Kyl1xsbhbufsFK+zelguYu/M1gfPziDUWfW6+aGQ/o6W6B5aHbwduX7ub
pt8FtmRhtfQlqHHVVZB5w7Bd4GUrwhvGNhl7fKh4kje39xaEpLA1qYibprxa7nh4h6M4FqD79sxj
hw5J8a0gr3cio8Hh3zDWAH0PYkuJfLT475a9Q0CgIdr18qLh6Bs0+HfXh8uaN47hbw4rebAN+Eox
RqDEelXsAK4yZQ4LyATTgOTar+a6wRdGqZ3h9cbnKIJxA2X+X3vTjge5d2js+xdY/wl+EjyDN5us
cW2SLhI3XFVVLiXYjzHhV+m/x9Ss0w4GLIgu287BSutwMjxSLADjIW17yPgTxzpXTo4WTy1gsVJK
qcJUyd9B6Kzghu++lS3MVDwLdrN0u/KZsdwrVZ66lqFSbPNrGSViFQ38JyNWEgNuRVcVcvbfKV6C
xKpZIg80Pm/s4Io8ebHgEeDuYR9SqkJ5YJHPgUdLEaNSFhDe/CrJt9hkpHB82eHDdtRlEh+YhAC3
v2e0mD2E0yMJ8qDK16uAm4Ijgj/wc4UJ5DuV0Hl84OFGW+RVBSntz3IkXH3heFopAbVDM6BYbIO1
yo0AU4PAYIfW8UWV4ChPOCvgc1dH05cBUpcKqigUZvwIWnS9wlPW8mwkEc8zl5E303odrtSPVd+A
ZlqrrypQNGdrlsBf0ABzH/mTJZM4rvvgLIRvfyVr2E0ak0UK+gb24OzPPmVQJJypOlj8xI9EZx3c
5tsbE8tU4+kxm7an3sRTDYrZ0xadessogWnWXp03JOZ+7JFJgt6I8waBO8ukLWsv7GvhE79WsS8G
nO1tvfAXwvjxIoDWLrgHVEYWF7NQpbkxa6WO8jHNCByikyIbq4rwR4Lj7rjo1BhQIWzm5cZrHyTF
ClxXlmKBQvyrOCuShrWMKU5FwKZsFQRwAUANZZv9ZgSfLNQfOidf0ty3+JFxiFHRXPnKAhrxmdXX
eRVXPNl5pt8owsFU5Iihiy9yHQ9v22GZXLQ4D/4O73So32aaJK/BiIO03zchUY81TDEZuAABEd1c
rkCo62KI6Ks0GFIKfJ9zr7ASWyymXTltzWYu3/k1pJB8ij5G62lvRg4asH6VqGkZHCpk8eDOpXbZ
YBvsTB6HZkCcgJHUbejXWG0f/EkAumJYnPoB8jQ0zH2emQ7NkTdX2AgNEcolmyHpxXS5uZzAKfsJ
DmGVPpBjUTB9V5UPZneN8VPOfr2IyR+9+qRtL8d/45tgIBAGuP/0CqNoosN+AKAzJJkvL3u5rFHq
wTO76SldChDY9CkTxDve5nlAVru1c8wpC0trQ5xx6Sk8/zjy6KVMq1l9wS5DxR3EbBLgZz9M2px1
lBZHf9CXEy7FrggFDGF8vxquwvsDdJZRT7zTtGWi0MLPGcsqMH8zgSbMUpvju7TUcIjMAXLpT7Kp
TNCGA2GN5j+0jt8K9z34t4qYYFRcRgadin7IV8GFvFV1Bdl1LZVpVfH68uk3/djXejswJxwKTWVb
sgzTexwFVTZ8B623jmq8kWRlz47V9Q7tA98a46LWtu57pqkia7sZd0yZWOItKKIx6dTv3B0ltcu5
LkrVPWbYDz/y7O8DAKA2/E8qv4zUI7ViMdvkUCTlLPbf342uA3+0sy77bAMiD9x5nBAAH3wxUsYp
oVVAnY11J0Ij5awdpFAmPr4YHb6v/M5Rf+4LlEtOOrN5cHn1rc0364/zUkpUmqkpLN3Sa43Zin+V
XyiinkYbmqB1eHRDiuMKxpKMyI6ikcdrIS0iqccRys9FLOKtpY1WcF+6xasxoMmoZFlqAloV39xF
8iBvCIs6mCVBaPrf5AtHExxsNjuht7PEX2vINSWK0qwbq9nToAayCFPluOglUYdbF98RVr2Lptd0
rSCIbpC9IH1jAWm2Lj2Eez4n6ML7ah5zehMuJMdgQNmZIaQVFnfZaVmI3QgEHWxKwyOnnvw/R7gv
LPl7xw4Xrd3eeaPUocFp9xaZW5V5P3sSWhLAuGH7wHXd7eSos5j1PRgG15/TX3CZBv9/a7+p0uZK
wzc11oPgGAnGdSzU303zW3IsBWvk3jDewTL8tKZ8aAM0gB1TVOnnom0WlAtH43Lyjj6xuI/ZtObs
pnYEaz+xZ+CWRNAMJqmiqy1JipisLW4Hl15Crh55sVF4wI+qC/Nygsrbd15wIw0S88J4n20E7ddc
QJxS1mcDM5lYwhb29LHhIBoVl22AxmfYBdRVd1ncPQUZs3sQzedHBAKfv9rMX+kDV3S5CUouhQyu
BPVoj/AjxkmTPV2VwuWQLriHPszFpqKKEPZcaZIhZQLtzpGWz6H2HQwi7UWTyTG8CX+/7rjyhDdP
pOdSOnoeYHOFq2D3tjxe4MY17EH5BhUgqkTI+jBnfnEMAWh20AwCHMZi6AEryWITolNBj2YT4auJ
C6HCAM8tpojxVZYV3LtZGOhsLrm+0u6jpyinY1S1YFX6v17YTtf9+8fjxiecWZGodW/rFsk48N3S
hbycCjrDduCJyI9nP6XwGqQZHLGMM0W2X19E+zWYg5QxcjyxxAOstTpDpXdLQBzsgQLqihnSnaN2
w4CJGdrhNO1TvWLXRQLqVkP0BcAxOX2b5qP3ZVZeW2ZRDob1FNTiLcS/vWcpMUckqvWKehlnI7k7
bK5sB9+2IMr/ngobR1a/irITZ1+OrkbS1E6gbuGWXvrurlsjUP5BleiBzPxzpQroSrl7eYJbgOlq
rkXLyCITRWGlJtUAJuTqLH4e4Ndk+9UB5IClQcKDHWuoe17lp93jvvZTpB8FlsFbTZh7kQP95oCc
YBT6FeX8azCdsxNbkb26DtNkI2sWmgDvP6gHEqM0oXMdTIt4SMQd2JOZf5C8iHUKrt9LswQ01I6N
Rsm8wRAnma6qiC2QonQbPROOiQK1aIyGG0zXyk0C+W+r8BNp9JdkKaMwDF52swkuwkeT6Vo64nYU
ThzzNqkNEocZ7N+ZJBwXBWGI28vAov2lbhLv4DVdhXHUy3wJoSRrPrL1f+nthtPHf7ZzPmgjOXXN
3QQ7vy6GQ8/ieFtIRFbISpzw1lu3HeL4ByvYq3aNaIcDA0S2dptHG7AWhGim7+QU5165wS1dS6dU
kEqYJQZevX8LDeSRjx0pDgSRMOFxdviwt3xRCck+vx3bs0Q3VGUrWYxPhYt5wQS1uHpSwcMbH6Nu
WPORH12BBUK+Cns9FH5xWolk40niQPpLfNKK3DuL0egYdQA8dw8RStTo0BC9+o6rlEHrjbXrwZh0
dgMlTSuT2Lyga1Esfbk1TeEIIveGI8MP0EZtqXqcHEM5/dArAW3un1N2G+SKCHT87WjfG99m8k1b
W2nEnD7ZQlaFKr2qwFrNe668ABkgLQ7NGlJe4lQ/V675YJYMKmuUgQ8meILDqIvfmhN9vu3LY+Tk
4+bz3c8iO79hGkm7+qZHGTKNCNz7IajsNdg4P3subjqsNK9ZKEtiVRYy7q9UpmjgXJApBAIA4yJR
11q5q9vVHrhD+y5112qQi4QnV3DzzgrR+Xs/AjZKc0eHTmWLIupfV1FqkVZdS0fdQHrtnqUFjR/D
Q5g2RjClzNmRW0bdwIH0gcudxzZePsxHPEU83Q3zaB5GjI0N7BdrnYgi8ypzFn7uYgkw7om7mUTa
lhxLqtjJUsLUlTGAN6PmJJQb3gAt0U/Ipunys+3jGLgfZ9k0avqK+dOsQ0LGVZS4WeaSyizWsLea
Ut9KhsFp0L8MVDhd5/cQTKnJLNvO3l7yl072XL1rT1RExH8aWAfcZCnWbjWnfDcfPjVdOutd17y/
g2GjJYekAc0PAPmqXDlQI8gqE3wb/tW8f6R/PvyVibpXgBa6UD14oUtnxvGNOxUHPl43cqlCoKwy
ED8W2CnevZZ1tGO9iDEvDCAVkhFB/SS4gJ9aTGr9GOyF9+IOVLoDmAYlhOdtJBqOntC8Xv3DSX60
KHNYZrHFBBG/GXZ0pEQmFatAhdwPNjHjxrI8LwheMREmZgupEuU61iMSxIPm64e2TyRNWXGwBY23
TbCm+EAFqI8hJUoVHXsAVo49WUl21bLWsIU74n8fgErolUTJQMyqXApqRS0BZ2SAgSOnzMJQ/5Xy
4UEfB8iCeItG7f4019nkhC6HRA1PaLzV5ffuIeHCwWngJ1zPXu0Iski2BCsz+bM1pltiw0trR/Nq
aW05SDBZNzefSwhOFmKf94RTb4lKdFr44JJo4KRkemjnA/unh5fPs5kfKdLp84lNA4wMnGMak1AD
zdndJuZq0Cmvegq4d76p2eJmY3PbFq1RAJ0/AY1Fes0t3hbBMbXDZkelc4v510bG260BKa9eMwHn
ikjOcOdRPadYwSe3c4WTrAzGLPPkcdVPeGf5QP06USTsYZ6GsOM7gPecYslydHjJGSqqcspO69gg
OJimsDlz89iPQEpmETYkCb5DkACY9I580cfZ9PbKP+HsbRiCOSFSM/N3aWFHa8wm7DxtCM3SeUKa
eIUu3QEpkoa88HCJxoTWKIX56fQAMhO3PYKbl/cTGZ4x6sQvTt1dGSbwStCZYmGoM8GBCir9sEvN
W9rxKBFi+h7w5wDH5vk4ymqeBd/1b0XepuSr4BhzoS66F7AyObPzkt/LVvYTQgulGsK28zRhD0KN
DkLtVmS1VXlAG6M58fKBAijDptf4njkO4vaDx7p8+d74+japGuqC+SIV0Pil7hUpsdCENXhDZmI1
TZyhcquzdlfouMc6a/P0FJOx43ZtIZfksqtOeDe/S/6xrDHQxC8K1LkIIVMi+utfZuUFVCn4hdj7
2ijmuifrhysIEcUUgF5+23UG+pGTZ1Jr+zRMVRSrUTidqkKpz2PQDHtOH1S8RPymcBhMZXAD1n6P
MqFy8rnzd0wcjsOc0CIC/FWqnnZ3MYt9JYtOoY2I13JEu5+5FU5nJkxQFzVf1ImG5FuG+w1PVtmX
NcxNyCvYeFnc7nRjVpmgP+xlgbe/676fP5bK9Uag6PZbwYODsq2Gw4si7qK0dRLQeDWlz6wgBQ0K
nhMVuHOA52DF5NrcZGeMF0zrCz7B8hlmPSmuKvQcJNyUOQ+tP5rKYmYhTyqx9dyp5eL4NFu++Ea9
Zyg4abwEubeklqZEvWsX0yOOeyR0UNS4Cwy6FeL6FSrTFkKhvlS2mXfKLYS2kKqb4GDDHuD3m2Pu
ke38moOdTfdahjcWPZgvUBiS/URiVcP54oLEpq5rwUUdES0wAmLv3o9dQG6CzcFeghW7rrYnX35j
FYHdLMYZQanwqD4/7HSIbpeo1Tkm9enSKqUa37CavjGCXaIvmBLyx9d30fS48+spAbH4Q3k/Y6jF
g0v8fohqUSZgbAh9BFvoA9J5edWZQiW51QV4QSb78m36fpa/Kzt/pBqKEeyG7ibbmPuOvbauMfAa
dlsTkr7N2dtYHQh1umF72xx0HQXMNAuvvHHslEk3/bHUZRBrfwG0g7SxFlhwxcJ+s7GoejqUMIhg
MT80Y0BwuQSpKZGKODsqshLJba5IgSNbnJLjMh0pa94N0nnSlpU5Pj+4Jy8wgaFCyrGCTwn/d5Pj
29FJP1v0Y0vCLrnn0hFV8SuwrXA2FPiWL8pvNlEwq6lNFrnVE1CxT5pBdM74xCWONUAa0F3u9EGh
ohbA68eSpHSh44pR+3S+Qm8PU4AsIVkHUd0PK82dZHrg0snnHQkM4T+WtLhl5nyqUtgNW86kUq75
ag90/Hm/E7G+OBueKr4t5d8V8LKV9mc377Q5S0wFnCydryk7rb2Ft9bd67xIwRoeSgBvKbGb6vG7
F2qfuuFZP0AemXh4i0F6KwtEICtCIyEzc/mJGcQwPlDXZfpiQm80lLQ7Rka2KWrgRbD1LYKo47xw
KvA7bcCXZiMju1rnMf/6rMHfkE8zY6bHvOgUXe/zjkA7bCjFRSZI0cwTS2x1lJLBCPR0nPs/ls5E
yl0Qd0RLX8Gs5ucpOT7KEiA0662EG2nrIVJ6RyyHAzXm0F2PwaRQe/342D64U8ps93EVke25rE91
KeWugPJk/vpdp7cs+eYK2QKlJraeLB1IsThyb0puOOssiCfCI9Ge+uo5lgW7VFo5XJpyNOZEMQ/k
RJJw1cdaZBYZ4K0xIOwo9TAhGLGVUB7qK6VDQgotE1ppWtx7DHTUa7bneyF5h1kfA6jOL1T4NYxf
h4+oDeD4b/bjb56q24pk/RQTEvfaUBHPKTBXkm2T9qrzsBswIQag+rjc7TpG+ihqVnIKDyRWBVVo
4URot1ycQQ7S/6lJPUQ6dI34izXSTuamBE8R4t/WRrOBkjkZ0F+2u8K36/P2gwdwYvJF1sHomolP
O9FQa39jgGX1JDtE/+mD/vvYRNdv5bTW5MziHcZhfOEcRMRJS2p0Ttna1+2K1C+c9Gt3ZuWGUiVE
x3hGgY3cTSnhXOU2deoWFJey3PuGXE6E1WdpWTebeG/1xPjX7icdYiESPkGqg0Sdn5YO7b3YW+SH
kzYtp0yNMojIzMCbK3u6ieIapo2VmfMJPzNG4V7fhdMFA7/MCqetORikZr5E1QRGizUQQwdINFkz
9dGZlp4Qz73xbjw+0GJAxgeTmvIylQI/mvMkJJOYySyj0EilHigvhAlg9dnYfeH4kJkvwPgagLTn
wU43DYmcz4Z+hNIlwdJfqT+SnuGJV9cVO7aryb4mZljK0lVffsJKE1Spxc/jRV0zThlh7dOEm4qk
IRwlj628kwn8MsI5va1ARH+Xvkib8SeBapfeq7O0S2ajj69TEXgNd+5QmVkNQBjnN0kBSmIVgWAB
WQLYO325aXh69GQEds28oA+C4f5xtsfVVBXyR+e1vf//NU1RVqgaYQYPuYJhjMhZnqtDR8KGMpq1
q6jsiC5BupDDSRSTqG1xAJ3tmi/0gHBChjXbThMdN2/Erb6cYAhv1kL3YHOLvyAjCr5GGwP6EQ+X
Q4n3JyDlHGie1lJvMDrgEzjtNhFpCXtgA5BhNSc5wTbEWbFg4NJS3e0XxlmKimg5qVHy0si9EzqW
bs37djarU3SCw4D4RpaTv+OMNZWhj6UpQ6TQy9FwScqihKan8Sw2sWGgixUqysgQJmUPccxmx0t7
CKyq1R5A5c7mAofSESJ1rTMYeKwHxXsDd+8YbPWHQrhWsq6pVAAGuZxGR4MDNziyP1Cvxi+RUSlj
I8sTg6tAsK/Lb2yG0bviT+Ut3/BrnREuW7RSQcRoDFsIfCagvo8WPf0sEqAFTEnMCTfGnrQnj3YJ
7Su6AObG6bTCTaDRwL8u/K/p1xbSl9Y05jq1/2m8aTKhN/4UrKkRYjarVAeDtQSVmapb4DHHYvO8
FsiW2Wcp54zfv4zacnQ9KvbIW2PN3Q0WGAAlw0FUOaKHGmIJCj9wSVIWVZ3XhavYGX/SrS5pDleK
sNvTcF3pDs6ZxBZoGEtfiSjM9L9N2+6Hq+z70XQMV4L+3CXWMqfBTmxGHd8JHAjC5S5iRSSEsosE
SDJFBzB2++5ZRGwfCemus9R4Igg0cTlbe/N8DAZASqlnJ+joOJv23izC3L+dGdKRoBFhIo8NUd/0
Eg2A9mrMNFyMXULkAM7+ug4VTSyGRSd+ewoVCuf3FWOi4Q3YntaxAGPP2j0P+LIsW5JOJZoFWgfO
PUlwsDpt3O2O/TWgRgQ0V3ldBVnqvzPQgwcP+r9wntrwgcTthKTKKXB5PwPeI+14vjy2XPq+1pxF
pNHINznYWaCH1git6JPbaLzhQkctAzQqNw9MWZfdCgFBaUM+40r99bVbIEFDaGJjIHfvWQq+Jx0d
jHJfOoKVzoGPxC/QwxjTvI05H5lxwI63diwdJW7DL86w6DJQAXYtyf/ObDBAPx+0LE8NL+Q/8tix
hmYp+qlt0+kgVWQ6bTaoS87P71FYORcIqYNhSvoTkv2CCkapqxfwLoZNYcO2qgnD8/rKvNELb8mx
1dqLJnUzfWIvcqKGrcoakua4P4NFzxA4j4+weoVJ7DPiDwDiIgdP5iokaUPSOCFSyJokO0NH+DYQ
CwU7t4JSTmF21MtwoPb/cIKSyFMJQDpzznX9Y9Et9oXBgosigQtLLc8Rc1OwzfDSEqjwCYBJglp2
hgsSTReswy8exuCSwL6Y5d9mLYc+M1fBy0SbqvGmrr/b/RcU2fdJSB6ifF2rnQ1ywdTnnN37MhAp
IRX1NL80k7Ij+5BYv1P3hiFikmh4Ufm/2ooJYf2dqVT7EMuZQMxGtN0Sp6LSTQtLOLHvJyTuiY5Z
Lj8v9/lJxDSLVDvcfQYK/PXMVA96/EwTtQEX6HTmeACQuiLi6uOBAk0FdqRoFBmott9rFz72J6SK
JSH2VYS9VPcwlIoFIMJN9puYJ7RrQbN5URMXzGta4ZIwbxb8hXN4S1kWYuSY3ZYeFz753efmrSbv
G09YLupKElmbr8fgDGSVnhDCWfaqIz1te+EOmq3GEWasZGBAHfZZ9oEFVGovBVi8Jf0vMQV17TTV
/T4ropaTSvYtcGpjtZZ+T/md4YT+WuU/EQj2KNxJtzPURYMVKGcSHt5VHKx6UNSREBD/PpwasAW/
IaXVLeEM15kwgbXyAp7fjpk7HMYpUjqyeA4mT+8RmbyXw5RyhbJRoBwQxeVUNDyCKMIoCAMqH1se
KH3Gkc5NhA3iFZ+FeDXkaSLfJlHsmMDSXRorcZQtqUlHGyyLID20jHgaNkbJZ+VA5FbTD8x47EyZ
pi1T5mE+Z5QYYlfYPusIwumSwtg6C77B2ebdGpZ1ho/+OIOQxsSOtnCIWwHgImqZpGbFUbaYI0W4
WpSL4BVCjGUc4wIXQqoKmw9CUqbNp6VLR8amBLQsE9Yk4+IfMsK3uGvF3PMwYrIlYxRs/WkB5nCj
nv8fpmntTLLXsyA9JPv9K+aQu4doIzGsOhtt0BpPJsbxt6F6fZkLyYv6pQS4BXzkfz9v9rART75Z
Q81txCCwRR+QFmXx1E1RElqvmJPF1heFxQIcEzqw56m4PW9I/hq00Fw9wUaaFblAgxFdS4eqVC3n
bTXGnmeFrC63vj/U/h1dBvs8H0k4CqY4xmfeLHYYByrDfOcc9HQSFggi8cucy50hS7J/a36Y7xIP
SvMpqFlPh/Qw9CzBkp/7XMar409BN/37zEi3rk5pPn+J041mgiBuautXRGjB2Lky2G55mHAXd+ch
7Pb8wFHoJsNskGqGuJUvYZksR/3y/Ddf54+hh3pDw0MZ07aSaW2sUjHvxt6WuzFl90YS2lhyOYTQ
xpzPb/Obw20NTYhhrM01Zpo2qbwDQ9Mfv8t+jpm8ubRdZbVGJiIZ9BGLvmU/ys1dxetYbVIY5r8R
AM75f8EwyenFvMvt6u+1lWSwl3a4Y1sDkK+/jnm0sbjZoyoYnFNaVi7W09ESeum8BFW4afheWkI5
7yeV5EiD9knAiNZ04KOxniS0318kQwZ7Ojh6pq8Ecw2NLIypW+R4oMOTkI6LRFht61pKZHlrGomq
i84IO9Hjc4M5sB/Qfse8GRYrW6/099RHJOyY0xHTV1S0c5i2On4hHqvoHWYzJpCBZzebjHvFOm8N
oIIAkleCiLfGdKuSEnMkfB5j9j9UwKbohs+66beU7z8BY8ZwO42cEdkszgi/6k3E40UtSiMkrJ+G
Ui/E5B8+an0ck3C/ipbMuNcU/mjBcFzbg6BVoI5Pt/nPFUVDbBBT06ho6EUkjSCEABjXDagB9sdb
Ku33qAztvLfVDXQaU1Yk26mdA8tz7T3iF0rPFttZ7Hn4uqJNfe6AAMW6w+sn7JY3Wv0EA1qqvedO
HI3Owru0YiCDEdb0HYCFVzSUOXKR3Zy9XiEBsQbgBPM4CioEzGqSxj0mb4YoqM8zT5RRuTBBZnr2
4oMfTOa7GGAycQ/oUJDsQZaVH3G6qQ1n5jL5JrP9/8Yz+gCIUSYn1P0omJCd8V4NtfihhBZigRX8
35x1ljVzpX2PT+35UPHvuWQKDC0IOF470AiYHHcT/VmTOv2/wN9eIK12fbq86enDqSesKkj+9qcO
Ue+yMvL8IPMATi7Cby0qd6ijUALjyfZwhvHZxNKLQJrglRiFgdoOVRjXQ4vcdq66x0F3M2eqERt+
pCfOalHsCLGy9zn3G0h9iWb8rZ/P+L5DiT2UtNxBdX3qZMFnXEbSG73POZeWuSMctxUDd7NvxpnW
Kg5nLDGT+h6EkFwdwl8pj1LSNaZxWNql7K7aTOJqXpULxd99r1rVJxbcyz/fBANaQwPzsRFUNpug
xMpZGjNjcuRYsMIpfxrb/3LmLUo8VkJo1x9Jz6wX8sFfAUqdaLwtCxMzvju0RngZOSoHIznGp5Dm
SQ6htRCkCrAs0iU1MsE+Q11o/YkAUQhhSPRzmdIAoiySm4JjajHaSGXeMSihbPg+KiGC3lNhGEod
nTQcJIIjUDJAF1dUCpilp1HGvBx6EATtfMRHYMdxdBaN98MEdZvreyBIZf63oXfm5kCYB0ALMfZe
mMjRBNNxWbAipmmnnoj9hSwh50M1EwptLVE6zDwnAw5ooLnbp5vk5AdJgAZbXRzkx2eBOZ0A1GKO
OsrjrmaLRLXzNbYjx3RaHIZMNJROV3mJxGbaEd8HcdsTzyT0hW1dtvXTu3nm9gmLz2vavj7B6tmz
pMTM/MUIx+cd42mHBgs+JShPzc4o87luFUn5QZsI8ajsRuHIphAMQdnXZOYGai+7ZazTs7/S+1J7
wXwoze5E2xAOUZbYpvGagxSxmTQbwNP+1wu63DNBhUT/luENQTTxubtFduDuuMLEnkAsHVy6tKJy
LBCoMhDiQELJ8I2vE3jksVc+rApuAEWWEAz4l0gzrMYadsTCLowgQ5N775eu5F5OWBl/yoNbA3Jg
t6aKhXdxhrZ006sgHt9M+1+PlyRPb2utdp1+SDIVpXF1nMLk/ZhQ9Qh60XMvEj8Fu2NPhlLmL09b
EEhS+n2B2EX4JwPvBW6Mlao4kwNlAKTM2AE70qadBlwY/NFrBL3UDGQTqdvuWtarNJZ6CW5IZt2A
0MUD0cgWUEqwdbXdszO6km3F0T5HrbwEYboEM4F1d5zFf4qt0blYqaC8pxo6lUj6JkwbOCiq8US0
b8VTq4J1G16cec/JGuGtNcn5MHN6ShYKPiW3/OiWQavG9viJU8HxUiJWtXAbM9xpXmg1KDJfttBz
L2uNMvM9LJYuTsVo/oozRkAmR7gbIObTWZd4NYOp34NGmp9uTSGZl+qKi3GGjHELa2OLRNj5nCte
7i2wCOjpAD21UvETzbaTpCpEVEUIBxC7REUPlIbFeG69soGk0aIKIZ8hcJIINOXCkK0hAB7zAGQk
kZzt/Db84n1h2tYOX6ahPElE65KNM7Q53RC/N1OGk2nCaDRNMJDOwqsauG6oPNEjj0WpKosWozSh
vF7Ehz1K/xkDdmk3i+MZ0QeaiT3lUBocPoYlmhk1+TwV+4BfCwbroz4HK8NCTsle3JSScyEL/2PK
PiMcUBnFAdGq650iMljcFqBFaog0uaOp3P4j1BYvW4dHlKsOt+sM7CQP32sq6CWKN5nVYLwBASSJ
Wli6FrY5wgpqFrxDlWpaWFHW7Dk6kOUKr47rRUNUWVup2J6dTOWDoHRLy1tAZXAD0me4n33gRqy0
Z5qi6tccmE+Q7thpCmQAkuiRpAHsTIromnKBp/MUx1I9bO31MX3ogO/gKGVehym6+nmovRcQRheO
+cJ2Ew4vXJFjl2r/FZM5ZCddGOGQHTmQ21RHql6RRH2XB0/kjJuav9WrbVn5ZXiJOblYooD+EYww
4IPYx8DvCRh/JkPlnKbP/9CF3OCiCmSx9IeGdsgpXdCZjsyMnrkSwu5kjTS9jsZAFZu3HlJKF1dr
lBhpuLs92jBFGtH+7iSl18+reJGg8RQbbVYU3/nqEFrk4Iq7v9aA70nv4CFrcg4R85cFvqyzcBeD
/lT4KW/ndFWr0t8DDmKcWYTcvA07K5K50e/MLvvQ8duNYCAd0zQiPK3hMYL1w9vLgFf28orHPWif
qDfkeZQVlUL6LzuZgM2iM063xSBnC0+CTuKtHo/d0x5d+G571nur+vR4Wk4iVWNf5c96cLBGNYqh
g7CGMwm+8h1Ad0ZuLg2shnNTG6962lOYZfblkA8GnC4hkw4tm6iFKB6IWxrddnrB5ukEFVU5BemX
j8bM/FTZRxxBWxOTG1QI7T1fZH2YZyntFLSCwV95hEW0nCVm46R1b9G50teLiOoLvUugix2yoniu
T0y0eefz9nQQQXIS7idA1Id5OtXmBv1OjMcjpVc3q1ySgI8iQVzdaKstc3UN4VoXYWeEQOhKvQGv
uue0cWzAVv43vNSHMG2vhrxHHOPgWADs1tWyJXNTHPe6EGfvj9xMybHxwpO1yMaQs0a93nXXZ8LW
r/MsDti3M+3vR508enLZ76oM9Z2pbO4s6XeH4ca6yHMVOaOdzyKhZf/6FF8i2tCzxtwasI4UmBAd
RraFoFS6EPFL9i4CLEtCv/tuXTi3nVTw2BYB8botVGCHUG/v8vRPNy5TDouJmVyJDRFjn2DIrbZt
dXxb6urlk/iwhX0qhHO1gaBMTDM/jp87uIWHcWncKqZDKdxMOps5bLKeLg/hvD1wUvb6f2Gkr/EH
Ea7XPfloLcLDMZRMKpb4lSp2sjY8HIQ4xCDr+v9dXlI4a97EbnXlyjCKTmbKHKw8tmIUxQlRBvSO
DxCPGiiIB9S/8PpPTpiAzE/rUshNG7rmBiAFdlH5I/vMNoXIkmC2qPHTuY8n2THmULyv3vlJHj7R
UrrEJHwjqruLB30WpQ3/CGjXmeyS2GyBsdmQJT1TD2Qz+ZM/5MFhOA1FM7DCCdN8GnhaRV25ic4x
EBl0/ISK/8inPp8cwIw8yAgSR7HPcgISXK5DbfXbk0Uyblpx0qV81Ybo07stFLN1Am/4KmDkhxDa
RFoEyEEbWz6zUBu1991lOrwx8E7P98sKCoatGkXfIllB9soa55QOlN459403tLW8/XgJ3ErPu86/
Z58JrPMwaFVYiOq/qeS+V0Fp+yLWX4MRocn9hsNg9fFAM8tL85svbfkviSshsSYuwqk1VGbFouBN
rpXKj9jlLZnE/A2x6zN68Ux/Hrb0/07bURUGY6TD+Db1cVHkXJPEinuV20qB50QpXc8oQzMRDexZ
rfshfbkMoRlto0kYpb/vrf4Ql07Mu5tK3TZYialx1jfbH0PijKueQHHQh1eV1/kROPVRYv0WU9/m
lmY80WixDGwI7nOz4iSVQtMHyj18q9/q32fnUv5Gk+aZk1fOWivi3Ed2DomMuUGGzJhY7LjCzHip
0VOYDiJKMxe1TNnKWcXR6tJt7yiiXZMOqjki6oUS3KB1zMDLBMqFsc+OIxKW63+0BwBtvSNqVwJF
/zAdkGmjJbjRPnZpy4AUqYQBsgjJNowmYTho6oIJ3hZHJxmxxF89NWotr+qp/KM4CdX/PpwGUhCu
zvJnZK/IrHjzDEwwV1vA9uGp9NycIrbU1Va/XEbELWG98lgcXTFt7UgnrTi9LkTNoNPkyIt4s6Sz
QC2T8ckQ8DX11aZtgi67Oe/BeGWmG4lRv9n8VGgbnO71gPo9YF/V0dwxd0hAxt36ghPaDahiIJ4p
ymgN0y/bXcoR5wim1sfSbdlgXA8F8Vr74iuVFu60f/UKChu7p3i0IO0Kbx3DRSgTCNsTG9qw9y56
dHX2IPw1+tsbE7dzKRmfmQkXfNXfNVwe9tbCn27hGcis95rZj3FU9slXoOUNsJ1gPyPLLzIwHJOz
6CWHlvp7sy5Vvk99a3KEC5gCrGRis3BVvedFfPP5ZEiH/d/kuhc0JMaHpVBWxtI2zO14KhLc3mgd
u0QFOZ+zPgD6ng0udZyTHWDZpGOVPwleb5sbDTqtJMGeIqV+EjaQMJD4+K+/YnFTMB3tgfg9sf7+
COFexcun5BTJsPhx4Pq9EKiwLGi5OYQqjmP8motUSeZOo0DKWsgZxre135wyqOOASRTcX5GFD+UO
1yVCQ/UPjsLvpZAKyvkdwgKwVvd1NzNx8UuIO/JbZHugbYskivdAPKSjWZ/XO6Qu85/wdwI3bTDV
FTutV/+w1pfWbbjvcarCEq/x15dtP6xaaOiLPY4gSEts4bs7omQ/mIpg4/n8JaK5mDmTQ3CDP6/J
0yyXiA2swz2ms3E3Z3++i7BIBVHgKx22s8kFRlVXytvQrJYoDg1w4j0mbIoySXHh2gMsPPXmUV+i
eP+jtufHOd1+MVDg5MZt5dP32fb3dLHBo8yI9q3aqm5JMaR48OI8E5H9Y9sOclj376Na2vkLtqVh
bnwu8qljaxOtnVGlvJQCuarVeqJY6+N5zg93NFfFu6mFXt12nspF0l+pjhLP2hs69VhRkilBo9Iv
sIzNgW+2HMsGEpjdXJUr2o86GFv7WzquiqEqvJvOntM7GGeZ0TO7W4SyWig4FVPZvbo6cd89UrLZ
HFCQNcFOxlPXFBCHC7w/TjpwEhnSBRliYw7ERBJMK587/VfleaCklS+k7cIsg5hhc25UevtjprGu
HDZ2TST4W7yR57Lsrl41PjgbD6+fMbqWNK9AiU4zmual3OqML3SCiS9/J7smeOSfCZLSnUacm/p0
lCwfTTrf6AsJjsnfX4yr3yKSp9pxMfnwfc1RwBDD406u8g19dshwdyjtrJ0OkRyPa9ZXO8CVKxSS
YhL4aBhao4rjx+522cpsjUO4CagGwUYJv5Bk+4+9l1TN8ek+WhU54WpD0PLjUpBEzvp/a2GvmgMC
MXgeFjIe32s3Z1Sf/6jfxgvtKgFrBdUMrKLmo1xXpHNspkfKWlsAGRlR3dva4VVdrmYETYneNzCf
MD9CtuLOIpY0AZo9Kj1qOU0o16lMrPbNPg9OA0VN/GvOD2633pAM+e8/EGu3Y2Y3ApANbPbnfRRr
5U2PSSVX/h0EAGFzmvo4oYPOILZ9jln37ziwoY+oELeGUEpB3OL1Pg0hwJP4BR1diZbtK8YsRtOF
vNPrrB6Oj8vu9rHg4yrOaz+eUDtbX3NpfX+KGriRgCq4AqcOG1Li6ll0V5VocyaCW4P3Bp3lvtPF
lZJWbpyH3qyuVjx+IXXkM0lhPMt4rwPeK9GTMMGND66jSNVtesVIBBmUPBj1QS+SRUnLksvPBze/
QLBvCZ2klYyEHFGuUZk+nSou7mOdgsBE7VXn+pp21I95Kyu+ZAeBg9lqKhl00QEBni1wHjsSX2Vs
AlwQNR+Tjq8DARqq+ATuVGulpdvaQA4TneoKRpd1XzXzfgAz75Q1odFbUGXEHpQQJj6num+V+7Ke
0/nq4jW56qJ3+lBF+ffXTT4/04pkoUd1043JJaIwXI3xQm97xwKpQ7MjlrWimsUPOPyHfGb9k7XB
vuxxwJNCSCPo1gBviLGSE3qCjO1w2XFaqSIWlOeMVCrwFyXkB9cLOtP28cTF14fwOeb5MmkecFC5
UrdiP32HBbO9Xgs2e1eGDb7rhazZmbfDUGE02Xy/VIYnBuG/B5F6xV8h4UW2rPP2EHzCXHpoYuEm
8I5CcXy1Y5/EBHUkcXGc3GWtPa97jutqSIk9TEWSYY5Qr/Hewr74giilYTt0ol8bLo7uMy8KTTOz
p7pheWUsNl4cHD3YGHk463K/A1g4EHAJQySO+VcTbqiHO248NdIUfQ5dxFzZLLm3k22JSdTSd13S
yqrLZrV16Vpv2e8yCD6u08ELiaT31zhLZ6l36zxx3vapCoahzaosDIpabr+ZUn6wL2qf0TRzwipO
3l8zSs6zWY7s/lphenZy1sM8sGToGoSI8pOnf0VjO2eHNR1yzjtj94Zs0ZbO2vrHiVBzNRr29sbE
LQIDXYobbxVQT+NsaM3HiwkW1VLh8USVcSkSoK+meA9qVbnUOU1QF2KwrLPcSecix7FRf7OPITLl
/6oRftZn8ZXY68DI4WaxMgiM/rXIAgpW2q1jKTY95Cwb++nCOYXophiA/85StlPkCU66twDvcZNY
D9Qj7lSHoYa4bdmQ8CQZMz3ZjhLJ45sSeEIV0mfS4k+U/11xN0kNCCHBsAnCF51FJjAXDrUmNGK3
XsFSQGeCCnuzyIpAM0gaJ/ggCpg45emk8PwQFRMGjUC9oUNL1c4xAnPmxpdmX0aEWF3SstOezvY7
LUS6GPkhab9BQe3m91cYCMggbnjIn9CZ6SAD1mk0D3PlU8BVAu3hOk3BXN6HtJlRd1+52A0uqjLk
JhWyf32C+JkLDf9oXp7iTvRWMsV213oIdLJXG571Vhbc3k5TFkDJIqp5CZFHAvKkL+1p6rhlW5nS
fBKbZ49gSgr9dXbxQkuwaa+lJcrBo28jNjOEcBUKIQlGxXUzd8WeO1J8GRTYDSswFooIxla1/3m/
QB541GVOHSMy6phxyumA834DpvlLm8rLnnd4vt1PZ3ijoqdwtddoiUw6zBAdS7sPLG4Su/w11rIS
XGZoiH12bRrpb9Lq0aDDxyedukZx5dPHf1i0a7UTDm77kXRzYL9XLv7/JWgN7Ogp26Dc6upr0a5E
QVUow4xtnnAOnoxrRTzpX+KmYrI5rvfEAf+ir7iOUul0iwCJOSB6hqhYpQ+UHlCeBZ1gEWZk+Ocw
L0zrIHbiZLgaYiz6shsGvih6g9jXIe4qEaATeyPhgnd1kc/ktC13fd+JV9NsLuW9wPmM7aZXvAZ9
BARIX2YO1yuQSmi7j7SB2yKzP/xflRQSc2E9M5cTSIiSOpYypgzcBFcl9iHpF/FaJ6YuRTSNPo8w
9UxWdHY/EqQY+9IHFb0V87Yu84CdCepOFImClv02i/VFG09xMphXpeEwq7LxkiwVsNH4F7fOAF65
RaFltcYToiznSoU6R6H1otdYK8s6v01hgFOilzJ54Nw4UoOhAVPCkoGG2/+sgFE5lInA37k6QIL3
OBjjypYd+ETDI3uJcRNPiT1M9NQ/R4kiqe22YnkCJ2y6yhu/H+J1zENpZdmDgcJhATnPoc9L8Pey
RaYeV5Dpj+snZTly72jpsQ4/Dg6jAz4KOHPUnRo140mA99At4JIIKn1Mo889M5EKw2HI4chy94F8
tDn0YqdnJ1v1ctsJwCgpT9rBfqQ6AVqbkUaqQx7JysH2ZLxcUIRq33AiJIKKy/z+9gWLE4ITv+nN
HzdflweOdvGiwMgKZbh2NT9+wQU+Lfi4YRPgvp6sDnyHtct277K0AQwETejJv0FFbM4OAbCVLcx5
Y5pVFsuTEIWbNnti2sZLov47T1g5DwLZ7bTzNXZo4dWJ6G8QHONsDkOxt/sC4IevDZcOfuDSBys6
HDgiESlDXAenLqFzotA8GkUMcb7Gz5nFEEho/bjRO55rKyYJ/UWF59gD5/JrJzqsgePXi/NwwpXr
eMNiUISJ7ff/jScDMtA6/cgCVQ+ju58rEyPmm5wUyn0q59aktJaUO6stPICGb40dD7LB6QPbh5sf
9YI3BOmnCtKm6Co5DTu+aCdkPifnO4L6rYmrdhowNAUyQXanbUcetT4tWYA4n6gikeWOHsYLFyPs
X/kew62ASHKolcpjzPXSMvneHQg10kS357sDReSV8jAIMnHFW7g6/ITZIFfkCdn1TZLqQ9uiMJR/
CxTajHWR5B2jEYoKFTwu/InFvTZSUUUFxBHPW7O345yfCeHiGi6nVyZ2mmMnZSWwHTVGL1ALf3H1
rna8dkF728ZytDaCJ+yl8t11NAuWuZQiYqhHiYsKGk3xaErMlPDOIqyyWMqeQeA+klW8c6wH4gCH
i/dUrnzATABxzzcs80pG+s/9OIn9LltrdkoqqI4MRGJz/rntWbJQwb6/gNtmPLHljchDd6T+f2J+
KHJ/URyLEQdflOp5IPhH8TVH5lsjgQEEWm8Em4quMjPbwTyeZ6hh5EP7kSKyhtmCkTrrhnkqwkmR
13j2b9syxJa7L13XUq78jnuPAU13CBznulWmo7JMRQSTgbb1QfRiY0iuEvSQqBgyAnuMXIGJ0hlD
QGACBa6gwSNVOaVzef7MqNkeWfs4JfbJgfEFhGVzejvkNpK1YMmtNnYhxVJD9hJGoaAB45Jvuz83
y5ys+RZkVLPjNAtd8abqRlS5qZIot0375GV5NN9qCllbBj8WXBFxKyvEXQIiJpGUFJ3Ti7xtnpyB
M/cng5TVmlro1+Yc/y0DyqYchungbnuI11JFjkkHZACaGcoceABpbYxxnS2mXGfA6v0aG5qgix9q
mJV7TPfARqtXdnsT/RdgfinPj14YnOSuWmFDGU6jjCjyklaZmlXJoxJJP5t/A1tFENvXCGjkr1Z6
H0jh74fbF5CumbHf0tdFpDPKCfd1ZKIZDgJA9SXXPmRgQaG0u9fXcNAfPkMbkUCvLkMP/5l+lSSz
iorE6alvz9uvv6XvkywQGzS326zbmYclL9XHuh47TeQssDWzcZElnKWDUy9dAbvwPy2NEKU5H6v/
lIC4LPW58A4nvVX2AiM5HDgCb/EQl3dvoE1NV74ghPTIluGN/dOVGNQ+JfafdmZoctyRWtmN1gY7
xvkiLiEq6uoJJy/RpK8o0kDkLkedsB7nOylbmxRqTHcmeydA7YMsBYntKtfFynJZKaLkOzt/sEiG
+5XGyMFcbIm1TAi3150rUvSqDXRRTv0HWrF8E2b4/GU/zfULo/Jx5NE70A1W/0GZ4INWWeTyfUM1
B5NxCk9JxzWNsUvHyyhHkUT7Fe8EZeR2+jVTiQ8sjSRoNL2qnIOYJlebAlWn9OwXFJgwLKcnegV8
YzAS+PaGJ/xeIQ68f3t8P3wiFkqHwRlAa+eTMFIqb90NPIxjUWoaPSjPx0OAtuW1IxyeI6ZitzgG
rStzSU+gXFdAWbgC2JnoqnEXqog93ASzCR53lEI90/T46NlyQIFv80IBwh+wy2Aoqky+HeCwIZWC
evGIXhtfSj42pMHsJ7EeCP0bCsqnLz1vEMwyfZ7xRcHP/gJyOc7PDBNihp9x0p0KgHnhsDJxm/bC
Td49/zSu6KGGZbABTnHuMTSvGR+Sln2/8/ZaQ2D3LBVWCZdnWZqj2TrMzh6NJg/j3uY7gvqVhR4U
Ax16UUXQ36qj8vd9d4XTizCLyS+B0NU4XX0nFpoWDwcIQGAJWLs4GRev4Dgj2HnrdIUA8pB2ZGSq
6PSh5LJzfLI/++evjZQbpYgS5DpjjE0fiCS93UmfOSckkWNy2RDqPLMH8sVsQMRGrjr5Lr3tStBk
pZxXzWA925cc9JAWp+fshbJeT4WN41ppUQmr5JJS4lorMch7lLu4cFR7Sqo4BMIOSQSBtizVZvji
GeWaCEiefPsImUHmcL3QrkmztZwbDqaXxN+HV+ZGZwNjqn3MYe3Nl7/uGlza922XmSUEw5p54+ZI
pv6mqx1GNlNeinbv7AqbEcUbw+BKkTZfiKq9h/4I0ZBHb6fRDMk4RRfFB+mF1+6IK2+qUWxMvZcu
/RFMfLgOw6P4uvmhUkDk+cC37y7ZxQuTCCdWBnHtkct/kP6WxTy3/IdkL6C9aI6mSNpmh/QX8rIS
5Ie+xr9hhlcc67EwuVNQ/AhjL9whOo9LXnizDAm+3bSz1/SIWnOjGl8ilpwqXgHVKP0kekqRWdBY
lQBmXO49/bV/A5SwNZ/6PMTlml7DGggwPx9qY7zqqlUmOfKtX19m71TsjrNG2lCejkS2Woh0Mijq
0ixwwR6zJzQ13SF9/+++4dPU31xdCHTx5SC495//SDqLzaRvdN6qfZwj837GLfAGciUsdW0fbIAn
vlyKHrYLZvGp5W30g+3VKgAUq/4OrCHuiNOdCUUdAPm4k93GnZhJ5I9+zYRmjy3i4Wz565WJVYdK
jY6SNx3NOf6pEIGezOOtGHzHVdUL8gpP7TexyVsjIhoHAkSnmXlmvEtxcgkXJ67/dcfTaFZ8zslr
F4oRaPrr1R0pE60osNF8Ty7YQxruh8lytHGxOiyfarp+8vhhMyzFn6BsRuWvajaKEv3eKTbuIOOB
d8PRx6juJhFkY4wIJl87pwzOPJBEQyjPj8Gy2srgkk78obFjASWfkUp+v6rn/9ia4cds3EmlDuNM
B/X/f6nfkCfebdEiTJfv80GHK8J3T2G4nQ4nNpQ/8yCgrU0nQog8OOiimPg14QRQW/nwFe1I8r5v
9Yv88DJcsl7zieARMButpvJlY5U2wPqoowZ6RJ1nBxAEfjj+FBF1QZ6t9jlyNOn8kz/ezMu4YbHo
CRVAH+rKsmLn/AZCn/6Fyyru52H0DuMPqk/qN1YGvH/yDziD+KRmUDM1mLjp2sCOCNXofmW6VZgV
cUio7tsJo0BPw8mqc4xKcufl+rzEzbnpDDRupplOn1oX138QFzjsU2hkCq7YHZm5B8vMTGn2Echw
KwGVR+Wpd09x+SBjsHMNEtH9BECDvh6x4aGwp9bdrcFN4rWO7NX6zIHFjWIIJMfi9CSIiJzi5QI6
87qohfFYf39CydkVrpvj/9tpbkhPiIgw5Pb5UjEftQeYxngsvmdHlgE+Wu6Ib4w1IIegnw8PX1Bd
ix1lzoupMHDgh0SplqcQEDj0fVhQDSZ7fhEeWrsfhhjAyOtwG5hkLmthUVmeC14K3vhqVvhSraMS
hwMuH2ZWb2SZDYIbXloZjL7nr8IdWgtkfFB+WyDjRlLzGLPlpyQBNMREhpjut1REpGCN9Fgr0oFu
l1Xvk2cdckTrjkA48KFCJe5tq9NIhYIO4X6BaVcCjdnJhgq1ExQSEFgUH5i5l7HU15UJEIaLsgdn
2WK8/2WVdxYkzJ4ezFZoolEMWVpE1ZCCbUXhuc3GSIijrOPE1DLgLYy2zKSSijuOD5+DYc5NJKB6
46z70HKykSOyuFwcvF/RDVHhVxCefTCeBKFD9EAr6iQ2Ky8Iqnd0s+BU4EgLZYiUt03w9vKodbwS
0DQltDQpGeYn3JuDaqQWmNZhyOFgA2mgGrZBMYFBnqPhoMmqKFKwwS4mCIhqufuQcATt3EWdY1bh
CZs6gRCXzrbwpOofGpz6KCxM1REQqtYpQQa7uV9g2rae3pK5q1Rk9N1LkEy2fD938355qQamxjjV
NZJMqXNdoFcW2L5/it3Lno7k8wpACF7hhlNJl1n0ae00McWjlAnGU8QqXjp+6fzbwwycpb979Yi4
EhP9GKRbnGdAJ+pbw0RCOzXmf/+tffXPH3ZBPJxXBEwRGQjLU/gDRvMn9ShwWvlgWf43GxBCLAeP
21ouU4b/ZFhkZQKabz4AkmcrlmJ3SjJMso+DV1KPQcXAFbQkEs8fSrXsU1oe1uu5sIRATf/zOnKF
AJlvVH9O4RFx6rU4/fujzGokb3nOLfQk1AR42IZMnpcgbmwHk/+OcHPYptejnwWnTqNATdBjAZn6
zxzVCT9SucmEC1QFjEPDxIZXjqJpErIbz9dqSIelABZaaAy0XKemEyUCc+iBdrNdCu3v755gxdRw
8ta3iIHyOQ2Po5fA0TLQn1yGF0YsqdSUuXJdPEw+LlXYcIYEzsJ0OdT7Ov5eLsXUQF7pTn7+MEdJ
7soAdbyVP+Zkg7q0Ue6TuFfhHwjKlbf0lo8/lyD39A4oY7EAkOll2DIWkf5ix4Y8EKhev7mJXqi+
AwRqCvaO+hgnj2JixoxKBQFdWuANFi+HF+2INwo6xh528WcedOc69p0CM4uChLnhIY644cCNBiVc
D8I/cgNrkr8GRQ5tPKGwducCaniOA65Czb5r/J9Dm9N8VvGk9SCopeYlShcPE9i/80gGFIDUI28v
DVSBlBvR5txpvDlolW8ykFCGq9SytwQb+jdWy8xgOlpmwbIkIve2FLsJOSLWOq3k3ozzan6jfSMU
33ZuWOoHIFA3a18Nl1XJ5IRGFppp+dmtOgmAa6AlXdU+ljV4fUG65glk8qQIKi2UR8xGLcN/tawO
VRKpchxdRZ0DE9MKGiY2iPGc63IPsK/fK7n0KazWf1h+MInp1Irt9k8g2VLv0hZPsvbq9wZtbmjz
F2g0zzqkIhx4rQfKVIyzgardUAjAT3tp5ew/FbFTIaRbVXaBD5AxZhwEFsFg3lt7eCk6U6fJRbLB
Zzn7izwB46JBJlnWrIHACdEwSG1sFb4My7bVv3XUv7h+XLVTsAt7ABbuxGQD+AWLdb4+QYs6bl2z
t56MivwgNyi9VzWvRCl/jTyLPmckiyWFLHKoU0Zb1RVsSpj01kZHItBOTEpIi87923fiCrKfWShO
EC2ROzL/bMLkrIPiakZa68E1RRm4FGX/gREIKu/6rtvKKLlHikl7KY/o/SuL5q/pMUwdxfvkQmZ9
oClyCKlkAh1JVZUwgrWSlgFpac5lsaiDQ3QqMAmwLnAVPuOYbkWYmUwECO/C7W4qcxrWnqBQzPVM
Wv0ua4WN3+DMx6vyDEsmy3WPWBUzZK4h8V/bP0iI1YDDMdJ0Z0X/uISRoC56akMOQKeNicykIphE
8Vheg8bH4y7oJbaSMdTbV7asAdIYWitpO35o3aEuDIEq9BHb3PnAfM4pK5p3VHq/7foeruYTl2N7
6QMUCgo9VDwoIlFDTtsI6K3ASRTt+VqXJWuaF8Cf9uuMBgnTcRzpyfBU5zigim3/XDK1pJ37PGZn
sHPlOtcpE8GcXMqqLd1q70N9uSO1Kch214/Jm5tV5AjdgdIM3/DZuvbkEiNSX/vVVvHKiPT8RrTQ
4t82WpQZm+vC42FfFG0omsNy83mUbNmGp4euPdQFtt61qr5AvbzwRtrCLNyXvdLvfbYrjMAGKqpX
5jwAxQSwmEeCgzA87PDxXNBJbiD/kwUTV16qEsAR1q1VqRlPQ0dTA7JNAZK11ATLnJzBjwhytD26
VEU0VpaCFMtBua3KSLYrTbbKE3BwLDPak8/CsGuPMn/DzVfRjLo3NKi+sKhAkr22oO8BXICo8MRe
28NWFtqupHaF2AT1hb4M1tS/6k9AgYcV/3OoDJNWkDn2hUbCcDxGh30WiChwUeFWBzCg8k2v1sjX
eBUdeUNYl2sEuZAn/98FtH7sqGAsfTesZcFla+nTiOAhRnlqfSR25328SkHITCSMyIOCOOyny25y
L6ISLobe4/JEI8Jient/CwSd1IkiLrNkhLQ1LIXbEdOIZCc+Cdk/j7R+D6rPSHlG6tMMbSBM+v/J
CMEwoDVAuNUFTsobxXp6BGke51guHuIE0lS4hXujQSSYPN0zeGeCw5l0unJezd3QzYXvHzu7Hv2n
1MmYw7QucKSEOvaxjE1f+g8A0Ly/q1Pwh/N+PhANARBqk8fumdXPXrrERxp9sPpLoHjy/6PwXADT
j8IhqC8XdAa7/Ox5EKeyLlu0fd6nc5ZuLucHkFfeJX9o6ibCVLCJoIzB6gMetDGEO30hcj5mzzLT
HdNP+AcPWRUKj1MzRsyHdeC/YFlqph9ay17NYAH8+YGfiWlMG3wi9Q7Ar/yuuI8wNvYqQ12ldz7Z
fJxUkehKAiVX0pKFUMmSoRvR4t9BNtyFX6hgX7SWsQ/AnGYl8o9P1r1LaA3A7aXRvrbr+I49y8S0
JJCZgbFeGbux3eUjL0wCMTxvW5E79OvPHjpE2wr2RtDf/eKtdHKop+EPfm99cA5HRn77+BxHSo1t
coykejLqJ3lDQDnbTezQaYnMAIm6zw5RsVFde0atHRZ8mn/olpC2dQQcKIDRQchUfnTjKeVbbw/3
JXtG6YIx2mPz7VnOxyPc0jIGtGKLE20H+B5VBwdZYaS68ydJt4SqFBXROYlvq0maxCdx32zGGKne
+d7YDNPrFkEH36AukZ8foL4fd/Kb63dXgJQTaFZBsIs8MzcfYBGrmSoPHa0AUck8vX7Uodj7Jk5H
EDv+VVYSfmIRnXr6vAhHPKznuC+bQjrawjH2Aq9sGdrwqaTxD5p0IBKPsJKbn+Gbfyryy2rzJpG8
SS/7x8f/PinvU6tQIfoECWsUGKs8v2mAV5i2g38+ThG59YvTN+ofsOrIjPMKF3P1WwMHWR7EFTWp
GYHQ6/0E+ObAO+0nMvx5NUJCYfemy+W7tKo3FAkgwqCzvsGQPGcaAwvSbgkdMyoGVgonFmm2k1nB
+j1RYasPE6k/aF8OZ/XpBj4qa2hV3onUYxDUgb1WSQDdU8mNifKcwPov9fFmb5hpB+X7xPgU6jDA
D90XuB+L0qaq8vCLiwvhnNVoupvmWPxAbS7s2lQ8ZaT0d3wWZRTKx0IcEH0TGXtdZvSQppu1yZC5
62f8u468x8/NVcsE2R/rABB5uALBlF/B0pu+CKA02zyaNL94nOrFEVP34mqJEbxB+ZcnX7EM5waI
oFTQwagBUhIXneAhY4Da70NmY2ij13pEf0xBbVXXL16IVG6uj172W88O83VhY5pC4S4YSTfa7uIg
AgNLEudIUM1RLParUXw99jajSE7ETK+rOoHl6VP6JwNKFB3UODXQsqP5GAqfWmLmB3r97khcX+7C
VcnflJ92PLPQ17+5Mv8aL/3QdxYobjNybaTZ5AwE4WsT2hIcx/nJSvjqQtyclDaT+mDBO3KFXpln
bJ6jgjA2SXBbs0KzsdHAezWa2PKZ/CyO4ZhcMyRK5Cg7ZKk7V9NO5ZAtsSdIhNC1eiiiLGGuZz/C
B6qhGvIKSSXAcdvxem2kvX3rNAnOsVUGN41/9m7oGgozXJNQ+d7mymGH94G1rg+VhkZKEY252Uhe
gxodEwqbCeOpUMdYUy0l83xdUi1EU0lrwnZPPHujQ7ha5Kxw4tCN4SbPk5bcv/SmI+bc2s5420cJ
VyXPE4rj8HnT04kKQWtsUzScIXV+XAVzb+ESd8KNg5c4bNmDyEbGNtaSkIXx/mMhRW3uBuvr4SGf
1voFV8KM2Hw2hbT7RR7JRrBTumU05QQoJWKFhymooAdbioP4pvvNsZgDIJ3KIjH6g/w3eNP1C3/g
PRXfsMHCqOH8WYYSE98TGjiRN4OeIUee0Z3kT/9TOP6NvDf3N85d/iKtaetxje5lSFhsLTjdP/8I
JXX7sYBlNeGWhcmh01kdJUTYrBVmvP2icSEWF5Ud7cMIcq7hyrUrJJOugYW4boFotcesHqRO82PJ
oHQvoH599Vmm4WaE+A3JtaTinaD/c0ZFt6X/Ac4HT7PydgIlaxh9jIIbefjZVHB7DhvJSv21ZXak
YweFJTRtMzasiYRnjA7hgKX1Y1GiLbh3q91t7cHmxbp3rfOUO/BiOLX3uczvdkFOCsFd1wboy7Ev
lw/9hb9mHd0CM05UOq6Hd+J61LM+4zrI+5LERIO1MHZAanLbDlb3+lRv0P7BZKBkdExjR8aSuWg5
7p4IwxDElSwqGwM4eQ4b3OfPGXYGkyab3t7OAKvnDgmvb0/hoNibcio5qIwZRbV/G9gwDKSyULoD
YC1Y45ZOj3kA5XAamUOBElP5iaEmAbxk/WGtloOyt43BOOG/QkThlSEhZHdJI53yqdPuoNjGDWy1
haCssbb39B+/hu4KzQ3sWZVgni2BD04KcpDUybR+NKjpJCY7YkMkVkOtpfLE1d1Y9TnHfF9lFdKk
FCS4r5oPeAurMNp/8nbaBD0JQrXz9b7Db1jDBuDx/gNavcrkoZXgh0cvO/Eg8K6trw6J6J7H+cSz
h1y3VcpybKiiyd3nN43G3WOBGeqI+BIv4dFh77uWUakOt2lxJmoPO1QJIkwSuEvxlc+UHJTjrNfZ
XCWFfaQhuGQE6OIYKZHmc0t0MsdcLbFziQRgVkQwDXuk0yGBA8xP6taAkZllSPnWCSJGvl4ZqrZH
iUbyvzywSUe2UFfnu1mbz8Sv+XxtkLpRNq+VxFJnBeXUUaAywzwCRjKQlekWlcc7FY8z3OUbt1+A
qoN7U/P0j8nnca5PDjaUYpWOkadVIz5Jcs5D2FqwAyQ+JzoIVl0+MkGnNGg00A86RVMkTnwJWiJL
H8aufeuiAxeO5zG85tHthC5vavRQU0e/h6FcXNHXNSS+Ng03igGsrhNUGl4xXJYx2l/RKP8pF3m8
9ayVqNUPlQbDkNHVFugIUgExQE0pMyNLiG1jhPFa2DQsWMFNq/y5Km3rUvCF/ghxRjLGYTwW9HYk
UulwKKDthp1XFvCT1SbRrR0+cFgWN7rE1o9yJViLWZSMCK+n8dJyjHcDEivv5oddfiPE8zulR3/Y
x/Qj0Oo6S9wIGcsTdLvxtSmmQGRy/d5Czf4h4y1mHNaBmTQ90whF5kdn/u2vEyQDyPx3aJnAsjC/
roEcOxgTFzoNt39MAh4TUtPgMDCzuDnBKq3ZVI6OLLPFBkY6puNBlpfJKbX+QuaTmosVh//IGB37
aRFgWMng7UUMZLJL1JpU+lXQvkgpwkbBFYaoI7DPw8F3+X0UMwbKfE/n3SdNRtI0Lh6BTkwM6R+b
NPJWnDdbk3bZOwT3SM784tG1CJ4yJYbMD9dukrCMgkXFAsSoWSdGNxfDhJFEA/TGut5Bg69ip76C
Uaq3h7UrIY3xAq5LGT7PUsYmTkndBeRHqV8Kt/i21ngi4g/LTVFkGZv5XieWlfJinPp/yZj8Hkmx
rh05GrnR3B2O58FI2rYAnjyQA7Zr7G4TJX7bN0D8WE3GJiqOIagjR4NWsN2R6DX/FXh9h5wpFvMQ
fBUXSYOKrvNibfOjYlPFm4xpT6B/ue2NDTdoXIsSUisz55MPWQAEEILre/p2bXD6rbUXcwNWvts5
Z0VV8tZnzcAms2S26pOTt3KgL0Pphg47Z0+1amftr0XNz2xJc3uQhNA2fT5aMAQFWnPzTntBeYok
eKo62O7fLGqh7Qm/QhdL+vWK+ZzJQStfDmFXvF8HjR2ggErYzT4Sd5yQoVenlLjJ6hWaeVS5hm8q
05Gay19fee4inMYGjipuhB53uKVaMwAlMKn1W0661LJBAi/s3psHoSDCARFpNm/4gfhuhmF8wV0s
NtCLgCWPicvkSNW+WiSktNVWN4XDYfRQ5ar5vaksYS+QlSXY4Fjf8KwJwPBjtAxl8TKQn+NepzmQ
W/ztCdHS6sPPLnexOOReSRHSMpxzdtoft04WCqJOSo6QOvLqgHMJD5M9WDlIOubBgBEgZLTVXy0/
/sBhqiFWvTznPhAwcT1bO1s5x64U7/gkepoZ4KT7GXRup4t850fnSCRna53oBq/iEnj6/ZhV8N/g
7o5k0gYB5Dpo2S26rP+O0IByT8eEN1HtqYLRfGG2TtXx1GpIGILb7Svh1bp190MBdYCKreFyHJqX
u33SaJVJQiTt5FqrhChGJksMUZv2RBpZKzI3ktedbbVbqBUMZ4TihIsiQfZocc1F3otQE73YGZrE
deOH8f6dZTLucoyUf28voupUIdvPJLjyfZREfymsviP/Hpx9c/GNJscYcwuyJZvpmdE/gepOl474
wBXhYsz7AcjdGMsODclU16cIl5zZKXucGr3BAm3I6nvoOBp9MfyBJxTEva7uefzf3zn3DteKIco8
ubwqFh3eG9h5PWP8XgF5r61TN4lU4GUnrOBNDtV5p91R0A0+eBgD6iTAjh3rOipYeKXp61Kwbzp4
Z8BNeoN59QHHPt16hDkhhSEk/8evyHirun/ythNJ9u2d7ngtwQRG5uYa8TXSKe//GcgvaR8Ldw3o
gxYixXLNvss3vzKwLlW/jY9NSZpV3+1WBOWB+mJNZD2OKGv4MQiMMdWVWqnUTMPZMA81xRGNwESb
nF+5neRrAVIy4ZdgGLFPi/uCbZCQU0gn+m3EthSZZdeQf4qzMiz1dsMECORWIGbB2ipAKkoVvf7X
5RPsY7D8rCflyiNOS/NXrqVV9BA4xIAc5O532lGAn5xOr/SF0vrFMBUU8LuVFqSjpEqOwICbmal8
n/SwTfXi1EE67XDX/eiSqXR5PFc/JOwNW2VY1ZpmwmHMXuZWyZTwHMJlnCy5I77DeukhVUxRzmSc
rwzOfRcmzTcOCl1JCKVOAhtajlhSRrp/XsS1jYVNEzc8jYwCnS3mWJsWVEDbFmafQcWilYe5gyM8
ikARFTpaXj1GzQOeqByWBqiqA92iQXepWe+BxousLmBuqUT92VtD662zt8WNtOvlsvUuPQ/FcZ6a
gVNkymGSgQhFF1GS0DKz82OE4t1qTOxSx35b6ZfBwOJTfEmmGLcXZeo7ZAKjP5ng/UmvmBEH5Rzq
d1bsrWe6yxB3wvm/JD1Z9C6mPagx6FXNcXLKrzN9bB3aVZVRx8wlUWehwfmho1kOiRYES0mRO/T0
aGH404gU9JaXVN4+Civ/jsR3AKf+K6bjCDYWtC0dM6C5pOfp0hcpNRDnvS2MKJKG+C7ZwjZMrZlZ
XlGtQ7G1SPr6PdNaLDxaCjOmbmFmlHt3udeCupLluLtLZ4bNu6Kqxgo7ZFUmdSGyILRhNYH7n6US
ZZYsL1iYILx3/+gtVkzjb6UalYAuV/m+LnzmivLmwUMElh3fbgzJzcn7E5W/nHRwaDKDFmgEnRjA
iFCOBTqRvjNbGkNZhWKDnPyYV+j3U2emYUX92huB4/s83ZrcteJMyTSlMLS2PZPNtkuF2DCPCrmY
Ivm37NFaJmIaCU5oDwg+FmKfsQEg+oJ+awd9JpcM3LTriLXZsa1BRMYPgX/oceMfPKpK+hvaoTSx
O0b3VyBsL+bWiTCslPMdrzlW3X4WMJLkZ8MNrLx3Xzk41FE91EIycQRjqLsyhG5kJI1QuJIUlTdC
YPxVCP40h1RQIvNxeqvj6bgevn3bLHOEUeDRjKdIOnEN4J7RfuAqRIIDGbHV+U39A5sJlXfE6AM+
IG+ULwxNsZ5r0XuDeRR0BrouYmD07RhTeTj4vyyKAn3lu1uKlFV3gdYgpK85kYhlhbEnQAqlrNKY
1pplTr7fH668dDyezhhEAwbK9jva4q5RrWviDJ27iwUBfqifXuAk8JXGPrNBM39Kc08mWFegKOBy
DYd8Y8aFbyHdIS7HnUGL4y4o86vqxZOkHdPHKMdBCr/frjxo7FfgeAjQYuackx32To+7GhO3fovA
u7PobSqGEIB9BCw4aqK/RG1F1hfigkTZRAJIdBNgsHEhXF1iCipXl4jW4nXEbcHPhaiaSN+kCRdv
YnaCFVOxvxXvwXoCyDyCGPQtE67CWL/43mivkXxaAgd2dn0+f4dbKMXEXjklLLsDu0etaZF1Hci2
3DDhJNsJnADJLqWmcE5vWtvhZpDhSXRE5bS8d3zuvSDdoGg2R4Lb70uGCetKc+wnlL5Ue2b2A5qJ
spDJwY5SKvuaw+5BsDS+ZZ2x54isVzTJwHMdUwO49CGn2oyEiAfHK8gQtGghZwTwdBS2QVxQy0TF
sEugkF/3Eu3JK7k2GJNlSFzDp/1flbeES8llGmOBSTHEdrSPw9Dce1mkIR2CuHuKrR3eDV242PQi
U2nDm7cKNydM3StPV5JGSRrDcxpVP5pod1DozSgT4/xaAqoQzM37EKAEKng5qN0aPdpU/n89Ku06
xP/Qzj+LOqtdNzliGnGa4o/cYKq5+SNBzmn1hS8pGGO3hav4/Qu3zmUvuLiGjwl+yPaRlQygt1tM
GzsiDWUYtNFGbFYyuC3Vg33K1f53TnQiRoZX4UWnJfntkp1pGmrAY1cUNDjaguggGkvw8FOnwpOx
3Ix0/o1DJ+dcK2EIi531qCM0UZLthX0zvdTXL51U51wGzSuZEKwFRU/XBGE26eHzf1v22kYK2o3v
hjgOGIrCb8h66Lxd6c45AUhq5HeCitVRvDpe0UzjDYyBaekJnHxivQhYBNUVBjnyGfPB65hKcP3V
VR8BVngMOwUS9f2lUCO6BCPkkwEd4x6h5+DXBUpxHm8gCGIugPOXtoJvpBuvuNhbp1t+eJV7T9WT
1Gm9CLz4dX2NaUQTxVmczH4Wq0VR/WV7XYe4VxesGwO/hqi0mp3ApyuEzw/LpFUjkvZD/QugNqKL
g1+5v9DSuUy7t2kepfIVICfNkBKAVn4G/hhKmFit4vo3qB/pUDnKjUOd75qPoNrXXsD017zScCox
5KsvCk5VePyCWNNcEcwtV9kPoNPbFkDardGofVWjloG8CY8v99GAzz7+KcrsRrG+f3p+J80WcKJ7
X5VmpZgQsQdNmoM+A2GUe8guBxKYUQd3SjvwUPHiURXJr0j8ZVo/id9gORux/NIkiopFJ/IEnn7V
RMnWhXq878qttFC9GcqZ2DwGBE+Nzk5okjRP6KwsQ9H3xzmNclEztJ+spM3VKrHfZBhtucJ5oT/6
vs5l5ouhYDo5OlsPqDKMuviIaoJd95M3QqYCXkUIIRKWJXs+5dEuyKg3oR6QwbJFRryoqpQjcoBs
Hkzu6v2KMqTxtPYq8bh8ipTUXxGvn3SwkwaMFve+p7Nh0B/OWXfL+VmD+riXRESK8svOuwcuF73/
5tHSpNyDvf6mhZNd/oyeWxQcJm4DWbhgzJGRp3O9cXB3gY+qWnHB90kimVxeDlYvqaXmu0oDX34z
sOM1Ox8yf3UiACPpzoUQh7AgJgl+sT79k6ZSY5NTRyKXfCnwCtRaWjFqcnKjemRRbrJojEMl/PmL
pjjrUt8Gwk9T9djnv5K0XWmZFlMzL9vUUskuh34/D2K3Yp6I/yxABaYFAT3U3G+AH7KnLVmM9P71
hUci3fo+eVG9OysUOI6npozPBlNyCrJWCvD2u+BMBc4nrZLE59N5bMt8jVIdb0ArNFQeaBomUXz5
12isBQOfu/1n54Znkl8TuCmZdZj6Cw5SSW1kfzYe+F29REnjRpPjBpBwDZ/7QhhT/aRlNOvClYzs
0xl3V9/R1S6o1uUGugMas1tpbz0916/CZQjpkweFNAGBCgCkA87Gg5ZsxcVwJuPVtIkw9CUTXed6
EY4UpW4W1Cji0veR5Xw2/HCgYtnUf25yBWAGAb2fSuARCK2sqsnOHwpq6HfVvbahMcG46rSe+0SZ
GkdYFBwLHr/5h4LjTeMC/pU84o9x/DhXOKHCHSBpRru/mbi+8B6dOuA1InXTA5NEAy3IvW7BobBk
r2eG3t1AklLLnpZNVI8h+ePbh2oD6dWVf1yMnuY9PwzYNVPKMaR/Q20ikF53CJ5+JOaVVDxu7uS2
C3dUIMheLKZ64oohWLjqkf2Dmikb6INQDv/HB5W6/iAKgwulXm/uP3xSf1ME5cKG1y/IwDVC6qws
IqwjGYuZzyLhQyA5rSM2zSqYiZjlNKzfRgWb/4FeIynqP0ExiQMo0yE4FzV7JPzPnaUusUhftpz1
ZW8i8xE+NX07VsD9rajFYe38CBsbeoAG2IAQHWVZoilasfKpYiuhgTB0Qw7UCKT0kDIhgdGDevyG
WERChWPe8Vq5ZpntMQk48P+A4K3unOhCvJlV85vwY5cFiq6awzvK2N/N3gYVxRF4fgJ+9PW3NaPL
avrhjQgPnEVrrmnlkmCZdFYUnsN2/WrV6SMzeeHernaiI2AnsigbQfLsLFtIdmTV+GbbhLR/AauR
YeM3vkzm7wba0rQoYQ3YD1Hga1s9sL0SfpsXdITzKYH87DUPqs1TUf57ATHwY1lRJsnpN1eFIo0t
vqUM9QP5NXQBzVxq2e9k4jKAIUoVuuMn456BIrZ2bL05OuadzAaBdnxUqXLQhhTfeLIReAIMqky+
Vduu96zaaxup+Rcp690K5vj8N8arhz34Mm/HZAYIkGZXyhdZac1D+vjKXSiIyKtMZyJXjOkK35GM
8tzPNSBMcGYfD68zMGTrkxLlGDCepYk6ldNUbCxWGEInowX9A4yvYuXgNXFGqM1IKvaO3KQnNPVX
qPwhaMrW97JnAKN7mM+eiFGI4ABwiID85ckJjaARIi4ywpci6vr8z/PCOqEWer8OvietphMoQVPi
doITL880fJEeXZt5xcJGBEWnRSn1/4zl/U474GJKfpIQ+3UX0t+rcemYrJQvH+KsdaPHSyspxCvR
qb16XpjigYuUysJ9BwVFWSzP7KsUiZ80fL8n7jAX2/mK3Mg4r/wyKu5fnEZ2MUJtjpvgtpeLwgH2
f8HNMyZyfuL3F+zbmIYwvaP/oE8dJlIWq/EsEGaIO1zgl8zr0zm2kGPd1v5vcyViKRM4+26JWTA6
p1LlujIw2Z223XU5moqQ0lpGlELeoG/XzkYUyOB0Q8K2oTNoeWfiF3tx9PQlRXuVrAkXiXDyKr19
ssRous/4HNNzpOl/KDJq3+40dqvKLX6KxRAUPYA1+DbuHQC/cGzt9spZIn9M7nNqqkD5+QTwDVHv
Igok5J6JhcsOAmZUNELzIIaBwyciyZ0HrlZ5yEr4PsMrNpzCS3+jJYmiQERNpb2yKcdH6bblnsrP
zVvK+3EWEcx5fIg6tN7E7EHvxbdS6pj7G3wkTYyqwfczy/64iw3/zYRmRXJk/9TlTUfR25oWpN41
+RhHp+aBcbNxKEJtytHcvOHOpvDJ8lSYrV6/dxhhcykA8/5jFLmccwsZtc//YdRnPrgRivJne+9a
kY3pQQjZU0tUH+tZha91B4AEX0ZUs8rRDtFQwGt+yj0m26Qa3o8lNCvbR7PHMipTWf0+a1VIL1ka
4g+/jTrutNJKIaqVd0eGDWanNz/Ptobu9IjEzvHyTkkFotZgAgnUjoS4h0ewL2pDYPyBqY/1rJfO
ITWBoMkpwbk8VlhPvvWGm+CAgFTNm4Nl3htFlcCdZnquk+sNZe028zVIY4vcTFhobsYn4VYIYqIi
BFh2M+pfMHKchuOR74pSIXFuWqFNX+R4LamAvSHPoARumO/hxl2m0plsNJOYx+zLNw4VEcflR2Wb
/8iP+Rek9yJWtmA0KOXxOThliRY4O28lYTuzacXTbRlGTbXjDtZ2hGs/XLXO9lj4nSN0zsatql3d
tMJAzZT/ALuEtzH3MoKDXtoGBOUOOA7ULMDT4CY4EjG7/e69ZsYQr5/ul8KW1M4jVzvGN03vEX6E
JlyPoTA0Qm8W7X391m2xjAqAQdpXfGanKyPVIhNZ3ptlYOpgQgHASgPGgmt1JuHBA1m0fN+09u+G
zmLa6ErFINYbMjwoKLYx4H8PInNnlJwj62O3a/EpBT1ziGMAa40r5BruP4yvBDpU4gJ+eeuwAYkD
e/pldM/OJJUuaGAQ9yzHTjSMPx43QjDfSCZPJhMqko++mKkg4qfE1RhkZXHm+8URgPhIWFFXHfCc
/XYz0iUDRJ8zX8RlHVKaG+zX1JtT7K7gAzzUIiFo5/7UnZua6ugOzFmdvNaZrt8pmPAYVlBnOAkK
NG0Yz2NznuEK5gfgxx2hrJ7z8UBM3oTS+uOHe7osT4JxI28ub9J6oSOsdURiCKnPZ1qZRFIFzyPC
wVAa5GyprK59j+HzKAdQW8WJ1OVtuwln3mbd/FwvQ+AGShd5yv1CGmKTDy6Ti/nqGIyTQfdtBQPa
tbRJECzbCAHgzgiFSD7eGIf61xwrj5c+k91U7hAUxOZX49cjDBU501oGLWDa5K4HyHf0kpVidoki
3ye/jatgdbD3xfkLpkWKdBdHL0WL8TaPMlo6SYnTWUyQugqUVCLZg1tfbNRvN9d9wKJ2hw+soWIr
p3aMjmbUHeamunCYLBoHTwQI9PLUrEnkP+XBJ0Vnof/KGLw1DGKqtB4y7s0JqxORqCgT55WahLy/
883Ivnq45cvioDdkRVLsMmRQYFeQr9QDDc+Ecbf3fCROBqLBhyapqKGR56xqYD4OHSsqVBHqGeP6
v7bq4OIPkzOSsHFe/DKCvFdbco2lh4BsIMgCs2vkTJBAM5ck40uEF94BWM7eAdgTN6gtqnOtt27F
5BbJBEThfbdYLEg1IQqjov1g/jk/WplMY7SxacBtmBWq6HfbT1PYnERN/fimbzqtTkde/Hf8CqTi
mR0+3a+zvEt1k2lFHXEBFUhISUvQk2O3SYTr3ZwqdRtJNhnquVkivzh0yAL4Qrag3sjbR8xkf2tI
Q+dhlGNP4cOLnMEtb0H/s9txT3e8sALblKGgLchqmBhFyOf5HYLec4NlDBiHFTv+zQy3KqUGZ/kC
nSbCSxxhwGMUh/wqnKoQilxyDxhdohLd6ZV9/Rq7KyoINsBwcAG3qQ6Up9bsEvXTnYaFESWRukvA
7GZ8VdDEfihZdwyACxNlSrtgfxgiBJ7LvQVUwXpPq6M9S0DPrjp93kNk5U9T8C8/CZlukGJd5WFY
4eD7eIL/2cb8LuKvfQN6qYJAl/bYAmy6sKVFyfWL4KfrgovcNBQuhHJcI+OaiqdOi6APlkUKk6J8
6nASpPuTJUGjwHUsGuodMMuzZxQF+Lm+1oSFZlopvGEvjrJvzf4eniPj+786Wh0u0WZ24s5TUnQ/
yllioIZ92YgDnvMXdy4VtHRvd63a3m7680xQdxB+kIp5KhXM103lB+cgPIPBPnOd23v/eniVylnE
HnGWTDqH8R4NB7T0m4uOWhXFhnf7HDAOY/2mcWnQk+Q9shfYI/mkRY4OgOKgMAAmkuKx9OImt9Xe
mQFLG+gRxaMqsbQGozjk8g/SoOj/zkozdQV2HZVu/B7Qpr2jmDU5mnsbjyUP+AYpg/YRz4lmYpHF
GI0SzmaPuIiOy5zoRr9H13fs3MM4ds1L3GCGt0KLWqRFm4Ri5/r54KxfdBVojUldKClUWqTWNpMG
3INRCrQHH0ZK8c+n17EpAJ7tulTSMSuJTlPrAD5g9Wwn41LWNbkf8OkogKDJvZYyJbij4P8mEYZp
AyOlZ5+xRs1m+cM8O4zaBCe5i9OyzDKkE2IsxIsIJgc5QwpNpopFq4DRwBGoxEcBTHSUpHZlHNjv
Lf358xEeojSGp0E7cR0yaC3JjhApE2zBiQlgQVReo/uXGQ/rrgix0MJ+tXb8OKfE8xOqdsjvqAnT
Sx4MQ14gPVx9yz5Qu+LKL8AwhSgm1/oFEoxi5wdLoz52AKhtg7QuNMXQKoBWBC7BJC0NIFazsNrF
jwi9kKywU/rDFj/DDix+I3YxQrnsGQXKH9/1UsIxY/HvvrlifoZ2t99Ksbp5tRwwvdtyEwzzzojO
i+9lyeZUbwDM6ITrta/8Ro+4tyEwjjwqwfQEJTumM6A7xKpfCptlC+2fleOOV/s9nsuEo55BLeWV
fx5590SLMxjeB6Ril78YoXRq0E8+ST76QwPjX77gphlqzgnEGt7SalcbS1YYZxlynbx9SEdPH4jj
URH/alYQnnYBn6D5gp5+MJGRmIV4o+am5gq+18t5f8OpFqJODNtGIo8xGYHA9k0eGeE3Jx/Ey3ce
IVt7ZUWFOilqwBVrgINDB/ggcRr1csFV7vYBW3EZSHKqoOMqCNPnli5LTRtg/7nVZM3IIVSqSGPH
p+CuhsPjFBY/QjyESR9p+JrQOqYB1DVL4p169B4QgGfbNQZAAUA8SVKjpk8xQJYQ94BJUSUv83nU
9afu7G4nnDowTNHt3Ffzzc9K+qbokZ8LhrlIgUWNJPCyiJ6s9RUwkEKuX1D5ZuuUoq5+sOc03Xba
U5YOxZ0VqAwsVAoIndja/TsbEUqvWVw1kwdSgAwZIogzt7hyt2Tm24MHzcV6/wfq7csIDYxjGGD7
TMDzlkFVHmd7a7ft8TQH1ByIOLLCXPC1m52h7tHzNqu9hPvsjE/XS/ivxl5soFb+3dDmktHp0Wyn
M53JtcP/7ndx15clOZnvDNdEuDKOeoVIVt+yl2gtklfDrm26vFzLccrwS1abfH5xlPPj9AFvJG+/
GNEf6UlZJorS+DiC2dVcct/RULqVNXcpuG8ZR7R8eK5mg0d6prHDXU2kxOxdPdakxMubRODtA5Fr
HgNGkGv9kufoph6hirT8ABTTWoDV34CTjfhkAE4frOUaf3+pwr1tE1LqjO5tgQ9/MliMmMK621W0
bWiUwd3uGhjE6ynDbvWaDWTIYzk01qYi6RWq98vLCm+aHhZJcjCzRHrsk4e1wMw+ty5OW9J4YKL7
BAEmiTiibxpuuRL9KuWfgUkcyCmWZj/NstbKXnPAo1HgRstbct3aU9tGBKF4C408TsxPvRVzxW2r
Op8jZ3KuMX4T67PGza97IFMuWOnbcaEtjJcJnWV9MSxt8z7wph8b/NjNlNPX4RviDnOOQp49uS92
+pLysLwrsIYGRJV5mduqqcXotyuzfiR8tP9w86Bf/AyvkO/gIQGoWy3KZds3tgFU1TEQ1DjSSOTy
6xh17PlayHjda2bzyAeyFOnEsqLaavxjY1Z0EmNIpOzHfZ0o5GxuB0L3Xd+yMv1EMUNTDZ1z7q23
Q6y8yELAsJigIFYG868OqKqGVPwt1U0KK7Rsh6FvQ3A921lwRER5lqlCNL20LfyrczZqpmuKuR3S
4IrYXDWYtPiX6YaypaWmyIo7ZcA5eY1RO2RyjIdDN7YLIV+L45zxaixkRXkJaUy/RA2iPyOmxZNG
uJAk9xZ5EaSa/Tcdtue49hvRrQkf9y/O3JS3ncnA1w9kd+XUe9icqNvDiu75Xk+czuiffgvHp/TT
EaUt9/6WbJ1vZWCD4Fwx8p80SUAyt43uwkfLhKoXxMFpP5//GjjAe/CysMKEBSkgPQvHprgnXDF8
OrZh30HC9OIO6fPAxXJwkvTrIvS9XLYmo42YB1Z8qvu1ATtEFkWrUmVal7kt+dWU40WamB6MF2r9
M7Rtq8EhmE1UO6inEPW1TwGSbukYyIU5o83BuJJyAoawcvr6WNs5ciG1gITZEAwQ3bwwb/zfkPqv
rD72uYXxx5N4HM4EwCi9jycpFhxpTf4jXKCaQ4SUbbEto/Sa5OdKHjffowdMaTbhf+qKXKKbeTn8
CvRRTlNVmoaFCM8m0TnCLIKFhQAzxQrC4MDPfljO+MBQaXFoi9JecFD/HjMnEXxvy5BFi54yX0OC
Shw6vMBTzwMYviRnZXdTq4/4duphTFA1z/RpWngup/0RPpMoB3YxvMCGCr3Hr/Ceg2V3x79rWkTB
wrUtCscNeMAMgtzSNzcbVTRS5aQEvFV7erHfAWsrTQjuYUZaWUf90J60RuY2qJPJ6qsN0OsSz/Yp
s/5bpJNjcXy1k2ztHmH9ZbBuT3/lFJYdYdO//9TBU9FmE8JEsDZfQDr5rvawd932VMy6DDGnMT5N
h724iKzmMh2u09lYbeHKrknQnHya2M1p7O8jC+d9s3ZJrfgr33BxWTDNKiLWYJEvbkFUo3Nl6+Tv
Ah8ON94mI/GixHUkTQxltelhWt8fwZYcaCPcs5jrn+NqrBY16oKbdjAj6RT8AqogBFtrtcOdXXKd
j63SdCs3nX/WRbD7u7PNPCXVsBOobfSJ4cbLPCLiQY/rMc6lqBh4bCo8GCFLQ9A2yYGOs8iSaECm
+LeUwliKBUfEc/sTk7qJfN9o3A+n/XPU5InpMNB2KvNhEHuxy1M4Y1DbnvWpa4dlVTwFu4gzOmCY
k9kVVD8Kf17mgg9Rk0uAxPaAvhsZC2hu7SJQOB0U51jKX10rDnF0n6e8h1izncvH14wUGKAPoRPL
sCj3Gs0MlW29neNiRTmzhxXom+tp534tGnBMTIOmkBoUe1oyxdzL+bvjgbFOAKLKc/IhkW9SwGqz
m+YZojFqXsNmgb0EPrXZqyH7w+sbegRJlCyGaXuqeassKmcmjciatwfxCqM7OWxrN9ZpAs0BiTXV
mu+V+QCBSdHOwkSfUx0BdohRsi6uSjRaEuRJRn0/Be+4cwfr4Q6SpcBJG3EGrfmp19Pkxv0cRrSG
a7yyz3bwcjC6AIJ0/tMUhlVK9YGNdRMWEBaAMxf+VVkKMUNd7M0InmhsnvDhpStTU5JIoVoi/jtY
1tzmyqKDi/s5vCP2qsFmI1mGMnwPmDT70DfZpK/0aKJ+uJYJxBBNarGjIul6qKuiX1oqguFhAeFl
nxW489yoDB5MfxV7Az6yjx2zQLZ7fcFKyAQKRZjnwW0+27b+xeEhUSl4xR3HQuuyams8mflFtaQD
xmmb8fOa0dpQ7EglqukNaNM39+eTXCtLFNj41yiGbp/bzbBIWou85BVg4UHOnTxzz7zQnsi2sfHU
HqU5WWiucsLz1rkWoB4XkWyqnQF9BAR4CBSRRS2hNVtZTQunGtsmTtVxZK7GtTJEEx1fBWdWROI3
QUiJcFH3OgRQAkFfc6h/Cp3vGKvGwfhPIhu+Qgh/tHDxZvNJpnfTvqy0I/XFq+dxl5V4cL0C064Q
O8n8pRfF8OPiR+o2cMlCpoAB2NhEY/urZch4e0OazfUoUoMyFK/drAve+fdnWg6EyEnlZqVRzxFW
TbtfPyqKOT1/oSsVSRrHSkUri1sGX4t1wwMN0ojf3pHRVhvk5Hfvd1WOC4XAJEI1R+RIfP0PYHdc
fcmTVqrMFmRdgnQzDzkoRTOYkxQQQDulDwUi9zhATJfe0uFgKpPmg78zn4RYBBrn3vdhCov5WlDX
0Fe2RHlm0PXWVqNFkQe/UsYN+PAY7O4HJxHcCSMeQeo+8GW65AjAYR4ofbxJAmEOc9EIcIrWg2/P
4qjwqYSt8Rxg4XdotiLpCg8KINqIlLvX2+Eroh5cN1W/phJak3QAgFVroCd70LGoOLfXWKN2v2gG
iAgIic9nKPlMos5ucX2a2FiB/Wyt833R+Nz5s0PbaYGCTSOuZj50g3zNNuuP0OJ4BqfAqauxhfdy
zvzb5R3xP50iKl4PivDj2g6dNd1qCqsXVPUfIKEleaDVcZhfV+8jBgu5ep96AAbdxbgXeZeYuzZm
l23CQJ/41QUNedqdnjRqr8QrzWZub3f6GQGi9z+0y8TcK4JYZPilVRec7oUIOzbnjD7psmI/apSM
zQ+DHGK5dFZvYrpJOYXI7fOyYmZXY+WF2OU8o0EMVM0pE3DbCVXiiTieVSrh1mE7sJ2gx1puUqjJ
Una62SB+ITIbFd3oRv+1O/CL/+7Hg9tUFgvVqOVC0VJoB5nz8lD5dRarSXop6ef4k/csNS1ASvTJ
VFmev87qFJfPt0zBBNt4vyMKOeeLywC2O0IYmVXMMk31m5yfQ/e5pK/MT7I9QmkWXQL/VJbvciiB
rNAFy39UdVmq/H//VvLNN8TRSyiGiPMcdF07EqzaKgrDmnrCdvNlvVzWRUwHz4NtauU2BCyNSDPs
ly9j1tWvgAXhiFpw84KqnE0mUHbK4cOuNJFuGM4wvqMcGKd6S9c3FWVBTURxYS4fk3ioO2pjiFD4
Y0hk9k17lnXCsXZf9lQtOh5wdvemoCO9ZYtLXhIATVdc/ynMsnbhS3XwcDxJCvbuqh3Rr1/uHXRH
f+2DNxUk6/nTpaqwRwxzEAN+7XKYSjlk7WnE178b/SULDlzYCim9gtwQksk6C4RCtJWuQuVmF1R+
y5PXqLWX6Jmy6iMsLMktpNgaJlN2/W+IRTZKcVQwbpxMmSl4WH2G54SOC4/+afQ3XnGiwZoMvnqL
Ct4yKEzDaKfE7fyO4CO6KnZ4IVtVb3UU+r3CU6w9kkTH/m+REDMMsJpLYU9kL97so9Y+2jipom6B
QGG1bXHPzjTKZtX2LPndFLYW5+8vz7RA0TACheuyE5pIE7HI5N5bhOf/nuxa4w5s0lzYP3cFHtAA
gUKUHGucciJt0wNe6+VVNzPFsBKFARFxZJOz0OM+HXsL5+ZOmj72O9+T8TQ07KKG4ty1C3UrTLxH
6qZzNpbcYvqlavrv8cwTzQGe0JL5HE7FhprwJQT2N8jBNTP+jse6xMpqdwr9ogbf4SLA39g1enEy
DRYCmmYaiAcLinyRDGEu3IYOZGhVcRO6fJ5XKORg4OVt/oeOsq8B72jjDN2iipE5TgFtZwa1qe0k
b9ongDCURJ/xc5Kd4A5A9ryS5C1FxPt/lyx6kTf+sxtPpaoZULhzUDGg/4jKvTDJThVcinyO9oDO
HaCSUja/xkTgVGoMCxhVkxHw6Im0qbhwB54u6b5lltLdSovxYNnyw8Dxjm0inwJM/cK/9SBsCiYo
A2iCc9V31efimBkaV2lOKRfHLTmef5w/4YEIhOvID5e5YV4xPl6rhDRdbhYW4jCQ18i/rmZb/OxW
I+XjfWFvIOo+MgXMQ34k+B8Mi6AnZLL1ctr8NnslNXlQHccat483ml4+i7rlpAcIRaq91gt5DllL
LXFUTU4wvMaRcum4+UwdUJdLyfQ5MqXxaO28lYnQrpzokdHFMruYN2zbDK0nJbQ5hrle2eJWnrv4
86mbepN6xTgqdRedUFPhEsAwJmVCjsIMAlIyuBBIdBa7dp/3PCxJ0xQtA4PluX851/DcKvxB4dpz
ER3KiwKROnkQr0JaureYsTsm8oapwZBiR79WNGkXyt6ugMhS9p5cTqltyHyRvsfqtC/WX6bk/mnf
i/TYuzYYbl6yHPDQcS8EYLD2zMUHh8QoG6gtzvIJceIucBOBiWLb/t2MA/zq9MbznQ7JMD0xsBEj
eLoQQeE/rXTprBqtLMJSdRC3a5JZFgs+1JRpyCK/xOqe46rMutJszTOJ7Df1ednCWemLbEbant6T
VI6A/nbcrPTKcFgcdp2YYAGz7XLJCoBl/DXzAirxVcpmepz/aBFGM6DIZBLPab5rald3fHms6ZS0
5Yi4/T2wqtvzglX414IVL82N+xe9ynSGAr85rinv+pxoC4YgS0+kqqNdJ+JmXXcIIyTv8YNhsxhF
gWjkYL88yMjqnR3C0Ap1R+M6c9YSe9OX66kpp3S8jNX5btC270VaD83mdFZF+zR2jzcBJ3YOjrwC
lyn227puOIPsqOG5ojTQ5oFNi0f6d4QRElJTofluH0AKTTFi5z76VTnS6DMck3iNZNhnYcSpBBHU
uM4FlhyWRw1HoiWIqMWaIy+TBfolC9NoFDhwUlQW8mbJhK1DcGwemYYL8Q7hLI534HaqGUpIJmPF
tqhvZIdVBw9v7vLARL0rM6V2ShJti5pPH86RnFHZzWPAhCJm8fF+u+s24I8yvjFj+xzmGzqSFrqo
s4KOkDMmLqSH3k0RKH5cY5BgckE4+X99Nsm2JHCI+N8JI6zflKlvq3UZGcQLWo4MLM+S8Dw9wNU/
BXRYB5DCc6Xj4mLF4Q2ry2nyPqx8uIBlV7Fxj0Nz7WSyqSKXrXKd0+xfGVA+b1OodMaugy3UVrNa
jGR3sJziYcNhqonTDwDIpuzqSHsXMNbOMBTNosIRpCWUfS8LqTA4O64KAGDODa7szrDSsiQgD5Fy
KlIoEpl4NvhHy13aFz40lRrJ+W4D3IH1K4yNnAnc4PeMNq8F3PQjF8hGSbfUpMaHP62DgmtQuWCO
8KqnLN1cyD5W/dj/F7xejH8EREk95JjkmEA8ZOPGXaXm0jX6U9QApIhzFIKLFZFizJ86wlW0nz82
rT2jqM2F6/2wQ8w72AeoK19vMqZ7uVxlCq23aPAMzKKAqD8sXWRgDkk5a3xtKRS1YliwoWFFvd5L
il0dGZsLD/XZMprcdViEeO3Lm82LtXMpwE3ZfL+3PSw9OVQzUXHXToXA2V7XHmZc9HfW03khFWQM
kwzraz3MhOk24qSQJHsg5k0la93fL4YzzNgIhwIgf8DCn7FNFbbGCNbzZVzLNl3DWAhLfRds49gd
xVFeyW5pvnpYuKOzaZPdoz7D6jco8XrObJY5/pqW6GLiDvdz3voqOHCyUdy70vUr5TRXdu8el4MQ
WntWWHtY7KnlISmT4bKCMGAKh0tJJJ3obhKV9sWSXVbgpORitiS7cUqgbr3MkIjCerqpVT6u+j4T
x9sr6TdF8IVMyVgsBQ1qzfvPBmtrYgK4/FA4xaBUmYx47QZM4zrI4kEa2NS0gk4y7mozHBa3YgoA
wJeSGwKYHEz3Ykik5zdpUYGEO0gOu3bFdTCIw0oPSEu6tfmktTs9t726KqA3yWrthpwAoL2dPfMx
rthl4V/o6b/wy7D2imKWQgBA+v1KT9flzDKC6hw9qHf6eDXOL1iHMhGnplqOxTRbpy5lbD3S+qpM
sOhcPodqhZbxgwGmp5DCMHcgxylvhgzoWdclejUv4+kGTYvKvuR1IxgejHQRXj5EctPvE90opWoF
2xGsZNnYq5KxOGWhhD3aIYoIjoMFCSjCx7ti9gjoVgA8WIBdx0d2bX9smZG+GBIy9qQwfkYt2Diq
i+0585P1QYRRvU95TLzRMoLOP747jxBrWkBoCVCdyyQPTluxpb5gz3ZvKrT0cPRWsZQxOvXMGj4t
2xWqJsE45+VX7iTkb76xSKE/b7dMyt4S0mEnXUJZQycBlfnN3gLPgK6cnlpOyXJA9t7rzLlChHh0
e+84BsffeXH0fq1KCOnjCbtdgDMVsW8jScuI4ujgM7P1P1uYr2VwCNdRuVGvqoSZQi32iGmz83oy
NEx6j9vGw6jJbqSHBNuZDsX/PZ3fweJVbhrW6lpu/s4j3wSQm51XJomUZweETVXenW+FYC9RbArs
aRceKq7JRAviU1pmTJfv0BEv5zaMTu2iyZE+3XhOjSfPRp2RPs0VJABZcyXSGr+bhJg5gIaZ2pF6
Ydh+VpLCCmoMv/i2dwtJi9jRUs+lCRLzqGdsOe5adObHFI8DImOzwLA/FUy80frBjjQlsAQybLmC
8X4WhKZQa2Gf+uE6BkZ5QoURjTNzjaQE7qYUtIvwlawREeKSJEcLbfkeZwFBmnlN1HcmJTaV5ysv
oxx8hPWicosFqZmQDtyiHUMpIVGfddD48QPVpqIdw5I6OwwEd3aWP/37dcEQcPSwGp7sTF/lFM4t
4vypbBxXRdtrHZedXsp7orvPve3VpwZZTPyReL7YswLWo+1wjBwFd6VYyDf7wmJWgxzd+hCPNGaR
nDwwgZGR+q9RILPPU+e8lFyqCqT9cQVEwzWdO13mebADpVMeLN5gA39iTJTetgEiglsIhr0dcIPk
r5w+WYJfca8dN7SHm4G5bGUoOZLLY4jT/QI1O6GEKiUeyulBUk3ByW2xdNnRzEgX/Ntn+fa4iFqP
Wacl3Q3hwmZdn94DKp9NRqjIy11S+0wAWhsMZ/HyZSfn90GL6wBmenShYMNoSONT03dwl/LnUlEp
qjOXExysagEacEnjc+GygU9c9+l8M0TqvtQAis+lpfVN6FFlk2FWBZap7Kc92EbwEmA/mJijzOSd
pl44uuPDCoGcwFqzfNKUdLCfcelIvDGvHvfPfhGXnRBA/wMdxVEOrQqGxnjn0jQ+UzpqSVwj+xk8
h8QaakA8uHYq1DDE4YzlfWSy9lWenCBymaDceBhqEf+rY1baoYzUcLswclzb45tJEl4H02psY9EC
hhggL6qQ60hZ74+30LTW6cA4L5LJ/UgGEYL7QEhNOWMxOpkZN/PJniBUd3HO4jST5D/KMpNFL0Ak
DwDtB2qzzbeOO+PlfqISEZXBdK3LQXvac/SZBkXIPCSnE1x8LsnSNsgmXJYJqyH8Bk84H54th9Mp
nWSn3tMbulu588yBbnfctKmSyrcw0utSoFmRr2Ti0A1fSqnmyqAUTyfB5P6/lojXqBIxzjP7prTy
4lK2l+0ZInIEwlZAZnAzF4iYgM/vZ4DCVjDliodciEMopWtFAfnQOI7v8ljVf4hJbXFKc9bszxkA
GJ3tXpzwdtJP92RHwlFQTqfm1mQpCdx3MctJis/Aanxyy4Rfz8Ip+c9eVsZF/SdIXpsFkv7T8yK5
XyXg6qFWLJmIW0j12L7XF3TDhePyRpkGpiDWguPqG82UjRAhYD7KC2ZvXWtOnB12Une8eMoVNdRb
gMs2M8tDIdQtKC+F6fQ3Z3YOxGQwdvOZOoO2EsVtNFFJJjHnRtRAppJqau2Ll2MfJqMhy1/fA2MR
IE4vT9kGXMpY21IsGuxpnbDjsAcrO5BGUAyicUpD92YtqZPRUIq99N7rXaaYbECjyHTUAH2qjiVO
2r1z1xoDHI2HOpaTfXU8zHb9d+KPHcr5ComTevtF36f61ydUfuQEHVUfiVUIy+rewjHeS06HyuPb
3gaW7pAajdqUDAMkR3sDkKgEUqkWz35yM+D8lvXKA7rhPRpMgMYmwmJ4w/jMfs/tc+ygyBzePrGO
r6Y8LBPWIjiOhIujR9rBFL7NQiBajP2SLnrLUmkiGrD1Im7ojCGmb2+AO7DrcCWPFWLv6iVh0k5a
/2K+hSMhqtf6LXy0zRKGxzFYXVjFpPv++WRzTg8UOIAQ6Dz9BJm2fON+9a5QmtO2RoB4obUM6r3f
Qj+zQtnzCZw2Jbc/GKQegfcoNt8bIuNWSsiTh/waYBynDCDMd0Z9rh3wN5rAp89zg7g+h/4zZy1V
MoSdVMgkzeMNbh/jforUlBt42wsUzZX6Q03iLht1S44FjIMrnkbwuAQ2XW9dho2qg/yDkf19CzAz
DPyScKwl4zcK3wZTbRigbepmnrSAnTfSiJTTF5gtv1RZFgEzsFjEIIhWxLc3iAwZFupn/4qLT5Xr
OFH8rXs3zqrW7XrXh5ulAXAB7Tpu+AaAW1ssdLl9HbGSDmVXTwjr6f786CkAGyxsps1P36rozTcK
rDPdJWfXDctpv6kNi0Q9LPobZ5i506c21tL1SZjkkcKZZR/IU2FjmAK5bqNDlF1m4jVfcUwsIlOy
nc9e0hammItR6QUW6AoQqXjP0qZdRdlF249wrrXEIxEQ+slQKgVpcp4Hg1faEIRPMGmxMMZwURfh
Ww2vyVxob5Hirb8ByE6kpnwbBYxJm5A9aF8cvoClNna8yQdXr6pm0WCWqpafSpcUyt7+x1P73K0D
ticS9jAGfUBugYg3ZnU2x5HQyOYCjLsIfydKG7UjcrigbNsAJ8G0ehBxZBcQSkxoEzaQLs6Zwuyi
QrEqlmvtgrlusdA6Ceu5BJicCs7FDOuIe7JGO7rngkJgngyKr27Cd2W/Kj6EHer27MK6I4O5WRP5
lhkxK46ejS5NZ1VSL/IvPjH9msyNjO1uOlCJn1icujdxVL3kNx/4bMbF/NVYHGibvxVuEqn2juxI
ehHJC5WLlrae64SIr67s8FTeYCmW1FwnreQWC1YavGwDrhZe0nfxhxgBzGNTf8wxP8PC7QmLvI4e
eOhsP6i2MXC9Z25EDV+/Y+7Y9+c6dmyzIr8ja2oTm+31wXkvAfEj3DuVnLZW2ez908UX/iAInaz7
Xb8lz1HU6umQHtyv9K/Zdve7+kIIXOktxshqdmHiDfoGu37XK1zPC9e+bZ0EsfXerYC4wHYHpg7M
p4Sqx3UO/DESwCtDCiwXhY7+aF0LKq5yJdMN4MQrvPMWSRqu3TWAMI23fBVxwuorkrGpZpxwUfbO
F894BWqFksfZ1nZrUcJPDZligiUBmuiP2U7Q35pZJ8pKeIi1DZE1SQCsXuggPpytfVXyUQdAPnfh
5wTakKcQUumh2eeaTicV9H9GceVcYs4ubDZohBmmXms4k7RooZtqLtwEN0Cn9tUrBFC9jHeFxVwB
QfkzegA8EBXrGt/TJC8gWOuxvH3o40LO4rY4c4+3HouOXpXMSvbNuzkOjljR/bbeVwiuWYNKebiq
TIdrNeKZujJxrcyyYDn0ZDtCsRpFjpkBAuW5vdAj7KcSgY0wioNZNqCXUra4XhlbMZxFe6bI8Z+Z
SVd/9/dfQqPzgrPJ/lVV4AnHDDzIpDRZJZ/kWw+DYHqn6Ly8MvSehUH0/ajY0uhTbmhoKmiNFj3r
rtMCcA5Qr8CFQlAyJEkiVMEwkouzxGdU/vjWZdwFZtM0vOaWsXvD7dlbhdvq87fYhYQ8Zu2ajvtT
QGAQmQmoGe+cPH1g/iWYlJLsNMURuHDiua13RcxbTGiPEqWJLEqPzof0HtR8j2FYLvFZ1F+5OYPv
yNVYQy+iZFqf71iDuz/8+A9OHAbXhiANOrA99it2qcaR1k1QUBPXqBJtpXM0FJDoka+ZRFjhnnAw
Jzi/sIgW2cDKe3Affv5fE+qk24iZc4hgWkpmw+SGlflNXscWSWQddrF/OPHA11MdC8YoHxoGvLl9
7GGw8ZpFTdqZyemJ1DcPxvPR8T2/66v6n6CmS+3+YpCR3euu1PPuwxt46l/xdEWiUqdC63cQZCXC
Vu562281+UwHRpY2wqRvz/SPoRFevSx+t8wxNwyCULKFi8bTkzhZjgy0ApmdmbCu4YXWHFkMK3/W
OhTJXTlou7WzcCLcHSZJnII0DVa9gZ6hkgpzmxJL0o9CMV7bTZQx0oZVWpapgGDqumvsE9iPtVwV
7Fx2cXn6I0i71E9lbevwaRGidxOn2sQR2Z4ruFKKeukgzs01UaRhORGG1ctLGY1dtV6RFb6vMwTK
ToHntWwOyTA28lV+rTSNXu1kbcSzyGLxhUajHehB/MiXna4jDooZOy7bNdrbj/waCdb4GyZy0XbT
rAgV7cHSmVRNGgCSINpg9yv9V8tX+XGFKXmZ1DgtK/vxil34QcaVORbL0Ufjwjru+637/p4PTf01
1JCqqdWfx+e4POLHUxTqAqZHaJhgHX9o4HNbpmDwQAepg8E/oYxTHNDn6hg2cZQwrTDD6/XNfy0F
02zqsu9OWsZMG/9cOxu2uei2lkYIbvtWf+W42hdAkFZtq+HNztQ2VI50gatgNMUlXVhA92mpvn2T
Q/6GwQLE7qNGyDa+VOhfe5j4VtolFCAKavVXwEEdx4Kmfcd3WM84kvLAar//gS0RQzHQQCLt85QP
7iAA+QJ2+nNjdhR1wYDBApMmXoeK8YTXpQO7sRpNZskZ1TTHiedIA9G2WCv0hhxPo54NqlRLSLXB
ChlAQlYelilDi2ewz9lRZ9BkYMItMJmOuFZWr9erKS7LNBNRW4bLeMtFw6mssrx/jT+LdquKVfEV
5yUvY0J0M2bCbOh5zuA6ZnwZQOpIJWrGbbuHrlk93Gwkg4PafzoIoW5qGEMSFuJ3bDH2Sds/jwH9
4NolrljumDgiHeFpjdjdQHlQhVqzKX1ajT12S/47mCefCzPcfspjEPGCKUPS6thsbaZ/gzZrCQ5o
qk+sXVyKlEhQJBjuzQBoECzymcVz/kromYUJVN/hblkd2KCHan5EnV8HToRO7wlmFuVliwMV5Pdp
Lvh1rHerg5nfpo2h9S0ZyUYJaRG+wJPbgcgjB+h9SpJ9FZZOwvEnIIV9BHHlzkbOc5b3l/KnlrRm
Wfj7OAOWJndLK4B3yxpoO95tesKGnqKGjQs+8YeHqBgxRNEGaM7jC1UgMb11YX2Ba+kd7P3nRT87
Feg7EFO4cPsXyf/54jeRV/hB8HRYlFr+/mxYayokg7xIPdjX/uw62t2hQywL6YhqWEYsRX0nCeUa
m1BNYvM0TaQnLgZD1k1o3tPZQwrx6Kd7Y0fSmSpo5Y9NT8eFnU6ZLVnK8fdVh3+pS9vQQJK3gkvW
KBHr22SokcOk5r7lxWuPgRMi+2pA+v0rsM1v4wivn7aQSgCgwLn5ujXjyvZiSDY8TctiCjVcEuc9
H9kYiMLQEtpaJw80EW93Ik6IFFQ8uF4U55J84Q+aAOArX2gDEWz0s4Qwytf1EMdNlt5zEOQ9Wsj2
RKNEl3zOeDX0azBm/vZ90ZuX5WFMhS0I5vZLuElnRox+qm7O2qbW9WhZFl2ah1XTGY89I68PrM1F
vKi4qylxeeC5iCLNdhgNx0QgmvO7Wwp3kh0TZsduo9LT79nci7JA93gUVGAUsA1LwcrS3b8IC3HA
MiabVFycX8ZC2pxH+y+5POYPzNd4yNJFCBK3lHSTgc5nki0/Jym52rFHNM5mV80YfCatIlPnxCdW
OvxbS+8YiYmMEB4ig9DSmUcH6EW7R7THmXkvM8/qaGBvjNW7r7P1F4FicTfIhbge9yY+OQBwHOxA
TCKUQOeqVBvL/y8h2n34U3HNuJ3Hfb/s0muceGmy5rYiZukwyZqhM0UNAHIbMMeUkIC9pq9dkK8k
HSVIkMV4T8uh/0Mxa8ZxcLCN9LeAY1d2fY4S63AG0Ok8oOmHQ86V4zTiCXMOXS0BCJpYpFoZhVEG
P7JHMfRvgBxPOSc0vOoHDIP0T1tJt3iIWGEGUSkhNSpuAbTyG4W+DUoCUJaUoTbL5e8Nda/9FyCj
TQoYosW+Jr5nNOlYUHCM4tlkc8PJSoh9De/gCpURs0Jw+Djt/qN/j3lztOmVn4rWS9oBxoXOlkVn
poL1EwdiBRObb5aoGrAefnTeQvKnGbeJvXydBlv5/mGu2sc6RUImu1keI4YHR/hxw0jTEopMl6ni
x1K9CKtV1FI6l6xLpMfhW+NwtCCHDV4JUqL0q5yoHCD2LBEmNp2JVtGGzTtA49mLAt6v0HaB6JDz
/MQTwt5Yfdhbzu+WvnSVHx1IyOR29mHjBrUtnMA+w/wkLNoKKX1OfzewACTJ2EN5M96ASQioRMp5
nCG14mYYVGSObGIDvIza1wrYy41Do63lRLK5v0q53YRZ3qP0zJeaF0EGo0LXg9PdyQ7S4fQY957v
fyzsnSFtGO5VItzr9ad4hz1LcDEsconX9WnUJAC6MxupOvrIlpFyccqwHuXnmKZzNb4v4bbfTLrh
D9nHvqFs2iUlIrpebeQd+AFuoCAUiy9WY+OIe4KAWIgk20yrvKXww3ZfsukZ8RneZHHleSMPnZKT
ZeneV2vJj9Nm+7ZDmwrWGApPGAjiSvmYfc+CzZLxa6EhMWkid1UkhlUg3VMOh9SSjTKa/NmcrZkA
6SGzlxAOIZWKU+1r5hKosAXoTVNH3lf5y82Q673UwMJ/30bYC9ooRvhgr75mwYb+0ig2bPF7k6Vx
e1qYYkC7LtiDKB6TxSTzWO2G4BtLCyN/n3v8NiyyzvFMshfhu/82aYiACMmvywOOrxIGgxPTO1AK
gYb7O3Z1bDD5isMwU7IOHUNBenyM71D0a0xAOdYZQuqEILSq3PLeder01WsD29yWVifETW3Rz4RO
cBHvn0LL9vb2MUGjRxLyDmpVqvqMD+lIiWsnTaQ80hAZr2Zx9wbRPQWV80bM+UNgJWXSaXlSA5UP
plzDKGDgVacXk0+kDYhplZ/fWjBhYHbHGUtC6e3g8K71xX4HJ5dGDYRls41iFzBOAVVmYlDKVDht
X1rg4qv2lLUqQ8S5DpSU2YOMV5KX5tp4RrEnmqRtJb5/kEgFkEbdVBtAJyKvz+2Lll4IlbWQFTMS
38KXD7yBkQZ9TKbrif72ua5pLlsdHIA78L5E2VGh31Oz4dPQzOrvz3DlTMGTSZXbjWYCSiOV0Ep9
02lJWZF0yvDdauaVWzuL6pXWD0yKpdXXK6T0m61Aan+5ihGcfyyKhcQo5pdagJdU1n63KFh98FFi
+shrEa4Sd4d9xiXKr9SkioZuMXW6rvskm+asHjCw8Sde92CuFIxZb+L3NR09EEdynm0pLM9Z1flS
RYA4PFVlRX8FlgcMfUNILKvsFbBl1Y3TfeW7wyCBbNGY8IAmkBKvvl2MbAyK1JIKmbjqzi1Ph9fW
eY0tWncP4MFBeyVQGXr1dfEKTyaduA4ieuHFrRGrcImsz8HyvPspMM0xjqpiMkKQmCGdkaIhYaN8
x8/KiJVRFYlgsuHsvC/mZJFnhKKuU5yPriHV/oGjO7KX7E9MguKuYr9mq4yDGEh+rlFoTwT9Lf5q
fLtA0WBFmoSsB6SdBWfPjX1PDpXKl3Eh/06lnwQdGOWIItIW8aeXLb+tbEEWbKC1Z/TNnrUic8YT
/u+oF0JDTSAys9xNQIuPJurAieQXfI4J7aWcHIwMFRDdM1ZclYhN2wPmkpLAtT4e6gCqC+plu7G+
jHE5se0qg+NCVA0OZhLgPk4d55tP1eAASxselLYyZbnc/xaNheu/jbuJhais0rprvqtvo7Et2PhJ
8C0DF2f7/GwinfuCo06/8lGzO6FxAJ0dZWdYRyay+QlmwdCrDY+ttGQRcAKTbFxuf14tCTPzJmsp
zkeracpwdLPxjrGsDV/llTqtBSyIjmt55pSyibc2zAymUPP/LQ+wUWfs/Mqol87MuGwe/0g+/tAr
MLTGzAUW8XNsmd8XK/dZjOt9QUNOtMIyuPTYzc8MtqO/yb8/rwa6NDoFstHGxOiToWS11zHQej3m
ZZBev03N9LzkKuTnxuP5rRe3plnfCc4TeSBMkQwaP7bHQ4ty3Tml1AmeE0y126nxrAfK39LlFg/k
Afy3oUNTSF81n7LnCJ/95HqUgTRGA+dTOCdNzZcJmq4tbWG1gNAilYsQelC7k5DCwiG8hA6e+mpS
L9GEwwIr9l/hjQFLLgL/IssQkijQS/LkzFdjCxvUYYfCpx+z4S4npk3RyXclFIkivWuQPhQNgL4n
Ikz3Vui2OhHnu4SCRAxRA9KdAoWf0A1LzwL6GtTSedxw6BkgVaZEd4ggpw9r2A64xJl1sa1yFnhO
nBnSdxjXHJezpQonmD5TQB4bwqAaAcQOoajMIe1bxrivC0zGPXR+rAcohEahwXHiTx1tjrFeKivf
/Nf7GW/CcaoljevnTAoGt0dRPB8cvZZZ0RxAZop9FKneHCFEcEAsvQOLw7GIchIfxQwSNsFG4ox4
LKQTBd2Gq0ozrYPVXVcqH/jJyO8SOBaKLN+e8FKBBLy4su/3QVpZ46N+eFm/mciSjJY+9qnHfpor
qgaOJKDEXXUhsLGvQP7DlwiImK5PrfJ8aDo+2TPPAFU/ceYN4TbI4h0f8xy9FHAqCpv95zalk/5Y
kG+6w5Bex8IkWfVM81ieidAlW2sTw1fLvmuUwBK1D/LmRn53xx0dEl/1FWVKIpDLvsW+5SIPzeEK
6pgtCU1mK/nd/7NL6+ZqxNscRilguT2Y0JOgmRRFgbVEylRoBVybVgEDv2JJYzeP6/SZacLQIYgH
jpwLEbwIb/5f3/iocqhGDt8oTs2eL45sjiAGy3jgFpvLvA/n7iUmV7G5FeQv3cBJNuRVMCRehJOM
vsqJi4kJvcUolyn/sCJBfbsWWULqOI7QxKm5yjQdjwIAwmIR3IwF25ukPMDFy+tWpVoqjp5hTIca
qk6x/P8ci7+VJmBHdkkNmWGocgUgZmzg5/xlK+IbQA3ngcHs8x28w5Sz/hjiUXOUkXddUp4dkCYM
iXAbwevcAvx70xV6Cb7EpVWmgZmxJG2uM/b1xyY5+BksCDVwLJ27gIOyNYYhzVCqaCaap3ONTEnI
8Pjke340SoyPLOSiIcg6jR6auIQJD4MMrMQvvVj4SEHPNZKHJJXHCMtexVDy/KHkfbF32raAa2N5
vngRpIhrUvGfj7/smL/Tpsuu1+B6T7saTfNtm04H3hI+JDbfLtZJd7lHWo0rEqrHP0nNUJU5oWR0
pMuhobGmFaorEnJjofb1FwFTr3kB58E+H+zzOGtbgHg9WqsCuSXzVYSt5BOMx1O8IBelqXyyAUI+
PfJpvSL7+4XXkR66eYSPabwT6zktMC0k58AmXQHzMgMYnxrUqD0h5Mhg361N3NH/A70HjceeVNcZ
AFnzxn1e/NWBEojpZ/gMRhtq1kn2FXnRhcR4MoFUSKFBsWQXhL7gYQKNXM/3P6wSQpZnDT3v/rYW
IlV5Is50Q3BApcBRX9obPgJJFkyjhxugSq/7oDcxRo25gJCm3gFz1UoBwOE4krhwgCmohcpRd8q1
JgXp6yzAUV8jpmYOjbzERxUZbTvSBsUibUi3uXRht54+Uxed6D392h9ydZikVpYBUN1e6PmRedfd
8tHd5eH/3UvXUnFfMkV3Jw4oC4225CutB1TeNRrPv9JeRJh5EejPOYmOROTs888L6etosKQgLR3g
ThAOkHgw2l8oMxZPndBxWDhJDlrE6lXptmrw5H3HkX3gOkP6bVswSOg5HgEjbkBUKC3R99XVPJU9
YuncO+tn17OncYuG0iGtcEWlW7OhrFN5rFkrakEL3Hs1rzMGoUMIA9HJyDjQdi30KgbGRQyXYye0
qunfz7ied+vFVk64SF9uysn5iDnD//UShi8hG7wg9HmI9dhOvzQ+/sRAvkoQdRqEEpp+5XkdfwQP
NyLArU3Jd+mIeP2Pr2wzNah2IFawXko9VVyxqQbwP+UFPcxOwbwHChYptlvRoYxHGkYAF2Vgvtmr
bYq/KLM/69KtTZrxm0CiGpfKiEVnzPSXktRwE8mJHZY9t+pbQR7S2zgdIZ1d6IL5H0rHwZ3vw4/R
1JL3hnpWhCKVfi/Akks1CPODzXuVnnYhOxN3UACAQGQVHEVfDgAJa7Cx8r+l5mc471nVct5S+ehY
roEMmwz2jDFWJLYu3I9Oypds5nfGf+ey5bT/UcyPcfWo/lCRasFRpN5kVBehTcUSp7VIPtSm6NaA
R8LyKewzOz26WoVCidPGdcsH9aJ4so0qOnWwX8Ba+DesATAPzqU8EtFs/u9QThw8KkJZdsX0msdk
+RP+uBbhKsmwddQCgdkz1hJ2l0dsVyN3vH4gkxMRjppLkQsLDeLgA54Uhmdv9mz/VLL2aT2CKpze
R4BlosU2p2nzFbr67jL0dKfYvTPSi0lz9xld4jPvd7jL34BO1b3gaM+3JUWV6B+LpP/4OpG67Q+M
QeS2Vvcqxh5qCVYhprdAxNsZTswcwQ6myMzxuV+bcEjk81wE0l7PbPVn4ZMnMSpqcHmnRCAiCLcw
dZcIe9IUGSp2vrZJ1sBevedJjtnOsxZ+lqygka+BrmED29nVoklMeRSQRwC3qykYR9PvLuZj2Nsv
E3UI2OJ7lVqNrAdrPJUr+BcvhgLPTs3h0B8bCt+YdVjvCPNs6ZA/SRpbX8gRErLZi9bY5PNql0bV
ZICrXjxrObhIGyGYBM3UC0bCqrngNaofiyEjYjtsfPAf4SNBeVaSLHtw2fdNzRG0TDi9t5XeQ4NS
SGb5/OAoXfThnRl3aoTQX59p8MhXI4EsS7B89skWT0SGRq6qm7lyUVux/vTQG8Db0WOTwfQLbuzD
kK++na9I5o4ItAb8D73YwhrsF9gK2nXg4+BUpPIheS+FYoJxZrU6ZZxzh25OBQDznWY2zPCj7iAF
m/Mz52eM9YrXJR/BYQVudZWpk3b6/upFW+qa6cP0ltOHKXFj3SNQJYXKy67NFzaDpuo/7GanREvu
Kip8BPjBc2IFRWOM2KbxlEfEY4vGWeoWxg5nPyCrI44i6+RPheqcstdvilld9HkDT1as4BoMOqLu
yPOFy6HVej7fYZ2vk2gSQowFEqbTBKXb7m6zVo1QMfvb86UW7PProUQMwRNZEmfMwQXj0uuSgU1T
ErwHfCjmoj/3j5mI7cJNLRw9O8Yin4GqyR5/obtBpMZQibuAyN0JGbJRG9RV8XyqvKUIqT80OAVd
v1t2BI9YN39ttJ6hKDRq99Au3aVixXgj+HPjChIWuDPcJ1ysAxtoq6pTsZldtzYSMV8tXwrXKyXu
hn8Dt9gVPwNGWvEJFctPR4g+pbKctgeOitlMZhlJSn0rHAIlCa6LWLaKz6xGPBIgXlBb4P7XFBMj
dPSgvDQq3/cyKFF1HurA5Y+XNfJCAgwUFQhq+62NyrBiTtU77HupoVrakVQvOLa5Q0iXT9n6k2CY
KdzE3OJ1qJQWPoKNyl4y6l0Yb5sP4KGk6lMnlaVVbWfjxnkYCQ40bXxqklYWdZkCoC5Zri1AVfvf
MymjMCP1e2uhN3nRh3TDKUOdRimWvDzOJB8zUVr83g0/0b+QiXHFKNKHHWisizjQJt5jMAZX11IZ
Yi+lIsQ33cY8vs6LGkzRdx47T62PiyB7X6shT86dwZ6xaIg1aHkA5/+A6ByoXQEj4qAJFxFCVn6Q
UgIEpKK8ZWiRrAamGAMVM6lIEKEkxfO0RZvWS4PcdApbdlWWpa4d6fnnC00WBHt0Dtami0VtDyLj
9fDbGRu6MCONi9zTkap7cuxiHUh1Mj7yyw91LZC0+y7zEGJI4w7Hmjp5Otm2ksuL15sseYCnDB3L
jsEt0uFr8OAbt0EqGXdV2E72IY4DdpPj2fE9BZWzhjRGDOugFWx5h4sjXt6ffX/Bh3Ma0VzYCxD9
6/43UIWHAVPz0/gggYONlRnfDK99dV4qR7HTjvRe2c8sMOyIhdHIwc3P/LbLtT3FvVh5vwsA5OjU
n6AvSPHKeIi8222I4ZbEOLTSw6Ay2Dg33C0XkNSMGlUHlwu3aKef104dTZxpuYOYeVLVSKNbPNpZ
mYTu2bR2TYGMAlbLmxkDitKwPlT86a9ljBM4QfKs+OmyJOt70yeRneYRCdhf+0dknaLZC6bds6X0
UYz2Us9hu91ITNmZOH2nhlaCPRUDXNoHoJlZldUklPzyjpRhfX472V+24iyk7M4Zien/NPLaurBH
6hK9Y9X5e+1GFTDcUtJOeFS1FaAxjMcIy1/69IfuKZ+VvAmdv35V6Ef5RnZcrBgwNSNdsRPcF8RG
RN6xyBEGpKLEyQZ5ba3GFiTCPnZWyo4R2Cldec+zTifs2zzPLs68kqpHqipMWWQfv3DBJXqOh0Ua
nwuvmvxlW1tZVM638J84LElEtAt+1Kb9I4Vmg4NNyleXJEM+ZB+IGqxSen0PQdWT7nZLLvwIJ6a8
AKpAAwYQgJ79z2xGZye25N4IivyvdI9iuzwzJfzsPDOttz8u6qCl3G1WiREkbEk4VpWnyY0RhYNL
MC0wKfI7lK/mNhNGT5dhvQTmg51KNMGjOL869PdWJxnegcmBgZiQ8taXSFXLHPQT5X4W6CUauWga
ICXivhk3ZaMlpICM5nE7gDin+7q+xS+KNxOBfOA2lrqIyFH/BFZHgSL5aJv764Y545xCfLf/MOZs
dfMV4oUhtdHYeBjwj+P2Zji2NU9J/2n6ENiTM6WWB7augBasCgLTnVVvIoO3CfGDuFx1lRvCBq1p
BGJ+FYAz0To8BuwWx1Dj9m6IxVJntP9vLl4X/2gtwyPs74zcOTfffZ9VXBFLFbe/v82qkrizN6Mv
HEPw/CpFP1w68MBSwUCJHM41ccxV9QzKWl8/2rfjWr6GZ8TXCl0++v9gBHJoBr0Aeqr3eeEho3aR
UhCfPXMvDMpYG21Y/ARgI5QrsfXynz0qXf/lwbYRk5Uwj/NPJOLU6NbG/+vLMUPErv7ND63iJpi1
AXT5lL6W10qzfO9XedLNchHf/zZliv7tt9wrFrm2k830RH1DxiEY31okX7VtGpYUD9CFhUdNncib
a4Ab3TZW/AIJdb/hCRhQoLqpWkt83Ul0cbrLc+DeCcGij00z50BQ8XUBTj6cQgbIJi0tv0i/+MTW
vbZyGGoETnqgttOB+mdW12+NRvoACvwnQDJl0Ic1JKnD0lDigfzV+uNNDkJukBvFoml8AujCq/1Q
WNTWTbfiPS2mMjZ8tAzgKP2iRVmq14SIpor5l4gZwdC33VNTeESbZ3ZG8CQZYf7IfOHWadIqCaNb
oADKiKRAXsSzDkXkPcLJKUmvKdLOIJjIbQV4UYrDl/EXb3dZNxseKMHwQ5NBxakUYkZgIOoYURzV
MgFl+zH774manFdpbOHAd9Icgtemq94xRnFh9bLOlnRZZufLVKyipkPXKEAoTXNBqx6OxesJR0UP
zduzDGspU8+f4Soyvr1eNz0kwzm76J7Chhmet24bWlSkFfwvSd15LD7JeAuDUkSGz9eZiKLcPraO
X3NW+yVxxDlAgluYBbOpoycmq93+ou8ES7EShDIfaX+2Drdur5NQQlsYG70cspskVqpsTHxdtoYB
bh4LZdjYDzx/7ndCQdSShOMdYJnJHXowDTkWQhZ8WqidKFVUvG/OjJOaf5Azoss/j0xqSdH9TQN/
w7UyTGU1vY47aat6/LR6ggoO3vsbb+gBOYeMU/zmV429UHliDjW92dbiZA0DtkfYu7ff/EiS1xXL
8lXE5PUoPU2gwe8nSgDCd1pdeQIbmCB6yOdaOZtesmAQsVI80QnaLsfi83qAJIWJ2kiNR+oE8r6G
6CqCCW0ChDealiVE9u89YGrKxRbykoxyCJ+blwkJSb1qUoje5Uf7lgyXaTP4s8sN428bGvp6TDOZ
F/p4Nhw+R4h4mZ6MIg8C9Qj7JK+T3q5G+LTV5cXMseW0FTPiPdHp2b2QFKGEH5QaxXHcYxt35Dne
i5kufTht6PhJhZ+tcyOCqwdysmOFfMLNnJz4cKxVvA3XaL0f+F9TMFZsHqCof8rRBgXcKRFig5q7
TJwIsy0d0SUjDAfYa0mZf7xYjqoBVfOn2FhpR0Bzhkgx0BKRwDDxe6rIJzI0yEsmriAlRwI59BAy
Y7uHyOwVq1L90+MXqYt+dPgcwnCVeSRP458MjIa5OhMkkn63JpEcu1OYYPaxtYmXXUHB+RhaHQ04
K7cf6m80SxY3LGJr3m72pk5xi1GiYadKfRAV7s+c777kmNTDC7jFpS355JcpC+5eRmaWHXPY4IXS
EyP8qm4Q8eXfePzf8TmVpImiObCxaUwiVcE/tUezW2WriRCb74ysfSI4AEfan5GBL0A6F984FxHH
p/vGDU8MzF6998CWabntj9J6f5AnFTNa3vt0SVvsFC217MDmvRo2Xh8/j7HgTVdr3dchAj9QTy9A
aBq7PzSpXm/bcFwa1szyqDZ8Ut06bNxSS24Rbm7zZRK4xq6xT3FBU2r6ypIhhpNaVGpi6IwZuZEF
jLvcfvR6H/Y+ZU6FLuN8ZAxMEnuVbSNgghARGp6eG52wgMR02CsL2N+r35Nmt6sSMmUGQpLt2c+Q
B7wFvNaRS1VJ00lx9r3d6f/TXt/k2mMQbJu9bUZ78FsFEP/e8M9bXWGZGl9gVUXQkcsruKoUFkPP
O/U+T1SYojDD0DOde7W6xIU4k+CXDFfURdeIBDckR3QZr1sII0Om85Qdxc3ILkuMguJS+HXUNjun
zDlgn4ob9NGjdLk/cjCMoK0sTxsiTsQ5Nh/9Q/ogmL+NB32znQZmrmfeMVz5Ft81RgsfB4WNycaw
QD5UJmX9DNVRaEC2hiqio/sv6SdOIPuZ7RkG0EDq4VQBrwUTfh/Xwb/V8d37N9JH67tI87IsGCjS
pQbMW8zCunsoYP+y03YGXUx6LJoEpquLrjW/RVR8WjSWEPRJMyaYjqC9GAf+pdaed2l+/nfkg42I
FfQGrqBbcaelpPAEvenUq4OuF3VpLc0G1ilyv/e/jBMp1EOZJbjyV5dIj5EpBDWmAlR9MN0dZzKV
qji3GmdrQuuaHOnntax9kOHxf15u2kufUoOJ2jd37+fIDqoeL/DX3zFj30/sGOMwKZFu71Np3wMo
fqXFTIMHo0wBYlfLrKHeXo03LZb1IaA2cwnh7tKFuw0muYOf89iiUTK0ZiPgiMYx/aG4bBaZHO+A
Elna1gltAXzA1KcTKN4eehGnKcG0s0eMUGAxd1DOlwRvkWRQnDqsWy4YrFG5gQylIqKnI1SI/9BY
uYIicP9P0nPT0tpnP4QRww24ndvfYjEi3TuPlUcnVvhpx0TEVdzTLWfDnNDHg7+wQa+rDJR9P0Q9
DWAoLXN7fp3zmNylrYeR4TzP8uJa/YAYV2gmd3HEkOY90Mk7a1GY/yuz5hRyanf4X6Sgug5URJRE
stQHppd357/oNnUckSgQGZ9D1thcO+j3cCD+O28ZrwpvzGDv9eaw+3vQb/1bl2Ocy9UdmKQggjyu
Sie5Hba2KpBLBhL1127BqZhM2b8A79iG0YXX7ea2ZlHJz64hJNsrLsGRDaRn0KKrHq3xo6jzAZKS
Y2dvM7Sd1yktkekjy7GPKC7AQAiBbyEzQslaGE8/m7WuJbkQKKd0kKAxlF7VAWZ3ARch3W8pyWoa
BCQyeONR4itS5WxUXk0b5w6pIFj5rP9YUZHWzssA1nwXf4+OK4hsjG+JJCM6lGCLB7w/ChappJLq
7VqAm+9cLkTflyyDRIsfJkd0GIeCCb6G7W4bq9EDLZRWWUGp21AUL+tTCNuIbVDUxnjhPOVEDKn2
QtvUyiEMbTWMfkmbRz0wlwb/+r0X4KDSyfFAjqig9AUFlvHm7HFn3uea8B3d5dnWyrS5cYoeerDj
GrmV8dM3P2koB/oIPBPZZaxBom2/Z1qW3lwGK7VdBMhUKsyXXHKuVyM3rchCBSXt7YrBaruC41Pm
IWHc8wLKt+/8BlC+bwCk7kkuvo1Ow59iMhiroKH5HRz9Tw+eT4QJPzLN+W6qFmLpG5Ar59pfcPNs
m6VBIHpuum/u2+P+WtgQXmCnSiArNXBrhpbuZ7X0n7MP77Vd61QRVyQtdRr9IV8csQ6r6aX0vY2D
mS2suhsAPgWYaVIqXw88JMTUZzMeSr+ISZhQZSOw7f7cEKu942G2yTwLRvScrfIz5VDaa/6QZWnx
TTYHTDFNpUi1Z62ac7JZLux+nf5kxWsPg4aceGDGnci0O8kGYvB0LQ2XV8p7xdvzMKdlJvD9AI9w
/Qeu/5OW6ZGDzNrnlcApA7s0jn0uEE3PrabDqh7ZEXq0LI2MiFIHo+JfbjJa5J9bkilKUGcRR1U8
UGm+lztW3uWzg7nMpmfADN3HdyfrgBISXIIlrm+KrgGLLLYMEmkmC5vlT6USqFVggT+TMsTsUToH
V1hoBETA0/t54HJitHwjU1x79TbWiusrQxImviXCdc5O2H1F4eIioW9dLIQWkAi7ayFuj4x/ufzz
SkfxddPZMKF5L9juAQ5auGuCR1DmMUCxkednbQMVMRDBaCoiJxUKfkWrNrVxLOBY5K2NlZ3VymIv
T3tgMox0pnpnVNEg/HVG5WsycLpmYLN32F5EnLG404nWKGf5bactMDERp4roxMgGwPW8iCVHfloF
9fz0/uSQH1G6MBM92uzw0vkrjxmGpJG3vHoDYO8lgm0foFm32LUi7bFlbNMkHRi/JQ9McvlKWaup
2ulYfqymE49Z0NNEJXffG4jcVVO2P/8rf66Ag9mPkZ6YXgQOwreFBQw9EpHMQAAs4TEE+p5MJ/h5
zONA648qpfkl/4lxnWe0VM4Dy6mpX8EVZW7EURTN34bPUNcYU89O8Spld1wa12s00COVaBnnpq/1
2ZCU3OYKMHx2QijO15QHmrao1rYnLJ7vVAV+9F5MtkbqfQgdEO8xQC5f8sa9wv7O5FPwF29GZ39y
rf9JWjB8ulxrpOJm+2CVZ52vh1LyeH0plVtRIXYS4s+2NiEAXLaEX3jLQogdw233UEOfT8OMUrFp
cWqpzIdZWbfx7l3Ca524lzlwyh0Ex9o+xm0lQG0WWF71bw9KsTKwhx8gkQkJ1JTFrxAm9lFQZMDe
lV32VEIhWvtxIBDLjDIbDYvpSozXtEVI/Q71cjQRxHnPpSZ54LYsva0TzXN3rGmSy+9lS7SYChQU
/K/JAf4o4zudeL2jtSTQlKhim3mdD47xmE7lvXXJicipl7o9JRGxQH0N/l9ZlpWEusO9h+zdeWFN
ZTmiPn9QPsk2YIZJhWcuex4clDOwdm+8hsgIhMeGxQouz+AdRetmjWB53zOjMZ1XKm+pfLG2sdph
ueIkg34KsDTZjQ2sgzyRkhEJS8co3CzrDR6DyGust67SIHhZUyDWmZS8wCyFcL2XFQtvM8Z4nG41
KiAVozT/qAnsKmgCj2wYw9i5MrF2v0q4x5Gee2UrE/qeO4lwPLSXKqXX2NLaA9gYa6Jt/PrfyBE/
1oAUmWctf2LCs5PuM/CEZiUFsLhw+XTYP1N0LjmBT/U9YYXg+OBygb5gcG1X5mcTdBXVFo59MN5t
Odf/8snXDn0neFnJGcwdR5sWdnxQhzgWtLWRLLLrSRMiglCtHybSezdCbzfIzqTSflncNyv2yhLk
9p8EsbrO56FCvOLZm9O24QSeCUqAG+z39nSNm+e98S83TphkN4dBsKwIvLuKXY6ceKQqFEJmjMQ9
YtvCcKnfkRvMDQC4UZ5iao/ymanI2Xo4/X6EjFb1WT3Z5UxCZv9wUXyFhA7Ux4ezMpSs5ozG11ZS
Rz+bZpaxu2Uvqgk2hCQWXUVy+S6uBeYGD/uGtcAzSWVqOUgcIQMO+hOrcyerzQNLOfWEZzP+HAve
SREi8Hi66Y2yLchOzqWZTT1Tojyz1MqTrBrQGya53tKZ//iCyOptCXx60v6SI+Kqey80FXfoU7IA
KedUsVWbUHpyPTIhDJALNic8biJTrpBJxV8X2IBWeaUQgtWyf3BOLxbmkEfP0vr7T+fxjpdHF054
sMRwAa3vF/Ss4JLpJHealFcmBlcI1wUxnGQhCci4s6KtUbSYXEbc6m6hxQEy5yF3qmE9DhCWp9Vw
Y4SONac6raqN8elL71ND/NjD+ihpBTfX0pw82gx6bs+r0lRtZXuZ13F0/BUddR3Us906TSo5QjlQ
JPKXKovIh4wMr0SCSdjHm6VsNUIxKv34MNaERHlSPz70AEnHLiltSniL32C4iKWzV0kuxrXAesup
Y49nvDV8gQHjAgwCZECyW/dM0PCexx1MtgJNdzTdCtUHR8KJamY0dMKL7fxS2Cs/YIbWS51I73Ek
Y8FvFHLLsv4YU5cc3Drk7OnqyrivayYXrylKn968TfEsjYC3+RifMcVw+tJCx0foRJWeGyMQvJg9
b1O8Elm6tspMbS1irRBGZhJJDnqfgJZhQ48QgbcXxOKy2mPlLfqAxrDjXseWsuDkSnkH0ngJ4S61
JP2anJzzzh+ThQWeFP6BhSlo6rBxVnJ+Nr8a/5VCJVioQxryy7FWIdpustrBEudtutLvflEimW0C
wGYOnJ5yKaJU3FZMDiRUZlxm1eNibFMFyXgf767acpVMW1VmpVncrY0gr79ZNRuuMbwf2OZW9ekV
LtckjxDnCOkj2aB5FLW3IhLx3fV0Oj1TuIjrRWee3WQPIeaRdrfDVKVMYJYpZX05yNRIiLW2Lw3I
vyNLh9l1xxfwfiM5h8Ly4cqfIQVYTWCR8dJVBMtlgPdNemNhKi0qexRr0YFLWcUaz8pE45Jd3eVY
PQtmkQ8UQOUDn1+DMO163y1sqoP7yhU7QRV6M4xqP7vGvrblBXtHX8vzQXN3Sd2vdSxbz8/Lq1gk
URaaYe2pJ3kCPwjmPyxC4enni4Ma5Htj55u20J68JD0LpATIYCYWNaGchObzo1eej7mTc5zxnyxJ
M7EsBjISPfF5roFIDvU67jTsIWgX2sUYbXYyBhdwkcYpGlZ80QvoRIabV/Vdhr1+h5l50kOXP4UV
ETfTBKS6mnd25TQQrTc5GyMRJg10cCfJNjyp58V5w4CXIPn5GpAKt5pNK1Kn78JkUdDox1Z9KJl1
QUNTv4K3LIqWARgGMoOnovtjpq9whQ9VQBaKMf7M98FQuC5fNW3zGOyWLyAvJDVM2OxSYDJW9/SF
dOSdUeeEPfBI1CIo25cSdXOXu0sh+P2rBvz59TT8QMg0oBAVamGEtfCYLe/1qFgKHuthvx62TsCa
clyI6MIMkTwcheGYmYWnpvpGp5XbVMGprjnfbeTVTGacXVpBY7nTQeotcK4XZybOLOJUHKNVacbz
kNa+yxGg4oH3e+mvGssBnXQ8hF/SyR3XFeGwNO7l3tsWSlPhXSVSi+Ts1INiE4hlUmK8YcqI0slJ
RTFQy/EyYMuJru419DxXbqHR8OwWKl6ptUnhY/693qU0nzew6KT8+7eJw1KfpyBOTPlmkaU+hh3E
MZMRzQwT44BtEO2b/Qzwxr86EcotkhwrnIdkGotxSdhQAIyf1Q3qoZiyz3UncFpFO64eYU5AhPw5
d94+ueLMGqCYSXGITtoqniX0wmm7YlgIoIRxIQWL6cTvTnmMM+aGbmPgbEYoYQUV7e8jeRQc3PQJ
fG89W58wSocNXQ80b/udM1Kpdp5m2zTqKtQCHLIKSFGBVt2tisQJ4+RUo5BG4TUTnjiHckDuAjW6
mFnPZ25fNnk6xOF9DorQ9ED0ayNcqXr6LCWFyBxdcNFP3U6Z4W8oXW+YE4ixi/LWs4DGdFgWn2m7
eOBarDA4hfyXfEQCJ4LabUEKqSFI2jn113OM1QjfI8cfIYj9P7i2yAslySJJW+Ms4kYFfhSX95NU
vsvxntCzv9rEG2+cgk5du5fvbx5iMKbT1u0fm1Qn7c4/slbarJsP+w4wgkfEGRvO0/1IMLu1fdVs
reTp3GYSY8uT7XZ0WgP3zhqcomHx8Ndtb7taM/k2oqQH2M29fZYnPqg2u3iB1/642OzrgZhAgb9O
LPotlm1ObZoda7eVU2JlT+8E3Y+5Zr5TOHp90loYfAf04uC0hHs40cHkd2ZM5/ZGIpT+2yWju3nZ
cWnVRmBjNjkc2VQT9nq/nFpQ2Zn/3GJQZYvPoORL7qaO+zBRgLMaa3nsWqQgojaLK1d+E8tcc0VB
ua61jvHHY9DC2OBGuvmZvhtApkGtC9PDZRv1pLXf730wWcyJ/9lPeAkIDBTFZb044WskGc5syt43
wzJctbQgUCWA+jWJCu/X/oHrjBLox4bRy4eL6ImjHFxew1e5WAUGMI5gb2uPD5wke1FaJwB1hAxX
dfPtJQvMyC+tkpaXGYdTC6P3FEKv82l89Kyn07jm1Z1uBOTu7G1ysmXstOjNvnV1TXAOohEetaOX
jjmPw79wAy/UhpxJp+WJVtR2MPrzjELsgrD5JQsokSoRyO7U0QR05zKztgXQNGPaOm167RAa9shs
7s3oy8TECtM935Hh8C3rI82Y7ard/6HeC2n30ZLyUd4SqH0KuDndeZvfu1Y9FHzWlG4nCDo8G5hN
X+HNu9S2E+0NLcQu/gT0s9DHaH1YwYLZ6kdFr7qCpdb3+mABbjYfD+jdrLfZrXSH1KTY/vhyQrOh
uNKJu+mIPON/kxkAok2ala5BBlB74im09tO88Em/RLoY66XkR2AhQcaIRuYp6uB1wIKWc34qekdI
KO29ln6GBQqx5DOqR2mgKw/xFdmJ3yFRwpjq4P+U940LO1oysrwQ/waeeQ/23JC4eEWy38DIJ/LG
8U8DM80B7WWLr8waADqAwQG0ChfXxSC++5puNiEg86FzgkTs4YWhlRRoHZaNAbB4sfFApE7++Tip
3qMpWa+zhtNEsqN8fNRU9iiSSv/KNMINvRef/reAyJTcm8Vqb3vEVz/fkKGb7PnfWokpGxFiXyqH
UYBwo8mZ/IOYzXTZyoKi2x4kVQrLYsMyYhfpGE4rk7S2JJSjJKQr7Y5Sl/NbJX3mkNvv3xB+PjpU
sgWih4vI+J2YG03zCJHt9dT7UWZZwBhvlWbe4pJYgAIP6gjHXLfBJZus50qa7ii0f/iDpRiTCkIs
G1Y7Mxdbge94qmEaIQTA6LLWVG2Ew37akyLa9xT8ooNzBgFLC6B7uWkL0OeQPtA55FwXy8SeJSAf
LSTnp3NoQtgrJAD4TfTqrTXyrTaemv4qkHT3VlYZLBMU+h8duWQ4C/PdjmACoqTKkRpKmdDkgE82
XaVuTY3SJTrWPq1gRWHCVcQvv783ycTsV14sUUwZr61zqJDwasBV4kWiE12eBzyOkHLfgTVskcnz
yjnN0mmAqge09eM6IJuPYu1GImToaXGXx6HQtoGxzzTaaxRSUVpUDkaY5qEvGHGkxtxFPYhg4H8z
Z+1qE1sh6VXxgK4z3YNcGbzCPFBhLaZPsroCXPNPOmVfutNxrub8HBmro2mmw07NDPtkregAEtum
toT9ZO3o2Xfokvi46pbRiPYwumUhqnVwwnkEWQazVc1rLiFW/pNFEncFXmdWZK9AXDDG7opwM77S
YzmA6CUvNp2G7XR5F7pYq5DWS8ihqwp1WtscVf1nQpx6StX6unkbRy3hj6Wwo0sOQkDkUbDIEOrr
JFENp3+iDSctB2t4bOQoNdfAa3YNNSOdYUZPMlRPxYdVfysGnQ/y0iGuMxmZDk5oqZfzwKFYto5F
/UbuclKjryGHJlugvjEom+U4TKma9YQ2IaMR4XvM031MyJCko2iNmXfAQnqfWkZvvNf6hGxStpwW
8tHXdq9X6SoqKrur0oE0b2GAOmu7fiDUrR/ZFLBPC0+v2YrkTHnnuC7NwZR9AhFn0RJYVrNzWkQX
vDMp7ZU+x8LDoD4g8uL5iSVtpFnCIe/zO6S8haVwH2RunANbcK4KwbpvUvp10CqtcTuuT3jvDrrd
Nep20rzOF1jy/CngRGcPOmtzv9XkvsEFRnbnpNUpZBX1nqkOgh4Tnm9koJcSsS9lgKfLvC1kffa4
LO7FyI9DWtBWzszJpw6QXjiqcxKQBaz9jl0Bk7aOYaLXAr0q3aMywttEmuZmZaH+L4heSjeFYEKO
fTuqbbeK/qjUCjyP1Rzwr5FzZwltAbO7i7gj9WHCRedgb3nYlfFvH+Qzk4C9xM7L+ONmZ68MyCI+
WgDusqzIXM3BNYEww9neVsiKorWNoB5DMsla80haI++JtkG2yLSPbYHAma7R17reIZkuWWp0Yv6w
21izQiIWkDZvA0fZYqQlzErNNi5T68xaSmehUXYC57x6lm1c3OKTqpxdjGkFwLG0Qx52RpFPY0uq
iumGFloVuCztfKX2FajWl3+1iQbzKDW7/wJw5KimDrdWuZIBwSFnCMtp57oY7joUuzBS1S3f1RTP
U7P21g4+izjmvhrkXWRh+dChDAMvmW7fCLB1ah/C/t7z4letY8/pRuwSCe+HHyVozOxy/O4wB8Ku
Brfvy8e/8ivJX/j7lwkk+fe8x6mFjFX0gM/1CgI3GWcxklKjQ5XvSwXnvXf70+tTXhv7CsEWULce
9H7BuwDjjvgeoqrKjAstkO0kc3wQEGxTnP75uCi08RCGKu7QywH13A8l9VzoJN0jrqy5EL0KEXzU
9L+UKIhnZ5mI2PGq8CakXAfOPij8ZB3AR9mO64/qIpPIwHK+G2mEjZ/sgsjQgNZtknolc6cFYZjm
SZNxZSMCp/v3eh4ZIHwObDGRMtgP9lvfl20CdAI+uaiTjfqTB4Po+b3ZZoD1f5WIT7xbw4569JQH
ENTNUA/OE+CkxkjL3aUBStojYQ0hE0zQFUGtqGhLL5jbpsiVTWk/2WlRJOtKcU2mxKiKmhBIL4dZ
V4EUH9asTXWEl53mZCqg6j53yMAE5yrhTa5X0HZajeniFSBzoy3sMpA/aUczlygDkkqvSMLUDARH
ujDCatRiCRtONF7TPg7alOXZRhvEmFe5SBuUuH3Ped79ENep6smaowou201xTWN8ceLNijqzF8cQ
468fnw+ATIN+4sGx/iugar4srEJ0X2mH7wh8/LoAyOFnagLZXV0oUjDeIYc+Fm47BB7AkchD9Njy
D3OnmZuGdWmpFXGqSpX2PODUmONtaB3aD9oglFm0FLS6+AZZjZdY0iARSXDpdsSN4CWk61i0ChDf
SN6VIPeUlKu4ppgKisVmJOt2+MjaZ9Uj9C/XRwg4nEIoZnNerEQK0+PjOgTXce4HtldBDv4/0oOg
ETlFBY7xdvkd/cNMqeks+67/XbudEiXTuwSXDk5LcADTDyA4EBKZeIGjmW/ig3jD/OZsN8x6XXkE
uvFmXASszJrfZoe7qMZf6YxkH+fj0K6tgvh5BQY6d5WcKe2SHPloHBDUKLE8az4muEl5XmvX0Bzb
2dsWSe0JU5a0+kyOx7vw19XLWApfURhFzQlCe1GErzLh3UyPGGc087hKBod3e6jmaRXNgp7IjoOD
k4X7gf04qQzOLO+tSOAUD5vHogcWfIZyRyZaWCNnsEIN7pGSq6KZR5pzs0lxl8Bzvt+0aRQPEnhk
tTcjxR2+TNYIgusD1B/WI89OYySb96enZ/RXPiKiOt9QUzbd/mq7HPocClxVf8e8KTwyMi1VpDY0
GXt/PCJfu9QIsHDXHKfx90izxOcBDxv4O2KGN03pwb3LVtLnUh92w0kXbWYf/pCoB+C+wNPzb4us
/fX+zxlC6ucoJ8EVDFeReln+n4r1unfqzSSyGUv7eg8IbIXRPxTnrQx7+OIcZqdOAZTvFss3eFNC
hswzY4PsPLZJUOGD//6BKCxuIgCjj9tX8rIAUJbguZWzATfQvqFEHcrtPS07wj5p5nqV0vXmxAcs
8JRoFvgx0cHFgAij/qxyN463Ylcpj/gy1kGxZOaI9QSkJ3GZC4VbL3iDYXrZKGjOuyc7G4bTIh5L
wfsuILtRnSTo2iGLk3P8W47GIJpEp/GijzZGwIU3IAlhdPM6K0jYf9eUij/Du2Gg2BT5pD1d/PyN
NBq1Kre/9xrpuuYGf85MuGAt48GTQ7xksqNJDpHPFmNYCmpQ7wIiLz/2Y/gMOTXoSPimHaPnMLcr
9lwZi9se7xbX8y49Gh9ugSI9Kgoeq1PHGpcST1BP/ZvEsSXibahPKQibT0nq03xPExGzwx3dL/de
QE4Zd1HoYwFxM/YURjl6cd6IaBxRFjLZTfMIfP+ZjUm2pufzutrQ/C556D0fN2KObrhfQYAzAugN
QmafmMPV2MLjAeSj0ZWS9Cym6LWyXpaJl1tBMys8yyaRGibB1wucAWI0qYxytM3N48ymmgyxDanN
0zvfITYKfnxukFvLEUUU7ELNOSWqOxZoAqdcSEZ8gk++qPH2Dj9yUBZhyWXNugLM+GQTdL1Cg3RF
2uljPnByEqaJy6sLU+Vc5ahNy/ZLCV4WgRmofRkWblkJ15L4qjTJeHrovZq7IbTOkksFntP43QKj
oyRxrRH130VclROH9K4fEPfPS7eKaBzeXwNh4kDVdHPzZmkErkPcubs7W1eHgYJb7ro0ouXG2kaN
VM6ERq47dspKXNznKX7cl7sHhoBjrVeZXb4Ad6Jm8XI/cTiHPvzL8Su0g8ck1uiipB4JaP8XmR7J
MoShyo9GuuqSWFTA7Do5OR2lI2/l70s38ijnOq/nnP2aFg2/CmnYkrb9fAJxLZ7mn1bHHLt3GCCt
Z/R1W5IUzOFtUh+KNp6hYrQSFaIqwK466uE6+SZo8oDog/DtEgT1GWBz5H74ggX8lr7hQgnlFxzb
qHCVImsIjL/X2acX51IY5nJHDsupZGKeH5gC79j9DfiJhA1OraV4RLgheqG0C6QbC7vvnBaYnuWf
Hx4gUR17DhJGKwSX1qwDfjSVQZ7RUz7mRT16piVSclj/qHjydlrRe1/e9YjMcMM0y94hoNLYZvGP
0x5W3B++xlih4NmeUoK2tLf0X8zbDcjpUll1dK6Z9Z+SVLTp8B4eeEzcIljbuAqaT42qq8njhsAG
Q+s0B+yIQXp63+0CRWhtHs6sFoBEVzibHHniaq6FoautSYv3G5zJEX7A+i1+IBruvamxmqr6TZ9Y
58f4l7hMGMvLot9JTSl8Lj/4kZUD3Qza0PCmyzJaFZEaC85xaCIWozu4r/tyx4bBB4wwhV+pymhw
Suy6Ue+8UGCeBHlRvGlH1ieJReNr+vod9GnSepsWIS/efuaJ46SHnk7DP2+zB03yWbLVnNroNi0K
upOnHtKX6nWrkzIncoo6itpEuueMWtj8Z/s02eYn6FLPXWqiWs+NPFdvNlSKKiwxUE2+9LK9q369
9FZcF8bgzbgtTTPYRIHEH5Yc81qXtZoHl3ROBJM/Kgb5/6GlHKlFXpUitpY2UCxXnwmMdcbDOE6v
YvWg2nTrXfQpbWJC5LpMnTS7EwxIjAwZo+nf1L75L5XahbSVy1rOGys47B8DuxHxUF/qCTSgo+Q0
C6pH4asOCxSUN/ZXDVektnEm7Q9hbdHjR67CmYjnRWrZ4bWAJ/VMfFwczDAOX7x5AR49YFTDl4x9
jbv/VQ+ddGEFu/pvGsKcteP3Tu+06+7WXkOOuLOK4LyfsQlERHgL+u04OtxCDfYjimc0/RDvicW1
c+A0lluGvA5NZJ00s6KanxIbSRYrwnSUEkRF7ap/gBTrmuEDCwuKAZUmhl9X/jMBx7QprOPNf7DG
TXzKDnPnhOy7vkQtfTmI+gHkAel9a7GgXuuRbDFf+mO9sfO70gguXUohF3SUlz0p7jmDchltAmwR
7X/Q4SgH/r4qy7A8t7lu263A68gJS1JaRbh30N61fF2QowdHXTtDnC1T3LsJxt6kk2oygIPtl2Sk
bmOkv6Anh1XaheftnLbhsaiOvE2y7okksgbEEpTJLp98aEXDrXR2tvU/k9ZGxxGzUiygZ2Tgci3h
dje4FGtZwDPfK9s5xy1xlJUUCd9yLhl7cLqx5yLEl6pX0fWnB7ddx2bYBkE/aZ182mHJpUj419+o
OEEyqvqKCf9rfD1dXjyWbrcLRngCrz54km7XSOpSN45F89a/2arnOwZOfAqmfPFDtuhTtZrDFk15
g5vwrBcrLUg0005Kf/to9lTqj7rZlWEB0FvlioEKLIdUxS5vaQ+doDXiFvbm3uWOS3vfYUSjUisK
0b2pl6H06K3iZEKATbLhgODDvJhjk3VcXGWSd8bqOe2VrAdI8Tt4LX9znePDAbNgZjal3W/HMm0A
OV9Q+hFSsHjtxtbcnyVvYPKI5MwohPbQtetzwxgPe4NjdWMOSfHaF+gUEXkxRc0memDziwto0el/
EqYWtRTf3aauWF8eglhXHduTrS8hzV3+E/7NB0LVdF5g3uvTE5t1cwe+LR/winREr3ZLtFpQeSsD
l4rP9cBtQA0Qby/n1jW5UXWdRPSOMdWG0BO8MZ6lYSHN9QUbYsIXPGyOcUEi+1exeDXDvQBaUF/9
Uht2MCnqixS63SYVosdURTLEMmrOdKElM700MmmxooZkkSdr7EdJJyAlEASGD+pKzgprvhlDYpTf
Yhosxxklf21IxlzqSD/+09dS+N1q7pjFSaYlxcidLr9kqq1a2MGXGziwRlM37GmY6JPcMkT20Vn7
tcZ80Nad0SRO6Bs4gsRzSWTM8/QMJmrxM36TLZmph7nfiQwoSZd5e7nVBuiTdxFkQV62zVCqD/mW
JH0fYCAH/Yx0iuz6wtW6VwYqDtZTnW5BYL2a3MgX0z8VXL95/GvrJhMw7BlsKp6iWybCBDZCkGQP
5G6LgTGL4iUbDF+5MJiowJ0hnGlZwYB1Y5eTzVG7rSumgRsywwS6CCEmgOgcOCtHefFGE7SSkjgs
5JiSCU2uvD7HM4IS/gadk5nP2iQySm3w955DUUbrT067ZcE+1RcDrHBRsgmm1i5w51DDL+BU6XQv
T1zzlP1YbfooK/CMsm4Uu4IkYwcQ9cO50Df5kwFnjWjv+iUGckKQyNlByjrV3ObsRitpWTn9XIiB
zGo+imd6tpynpCfziiRnTwZ1t7qaeLpPe3bk85W30l6zZreca77G4mRJvuI/2v+ByJPduRAHFC57
XQy0rlm0LtkTj4QqaxjNrLJKnOomQBJyJUfZ3SPJ8KYr8tUpmpYKNrN/6DgkpdKo2e5rKW8EWn19
9Ib+ZJDdIHpCXvjeVC9+pZhiAUCE1ck/4mJrevcZUkdp8jUoK6ivOL5JVjiA4HGzNA44yZ+j43T2
fMZqbD33qLO4EQ+IvCV8WoPbLAP5TETgk3Yxi83WbBdE7b0zRUg1M+FY//sZaaJEmCBv3yqsfYVl
mdaOylLyISVJx0zDkX0gmCOo53HiPFkcK0tYR2aOr3GuOQda92T7f68NSvooiEOflVY3RfiMzARk
2Oh84UHqhrX/hUPGRJwfIK+vNLCt+U3fwuAq03mUyIrJD/koCr/wNwxhKf8fFBwGn5dyaPW0rGKD
Lu4J08R6ww6yivWSRvO+n5lyzRiE+cwaVL55L8+dXdQoq/HLDF8yfYF1h658YAyErfUYZYIAzNX+
ZVqh3syrS96EEvVu+NoQgI7tIjiVZv4RLmsm4IETisVHzoptFRPlkoMkQpmEkCneV7L91I05bmJL
BUjyLHhKgMqZlgIovJzsZPqJ60q4hyyt85EEZy6HaqrHP32bZhppGuMctCZEpWB7QkCOOv29xkcl
yl3fJEJpaZkFn52c7cPn2lL4N7hUaIBkkoqc0tlPi0USfY6cwmWEKIUBdNU9sLV59sXDFzGHd2Wx
kwgYYrYvObVIMpsBNp3FSKIYlnTqCeZwnJoub2BpQw+/+QapamZjlaJXlm3Szptp2pQPih01P43J
EsDEiw9wNMwQYGsWwVxSPfOz8lojxkrrF8LSwWFZrjk8DTIZXfX5Zx0BBbYNp7jkRPXlCwdNXFl5
+sK5y2iQ7Wni4Tw/3GGCDF/50DVyn9F+lbet0GzSuqVDMc0ircSWFjINQtRIOvVTNE7wrc1AbXZs
j6l47PyDKmKb5WHWdWlK9MS19/+V/ciwl48Art+IBxiZSQVDPqDTz4bRaacvHmu6QId98W3RNg9R
YPHsO3WCDKZXgodIQs7GFxEp+83eoBGg+UDfap9cWRJjRikWz6x4XJHj9i6pa4/r6JagTSJTeP4Q
zECCbvv1ObXadP17E39QjCRLrOBJ70h4ZRwvaQsugJo6cEHTOylZsjHjbufk474brjh/J+Wu6u7W
KEtTdE7atTWH4S29Jmh70NVswYyB1EQhqTONSx0ar7wNminO9L8NrJ6nijdBMTidbwy7ikQnztq6
HDCDwXA/azZ38vM2P9bVBOxvRteFQokwVTskmiyJpiU9nfGJYLRZsTg7E/jHS/H/DdUtAjLRa1mU
DAIJyzaBCBW6TulilacgVk5U1PXdtasuXR6LlUTOyMnazuS3kSKufH3iPTq7JrYnFJivqnJJK15r
WpnCpzHNqmW2Yj/CncslfhNbPaLlcliD9gvWVmHS/rK1J4gUE1nf/jBIveqCny+W8I7hqlN4t6ey
d92T8PlveLstY6cqkk1d0bkW5Lao4k8ySi8rus8MkkPrRhtNFy9x64h5cSfKyx3YUydzvrIUTAdC
2WHJ0ZwFfDpd1NU8ykIFfF2b3vlsGkuqUrSAXTbnYMODWdXatpTJM8mQu/9QQVaSkNFmpzoU0Nnh
oaY+E9dfaSs9cTCRZ3aYosnthDnIUgXHsYfSAaCeUBYENS8/WF/UHIiMbxVSQXa/wyVztM2kiKT9
IHhyrSnJ1Hj9gvYFHb6F1/3sFk2h6Ctyb54fJCGlauGyKGIQcG/1NqVJamLWJS0r0i6wVV6qRHFf
TKBcnEPhdsVLbbRGK79zghVwUNhuqBGzvsQEjK0qjNEhKZXTLE736vNbdXooO+d/mGfNTujpQSSa
ShHEq5SQo9ljEbgdvNt+luBcAIz2I7711Ut+YtXOf3jDArTSQfRdrDPm9RkNVe+vB/cjlv2iG+A+
8QqFYrdukUl9Zeq1Voz0kFc3BIOxhsb9Pbp9KKpEEghUpWMVisQNSwflif2OsLPCmajeqFDuZQRW
jOjWJZRIr3LsisEdau19ZRadRkmppJ7Z7xndJ9jfmYbs6ZW9tVZw8PMTie8EXkxDmQPQ4kps6KZH
Dw5on5Qs6q3PpHyH3vWU2FvQtaYkB1KeOocgI5rwZ7rTdymQTwrlemRYTnMaWBAV+oqoAQS95RV1
qK0qNOBgBmEsi3S37urfRGZBjKUjTGHNJEycs608oPs8RmqwXwOYrfRiS6iA12qYOS16vNRQy0Ep
VaJpPEmGXZiz1n7MPrnEFL+1rQTsR1fwi+dNkZGOMaTZJHMLYMbDLXLwa1ntB1kARdLsGSWo1+Kw
2WzLdgpBp0QEAs98AHJXgQC5qVG3g/03VIt7kcJyBsIh7FqRHyDptYD7//KYe2ixu53QlHQDPK1n
fJ76q/wZJaHHo3vy2OSg5LiO4fT3WcU27/Ha1jsqdhpXZdvo409/mrqrtv93eLiAuZrJMlY9yCnN
0fhf2pc18AndZbFM8M4F7L2YVBdkYnGx3PY9YtAFoF+OMxFry/tdrqabhG+Y9l8AbgmJwrsc/Uyg
OA5Et8ObH3dlLBYelvqmWYQcuZp7UoHOOKbzSv5ZO5jFRACPAUi7l0c2JNVHCMpPlhHG4rMifiiP
t8KkNbBghGorSEaxYWdwZE+NXARpOU9NzDCt2I93ZkEijPcGhl67PW3Y7icMStxSTUE52mSjCG3I
K5ISbnZkbUi3hFU8w3hngWYCEPxTxiX6rBjAV1v5Rg8VQLF6ZIxRevSdxhdchGUu89ySNOhs9kHo
sb+1VzHfNrdrhbkRAa7hTVnS/6yxVQ0wU9RzatMnq2SGAIHm5LKWxk64QVF4C0Az3RtHm9w8ajX1
bH1jgTjEssQT11snhoBhdu9HVWn1KVoEtUpqIv9VI1FY1SkkCpAgnMchUlNaBluwEHvobCt3iXeA
2q90s6DINiCqgaXcM5b9OBmjGM7dmlG3kjh0mmz/PgKGwzIAlcekixIGMdrr/SDKx0niAEgNvuB0
VU0ZtFvzU8YWstIuhPxWs5u7RAWewnjdI2CqlThsPCF18h0cCPfknikEIddXijPFBldKxwswrh+U
bz5Muwg03Bx4CiM2jfrnF3qcgvY8ZSof2Sxr2ku4XS6Lg0M/cpuAcKz0+15a5n3hG1OjLs8xSmTh
NclgpgD7DMlJrA6zb3Q7wvUv4kzMqvswBj+YsQKmhSZCUbl5umUm/UnvhuUjGL5X6ySuzzlULhME
VKvN+nzgTq1xNOvzv80sEN9KYH4bCh1dxULaQ8k4Q1uZ48FcJsgXH5U73YNPwzmxTth38eFb5kFz
JsxtgyG3yxtBvHoms2xJ1wWXv8fYPyNVPocUpLtPvxha4vTou7qYyOvUiYlNOuSXJiPWcTATENq2
h23sYCQxih9MgIhch8z+oTtouP6cl2u8Mrrl0aUualnjpolSaTQHsFCqfTlojmoCtsP7dZP/apke
WPOYEPAwvntCQAh4eSPNOYBWZXHJBh/UhMEpRZcnzFCFOj6BxpscHSFE7Xcjdc1Gnf6WjztmtYUg
epW+BodhtLEopMaJEBf98/pusjeUVepWEXE2Mi0mHos64R4QdG2tRa2iC9I2fwgmfn10GRsVNXNt
jIW1g2pdF8tfeBp0z3heeyIGo6gCxNc2V0puolxnLq0lmr/uUW7StTkHJ+C/h9rzlTQK2MFqKovX
bBUUIQkeEVa8SQkNl69u+RyUuWAH5BbWM7saPvjSXhLjwk4LGCOZLFKWD/can+dCgNP6kBCdHW/w
AB9x+g5B2DTI6lzcLY3uti9QsD1rP4ziiXQ/5fMIoIyMhQ7hjFKbF7HNbgNX46EO3pc7vAGWnQG4
k1wTs9cw9sA0I+oXtXJkcltVLvjjJmQF14/q1CZkHggw1oX7oq/O4/WrbS+LiTrjRxZ5CfYP9Xsx
6Aa/q3HjLtDQCmwQtKLI9X03aurJ620ONn9q2t6LjIXFUHzT3HNIr4Ejmfwccz9ESTzBX+nekoqj
InCJDkWX8BcVhy8xFe+iT+8lJ3U045tRqvE9Zt3A6vTXbS1tzTraM0Fy5UjypMnw1C7jF3i1eCgR
8qHnTNwbby7mPIPqu5A0N47/LWixu/jZsH1LsjP9hjoJ1u2wOmHYpqXjPYyIcSp7TvGSq29UTGQf
grLMVmQ8kbMa+6KtFWwBiSVUMUvILA5sP7kpp56pUL/uBUQ9AAx4hgtU4N3heWj/yOJMGLBPZS8k
L7FK4Gso7gZOht/lgBMuum5V21zGYhZOouvlOm7F5HrN9PeI/yqwhk8/kORFEeUn75HsWg2PttEx
N7C7YBed+34eEDGLne89N+o/Zi7dtajN7Ne4H375nlbGsN2n42sVhFGZ0TUGNHZ31YCOtLwyPHfF
KTKYhKdNslkxt9VYTiPJTLgyP5OJwmzUfJWvflCK0RlwYy7qECG2L2j+IX40hQYn6elfeUO697Xu
aOVackcFFYlnm0gPrPaR7qfRxto79KgvKpDZgqGjGrko+6ZV0zyuARpKyvZJ5U5PbaSg0kfnXZ6Z
ZPEoLL/lEbtRXHx/AnjkQNpvr5dxlMHdj1fo7kXaSJ876T7MtHW76u7gwk4RWNFDds30Lu5nR6t2
JAc/7C8k7vrQSXQ+o0BUQXc51d3exQML1Wi5Acqk+M8k9eiqTAJBMUbPoapgnf32sBq88dBF636d
CvKpmmG+oTAqdHLmTKVpP4oKq5KWrI+okbSI6CmXklAEFQDAk4w4yDYSB6LpPxRV311nNwEmLCqA
DIrmkejk2BXoZoVniAryf4ZrWqOQ3oShhr47sgzeRfzW0yxI8MWe7VXhnHL7zAXChj3EtFvhFukg
F241cHUXx+4orTH97vZFhcYcsxQvIueD2HdOFQVLXlX8SMSpgrbKYHjrO4tcvWki7Z1NRd8SvRJu
V96PUuzvr6oXNESQvs7toZw6mDoKiee8xD78ftg0N5ONi1GZ3N/zcQ8XdSIP52BMO6WBeHXd+aaA
uWt1HdBt1kgXsQLM79zNlZKqO1AbDJsOV93iSAajhe5m3znlFQCIkwJzEr9oZp5jT1ZIOcuyEJGw
BUlyPNaJnuasPPykGEyqWxwAV0vsLhmnxqxeU/Ii6DeE6UvEf/AvXC8LEd1XP+tU5u+Wb+ZkU+GV
ew2d6yrG01+Cs3czanzSzu0lumsSgwWqIVDPexrEswa9DT/bSeMx4o/QJfHhUtMBP3n3RiK8C1bN
Fnwnfn+KWwK81gh5DnbKm8c9ZJwsC/KmIHEGxOablfAsMNTWxdX/U4UKyyK5PLqRrtf3hjK1FXl3
D2NDb6/ujmT+3se9sPNtdDzdybSZChJdt2NSoiybSVe5Rril9cTy0sLu76t0Ys+Rv0L4agjT03oZ
bzHUmUgAPUW8u8LvJx7Vt7AK+VR2opaydegKSrLBMO/A+8B03Xojp8diY4dzLBFBuLAO4hLazHWr
2FmsZJps+Ul42cz21nk8SWqJXH/71SvhQ2TehslY10vU3aLs3LH7PLpRxbIE9Ih/GY+2DN1F3GYc
z835XMrl2DhsVKQagPYHnXkQLcisp0ylikrjR8pGepJ78C1nJl+U2/jmwR1q7eiyB0cw4CC/dTAA
mcm6JQ4+ksDT1fSvN56bXmGmHebX9MJ3rJMaLuFWvLWBJoccMo0epI76Cxdq5ON2+REFDpH4NKlP
QSqDaUCpGiNBtjZcPkhYsmeBVRSNcwkG6t9DzTRaha9my6mHPaagc/JOyP/1KyIje5C/FG04+HQS
zo0Q8yujLUMy8jnSd84SqM/wVA1VO9o+oUpcTN6q9aaojOHBKUOw760LN0rbprIvobzE7AFWRf9i
XFlU/2+eaXjU6eVjqhDfrZgk5ZyUa/JnOx4md4RQujSKekFbGQf9MHDQAuUSvgE3Nvw33bcYTIKC
Hn22l+TrslbBtCMp1r24uqjHja0Sliqk4hqqxAtZyBZARNkeIKRkWXe/4tgd0OmHrrBDwj0nYWbz
vmE+chd3rF2xllL57ASVF97/51Xno7OOWKGcJsQALQHG3Ed9CsIOYeBvMKYUj24fJJRQxYakzfnf
ZqH6wEWPSa4ixcgdP0yPVCMN4BtPlWgz98KRr4aGM4hVzJNpbXkQyHHuqBRxtyPP7frrYp51M4Vl
z8od6MERzyNqkSnCnNBiGmpB7TXa0mlbqjPKjLl5X5Gm2ZlXaSfWTUypPGvmDbPIJy+eQX8H62Ri
bUtzv98Ix/ctUqBo0YLEOVXeksRZAxTkdAF+6TEGHWGtYkdIY2IpCnNpRUDOsqGkd94/RuR+4oTg
M8NMpUahvQ+RINChVi1vd4ZryDI46gcdGhn0TrGSwlcmJmlAG1qb92bJlUrEmThK+yHwWsfgDlVO
lAZMi9oUoN9XK2u10TcZdIjWSxfmAPssiTdsJcBxjWABTm/1yN4oF524Cq3n9i8QcK/jUhw8e3hY
53CibE30QByPAzuk2jEIXBZHRj+7mmJNOXnTMS+HbGW1VX8NlKC5QXTgUPTsErWDvoX6HfqBv7z1
/XT+UHKiSZ/a867WbkDQBW/kFFLk8ML6/TDfgeIr0GbGxMEGVS+WdhmjLgKVmHk+rHP6v2nuR2rm
9oUPWaa3+0CMzflbdevviJ7vloIX+Kd2Cwobx2sFF64LjWRVm0Rg7jW24bKoj58M2OCOjGUXtIoy
J4aG2sHSXyH8vJcjfMSRS/omL9i+p4a9B0dUMryisNY5HiFoKnJvNSb3RRO3Er+ih7VJXd+b/+V7
CmzS8QpqrA25h43S0PIqrmRBSmXPsyADoj7fAIsI6jysiYIF5eOenF8B7YV/+AyQ23/oYvZduppU
NYso6MpprGOvfnCKxSsiwyijMEnDj3IDZvg6G4tosagtQBJiybsnEniTI9cCChcuDFpKwJ2Jbmoq
mCVePvHjnVd0yoO+xt+wPaiV094T9Cfc7rhVRzBfagIGf3DaYdQ1lt4JZBjap9poUY1oB+102sMC
/vbOvkV/WtKQ2tEASB8xe4BXp+zD5IO70mTJHyranFGpuojeFkGwcB2CDiK0oZpOvit2cuu58NYD
CBHH2uFycoUCuPPDKwR+10dPgTSWRAeOGlBMgZEaKi+R3iwj1/lf7oLE1T0t5DzJAmQKqKh6D5Gz
XAf1GoZL8bLZXmdsyndv1l1UACwG1PLrUOZOF7SP2V1y8f5evxNpAfrMk2eX3JyMxXOG9Eh0VydA
EdyfPdUkMniv6B87WwNkHgAtNGsW5uZpiF8np6klBOPrBXJzwAIUtjovQT4hJXcVKEMLtVAWDZ93
uilO9HAmaySN2i4IpioBXAAhNGr5Nqx7UpIe6XoBfG1FE5GUV7HFx+3Dh5pqKX4gLWTV6JN59/HY
edhb7fb4x04IpYhSwkbIj2J6xRR4Tjq3XOtzdtckSToR0VEVibKH+1lukBgTaWhcOAE6NaGPohnz
Y+PBGMJLVsdbk+S5hrOybfqIGaFH+O49nPilfTbLSkWpwr56MGh51ATvEa2DA7M26m0UhtEZaqGJ
oABdkEUfoDrO41Ay/2Sv+gH6WsGRoh0684Gyu4MjScBxjkx8K1U5HTSEBQxoRTa5+QdAYs77VsAQ
tO8KKsoobmz26BmHNjEQFe9p9lRmpeVdpVmbQOkLOG74h/ohU4qGmAVllt5RpqctCcPHF8HS+fnM
cF5jvjGGGs11CD+gd0S8vIO/5mVAsI2TpPPqWKlbYQi63mQ/yQCjyhTf9usEijt5QsSIPg2mO9VO
7X/hRT8p3Kn6tvx9sh2bygQAxAQkdsL1KKK8bzkw1oM0U9MQJ31p+ntBLxpMn/Wp1U2/BQtAiwlm
IaY9jJ3FWGpQJja6CwCrkKV3v0i+x20E9Pcd+S40CMPUnddVFEaOKQyclTS/0n3g/0IMLav7ihYk
beCqo5iFwT8fSweZU481IXDvg3s8hIe9Gv9mjX0+wGjNxpJkJxZRbPxZJbbNxHA9ufuVO4/tTs5o
xSs/qaAA3PavNUrEuetv5dlivk2sU8dDYCGsj8kPduQ02gd+OdCqu8S79C4qYMNefhjdFfFXEJ7N
7FZ5jBRVAdMbbkaGQCyEFoCXdEJswEBASncvJSdY2vLrv4S3ZmlXDkUSb3OAIhUEECW5+8uDunRF
LmKx/JvfEtwVZjP1umHVkDzEYcMie2DfB9qwjOSb4ZMD5kQ2Xyb12RaYnQdGuYIwwr+YPfY5DJXE
DKjQiGJiEOYctVutBnjGZUtHduBYxufSB3obQklaRDvq5crRUmP7NfwOxN/BKlI5Zby9EQadTSTQ
gQeG22nGM4EyHaV0t2IPyfNnuT08NJYZhyklkGUrRre+axfg3x1Uy6+sQ4LUD8ZUUJDl7quhhQAv
uxamrKUd4ilAtxMcxtwfFYyjA7FwrrGTj9Ef8PxWGuPs9sbndwEkpk54wA4yaN7EUHrfLjO8C2Ge
cXxrXQKbu5h4N4FiAV5KIFqfKEVuQwcTH/0UQfvIoEFzAj1f2knXlsd5HqKrdpJKN2oaFLww5tyh
TnfUE7I5E8v3rZjwoFSPKapoGGw52NMvz4pLh+ZOyAi3dU4d9AInQx0gGzU3eWCHjDLqKqdAVggN
/j7aNKfENQs6B8mlZzjSwcQMuBUHS0yFfiV7Sd0i4xlzb790AF4a7690oK+ZMw/08eHxV8aq9fIR
vfg/F7gvtCofODqjwMn1Zfe3c1Gk2e2W1wuDgotXAMqoMWeRzEUDJZe2I2eUft8WtvM/hKkzrMBm
G1s/eMRErjNxDeHDL0ZdvHAiWk2+0bqdOdhBdkQ0yuLPRFoQ2hc6ByiGye52LF7X0hpzWqhZHsnY
kkJFYL7/RL/26cglQ9iz3ygvwvcC2fXkAuOlY+n/PYxs2ZRtxSa2aVU3rxskXe1tb/kDQHTnbJ79
MuWp/u1SGhevwwQPjW7dCWNVEVKDlnl07ZSvsKobJZ99r5O187+XOsP7IlcQohTZEdXSz0BbcOyA
PT5+Z78mMI4GZC7N7bjqUona/srSbGo2Aed0IYAH7mGPbIa5uVhgYcSLrOJexhy4Up/xH/2u+Dmd
fWnTO3liWDRNSTEKeE4C47SdGDgSzAKdQPtxIMyFGXev5WCc3XlAFgUiNsD/kpzxbiuuGjCR5O8k
2yv3vwDzU/p8iXpnVsGKe6irwk5bGDxPtwNxmxovuiyIpPCjGvG8OLuGeJcekFxxV0FVq29GJ9Sd
Zx6amdh9EWPA46WBQzgPNbnrGg4ocGwRNM9vfWv9w4/Nz+Wf9w2mjusziYn/QS+rBJORE+tpL0MC
s2WW8CyhIPg4bSyfuerZAAavjj172UAj4BHdTIOxchSKMbHybNOVQ5/ZAlct7t6IWxFim+Jj7oEb
k7wDxVeOoEmcoSid0zwrm7NoYWo7ZnOm7TGYrPyMk3ENMGxRzHBDrN/Y7E+Wh5ylRjk9EbPOwZJg
bn0tDnshfznx8F9TwWI7KsmAaQicoBq/pdqLNl6Sa0JVRhJ9NlA6FHHsoEW9Gc5FzKUSc5jTOJ0z
ZK2URSwpG9VkhEpIlbadigsm4VQDIHp5ngJHQ10j51Rd+pyByMXFB1CVrS5IsBdfcXF4bUYzyml6
8TGqJIJ7cdrXe6YN8M8l0kKZhiOCFKqanxQBTyaLUI3LF7I8H9pmKipe93I5GJ59WW3NAbK1/bsg
knJfIKY92jhokubtW/pb9fuPXW+C7VYc6phCYp9GGNxeWoYZqKpWCP4+3KwYSY+lYWHpVB7OCuda
PhHOzzqywagqNO3GURi+fWvx+UtQXIqzXwnoMasBcB9ulyl5gr1qzlrO80m0qKLisFroCDw+80Gg
d4s6uZhmEiTDyEvfneDy4CmlcUbxfuTjy0CH2VmvM4GMO82O1dwRJivzj2IKb6aIRNwiTtCPOxoK
oTIVPQrAinY5W+0VMGe4Uab1WxSbMUfSgV3VwbmE4NZtzQ+VVfDdlSTYADyoMvU3lVSbNpSnwFpz
sG4IOJres06N44ZbzG0ZwqEjLl2d8MTYrozbPJg+7Adb9HblKjVhbgRhxONO7D2/FE5E4HjH8/YP
H8cgmyD4R+Oz0DmRS3ZF/WOjNoblCQz4gsIs084ntg6WW1v0UHONfJsNmh+KWD2ecbfmwqP+Xb+N
x4s+wSCNv3fTRXOkqBGgGl6SyK9sm8mhBWWiFX4rWMEtFYFu0DaTCmIeut6RB708/R8ADIxovu0S
2si6aVyd+BMeO0/D78J+Eiz2geQQLGctS7G2Ks1satVm6WGEHgD2fEt30NyvE3kaLd+USZn3WxnT
oV/jcpnPaNWDzajQyKELTYpj6rbenthPEs3+2bLKU9MhDpBJ63jtIZXtcavLsbKjd7Ebxwd7vCNP
F9ph2kQJGSnoqntrXOua+qpzX5PkIvOiDj/+UShiSvRISsgb8WpwVChzi32acnmmomDjusSur7uh
8hxP0NHNT/lll+rDRl+nn8gdTKYbZA0W02JIet3FRrRjRGI6RZnsvH0Xj5jQTcCqmVTj3D9+EHks
S5Cm5zVnvTghGYUgBmRDGQv7/CZj5aeo9az5z1QSv2FysDNUygKKOLxAAR3+Lu00lJrr72IgF6js
lvHL7TSdJLOtU7NMWliH6rSSGkXkyEHg0Us+OUKdfIoZ/GDZsU82G0z+kDqye7pDpZ0tKo63NtwM
/hqvt/Nr5nhzOQdBaNYuBjfWWLBfSaK2Qa0kB7UA+CFLEKpeMrPpF8IanmGPfq2Ob2D9SuqszOhP
VtooyXPPeIppOUVrl2vMJUyrLpm4ptGYFANiFazXs+6KGKoTZly4xddPTz2Qxh6oHuJjICireo16
gABilS2dq+SVw6E6K2lKllel5zbxvWU/swUHCAGhTzvJJqjPcE0IcwP7gCTGLBBrfJj+P5YHNMOs
mggbPw74bAT2ztJpqW/fwS3OE0PIwG7cWUIlyy1kuf+ODbypIcb2rhd8uFI2M3Lh9nvvVWAFEreu
LQ6f3d43+HubsXzccZK1AB5rK/1C/UjaBqZfn5p/jd4+Srdvm0p+JFUjhRXheICswkcO7uksnJiA
77/CUEGVJSilOr5mF4K4BsXSr7BolvoqozzNU++dZHfaaUjkFWLtMDmzi3z2ngUfffyFWoa9NCrR
1SGnOIPtnBjqnazlDP7HUU2AXqN/Ib8WFVv0vpinjM/+yuLz0J3Sw6UtxnjH/5uXIZ3IeWv00jJq
kqZVhaeNoK9a+yUAVdmUk6g/01gWCjoGTefQ2/5KmNwgyAb7pmmqBMLv+n2VktEgshDuSKDRpjiN
fcDkWycVGi5PzHQQXXHECBc7QRTxYGJR9aYLrNFITerkIux0ET4CtEgSpqOdR/ebzHCBwZ9EUlKP
aOdydD0/G0muKDm8AwCO/5JTKXoBUg2h1d89KY8jJMTDHdeGySxMogR7uRl2iTCxc4Fh3G+ybMye
7prIG6CGDSnBtvHDjKW37z9uShHDsDy5AZg5wds8rIM+16rka3HU4Nr5rkwgDeVEEW+sh5GsqYH7
YuoGS3cE0Mlsu1w/u/opmrmvy7XWA8E9hVLzA6uF60I6blmzEObkylu40pMJ5nfFJKy1/rj5ypVL
zF6TMAAb00W51qt37fXb5ThjD1zqjwZ0s3Y4MQq30azjzNaVhf24UtB4PILNQNYtip7FVKDWqXzh
HxXS5l9jmKSwivV4xK+Wl1TtjYdv/SxBox5Ucq7OIfAwArCUcIfJjL7zRyxHdVftVe3+GS+TsGbA
KqQRQKiqnjEW0R94dfLj2f4oQsGpDYzpbCKwIqYy501It6ohXFWqxAKxt8WbmTB4Xv+cUxhb5VKP
UF7bamTxz11v9c2CJoqEKgF3jx/lx3AIbRtgDe/5vshBDzBCUNwtgGXcs0zjeYod3QWjQMCLDBhk
5qDBK/jHIsTIoEUraqQhr/NqtEmKLJ237s0geaI0pE9N582fiwrn58jEcLRKSPXXduSEU/gEY9pj
yYY/oz2YDspEKncSIiZA4fWjmPRVg3m2TNboQjuaHXW59Gtsu9IESJbf+U3zTnrv+87QZy3X5dqA
/rGDt+oiPVtDMVwihtJTkxy9KNCecvDYCoq2WKdpDp4Tn84bJiK7cAWtxiRO6fRJzs17fAqgtdSD
o0lJX/6QCbCK1AbUSbJJsuD0feLvGgmuHdb4FdEpsMfjoxwMNWL89B0888uNc2iG66rTQf6fhd9R
5uulnykb0uXPSkYoh9UJ1SgIfnx9kQtbtvz3h4RCS9dhSpJoq1BZ83C8ImucsZnDoxK2B42lXk10
gNPpOpIvYBhsHd3XKl4zGEK1CGdldpuQOO8PF3vdTJZkLsYYRArSUhYvxBxpevf3a5oLSMwduicq
5KvHpZKstKxRsdEpMbp9sjNkmXy66wLljUGTwUfhktRvb0rgVen+teZNqYQ6BhrLBZwpsz+uyO7H
HFQxBUle7VQ5tqGRvByUcRCyJJu5K5mqpjv7LCLz+KXZZZ6XqiT/SD3Wx7viUd1xuI3vmf+XetAn
1A2R35sEdBjI2pC4h2Fz9zBuH/4Gkn+6C+Zguz+chzM7ErJN3slkv39cp96kmi3/WPkVX+MrbTH3
K74SLv0V394Vbu/RBECV84nlslNnx4s7kJp7ttw0WH8+PQSeAtY3MzFfpRCR1YdYorxU8P3QHQf8
YOGrLQD8Vwej7PAgtOKyUcN0Ny8St61IMxYcuOGGNTf0Ju4IZwoSE0thmUmUPXaPNdbnB0+kSQ0L
yJqoptNJTNnOiFLoxgA0TrxbG0GHeOiiIKAGYu1wI94BnutdK8cy9OBmnwnNp14tE/IDLkp4TaNL
pmHucjV5gSm13X1OWALp7KwWUvzFTqhHtQRAKu/12qEIpZ51m9/zJOs0QIxY7AZZZ7BGgIOhA549
Kv93dtWnKNr9oWaD49q0U9YsINhFknTpyLp5Cou7OvKz78OweSWtrZ8odZEak8OlFbA8AaW0aN+0
eDyQCdFHMg1GKBxUELj4M7+PGvvqlMsY1PfGqQ53rK2E57Q+02gVQyJS+tJo7gQR25t70Bmc4L0I
4wEZ385XjOqhb6TZtOU56jtMJNC6LA2hBycLnkHD0hJvhADhE9ils+LnLiZi5RwzLlhme1xOuH6H
FuTbrgHRC+/xLCweZFhbWfEQvkbPfA8aMUNvsDZbIpr2QzPi801EhRJzP14g2Rz0CKk6lNmigxes
PHeDJyrSdkeaR7VFCLp9/HFq/41KqZDMWBcrj7wn1o5c9vjdgaQlUeF6EQMtTw/hLQTF4Q23JneT
1UdGJJEWyV3pSbRa5hkqfmugJXDt7N1DP7kFN4f9+ADoodHUnyGGFBgJkTpkyxnMeGwV0RXGBBsP
iYgYp3TGXjy5omPmcV9rZEoC6oipTAq6ViDATQwVFRrWfgfvzQLUOLYrs0u7ROsDqSXyapoFSloN
U50b/a4cSk1TGOZbm+UmMf1nUiDyBTuyEwEQckbkuxegYayvFvu28OP3/KBo7c+KnlwLfsZ1PM0S
rar9gkfbnD81IORrlta/1ZSg6yTgTnjDESc+Y9trE4zCiBxGtx5HSlIp6CM7aqnl8zAYbuaGHd4G
YrpLgWjy1dongFEjFp6f6wJt9kDrwFAe1GTX/LHuZMUf1kXOLHtBBuQsDOXhZKkh+RmgHgMrnopl
mwUyqgnAA77vkG3RKoes2D6X+AdVMLPzzSBS3V11RtfGoz99h8456OMvx9bg68uUmMn0TX77dC/r
aAoEPeNLX6hKD/kjhE6Gp+C2zArq0stBolJ2ol5SPOzfD7GnCAJvoSGb/BHi5phGBGaGGuaIKH7K
bi0jd+BZ3jB7yZIDZfTfzuWrosbMgdHIMEZbVojegp8ZtV8xRHgim1M32ftJ1tWlV34ycREQjyxr
Oyb8w1TTNlmunAencin1Mvd6B1rmnvra2hLcHxdnbY/MCnLAMlbYtRRGNQdqiiojNv6/RzpYvyM1
kSe2K2Is0ta8EJvw8vWtarba4leyNnwWwNRyM0KXYb7PRtmcsAq7+eR1u3LLyb5fBapXHQ7dQtiO
0zrqo9ycYDFeZvyIPc+rZDi9KsRNkhx8lpXTct6SmTPWD0j4rmqJLkaNYIXmgtahlZBpExVYFNIc
7rJCB+b2pBOOgkEgDQZsTmyo6uV8EV/6yE529E9Hlzcht+3WyVFBMBjZQ+fu4YPc8qu6A740sq/a
a4g997x7kSC8fLEOIfdI5XNfaEGaCVNyZzB2mBqgdQsgj7JHc2q936G91+GE8Pc1ctAdxxuNpFxx
HLjcIJuRtsK15KjEmlTHmWI7qNS3q/2GuCG8kJ7S6JPk8CkYSycrNgktzkTGfR8fpQqeGzmWov1P
bjUeBWHZTP9EyQntISFZ7kPwnZdDmHPsS/Y01rzCmptSESuthuWzeMd48jgmsbCLnF9xeqNAQh09
munDVIezem37SGXeLaM6ecSF/c5IF7asU/fUdedAQa+N1xdQqM+u7/k8rx+1AUkOGR9e7D5cULYw
Vyvgfclnc+TRaqg6QjmYxWbhcj0CHQJLL9SxffqEft+uKF+qtnVPpLOst/MLmZ9H2foR+6OQSL+T
qgcU7i0S0d1Q540+H2Ra21rQtnUDjb0eWWFqiShgS2NGropj1/p1yaL/D6oTb9feKtt4EXfofXZ9
7ujNDiy81r22bVi7xDzSG9jf4OqYCtlMoVMGQ/JB5fjwTDqwpRZx/4NgQQscvVpzgO3bFK86O1OL
17vjojsFyVxhHh18qszhd442ZpB+sPE3dEB+HFizUDaf4q61nPHr8zzzZbYyujxyrYwurfyS4PmV
GxuPRAjx0Nxz4QE148dFF/mWslq6JOx3yu/8c1ELHPF0vOagFPDHxRv7mo9MbpQj+KpRfewjba/n
53xX1lkwOeFhJn6reYsaeerPmlhAiQ3Im8DXP9xiFP9UiJG9uQMTucHPdUIudd5CVCWmchg0sGvF
m0KjB3VqpElMGsyi511uL6m2/RIxbpPo3gPUB1E9u536ckTPDeb2WdQl8PIDBvchOOD80R8HeV26
6VFeepvJlj2ofqKNDM76sUiyFfnNkeGuqr5jaoGgsh0lmcbyOu2GnspZ6jTOQAUaDuJZuORnHvqm
DOHu7UDnBW4qgrnaFSCjeZAN9ROMClaJnDQmsSppFefGg4xgFcjOB5UAoxkFYQejw3HC3zSq/0Rw
Ol1a750BEvk0FW3/iVlQC1bCjkLBKJjr5BAQj+qvmpeQUFDfB7w/Zfn5xF6TWUIRFa6s/wBDI29u
KKFP1e6A/VY2vlk53MKUSg9kPxBPBrmAXpTI1DWIUae7594NEZWQJ3oeWWVKE8T8q00VFRy2jX4Z
xYBHQ1eUS4bgLszHDlRoO2U2GbaOoVYiQ411tPHsCzl+rGbQ77E4iNidfL/9OKTdRFK8GZbTZ+r7
5Ak78P6QRVkE24gB4sDImMw4ylvd+WiIaOfxNagazsKPDtbm9d72AhIqUs3IJ1GBNI6MJP96zVAj
ZgbbXKLydmjNkiG7OJyDSARNPZLQpsyYciNrzvExbabcGo/TEuNFaz/6gNUASxA822iYNDQFc0vw
O2xavHwVl5g70xRO77vf0Cummp+KMFT6byBwXUgFjzqjus+9UOZdA0QwDbCUCNYx9E2s0j6Bs/4z
fHKzKfi2+NOTnPq2iv15EFA6Z/0SUhua7UhP/gmgzMzUceOmb4pzEGYO7cn7F+Sx2QOQKk2je1uT
tz97qF3ASrD9UHBGB/y6dHRVhmxHRa14sE8Z48bRUU55hVPL8tjVRxwqe5lAodZ1fgKy6irpkqA9
Lp3fs1dLvLIAneM6wwGh/gUVXXeQ/O1NRmDiIJPv5mg5lD7EU2k8a/q2NGD/bpyC0F1+8wcjrFN1
hN4mEFfgfLzRAocyTw+wGEDAL4ocoLOTmrMDnsCJV3jtFAW+zKUGo0FjswVl2QPzrVas5sFTuNY4
kbk5jQsMiwuT5wJMpgUWHDFxjSQYJ1mMzfu3F21ZKue4aNGEeyK/7Z9mLRZ7E0M9tl5zobC9H2rh
tGTOtNztMLahrVOU4VnXEbxD3cfzR1f/SWroU7I3S9HPpwC3CX5Lc5hRKHuCcGjn0PzGnxIrwZyO
jJoLNUBlvK7ZMhm4p4vURxvaapOa6MuyZ0pDuG7KwltZ0I0NimbGPQfQHRw/vNufOpXmEnTEQ5z/
BB5PtehpWCm0JBfJIprbb3dd1635PwuIj90c/CkvHzkBAsv13+sin1eWYVjpXNJ28/Y6Zn9lqGow
Vbr8W9HlhmR61mEq2MFqRqn+hkIcAal4G6GU4DnquCa35Xhm+zWWe1bBXk9Jpao58i1I03nOqQCG
qdtIAEvsRLHN3GN2rJCoNT3hMmBXMB9YM57QNuQGzNE/TFbbfIzUdHo94DqR3lddg3CMrcCO5sx7
tS5YenQbGPuLiyJEtfaRNy85K5oTdRCH1uuyNre0o2lvGjwT5Any2z5PdH2o/MeFHFI7sSLI8aO9
VDgHGtIzbnDb3DjihDXVd/jOQROVGukun5+jYlUh7E4+yqWYms/chfRC7zisVQ+DhCK7BQoqBb2y
kKqmEjLbQOoUDN6kapc3yt8jVsfUu1RzGNxPVJUo1uvM3qDPzMn/VIufMSLNgUwgkTbaUeYzVIB0
SKUyCG+qIkMgegCWxyXhrVcWOhJFT5VqQ68ABrZvh7McK2mbfmJKY2omALEv7ZB7Rw5QSlP6Aqu2
dggdOx/UKFHNfeIFMiQEfrA5K4lD9Nkp5ytBaBxUhzNT8teeamGiuu7lY1COwME+0DsHtUJBl8J4
b1PDa6CcvvqM+HcKFBsTYQJsjIYWsn+SAZow3gvKKWwOcrlz8Hj16DT7NaS58YsQnjfsutUzp0Jc
zkdlhae+kyeI0b4ELY+qi7vYB87I6AhNEBkFRc95SeyloqvF5MBUhn2rmzAtRNyZb8gmhwt7oTHV
xFpj4GDi8IFYfVGeuyR0L4Ew3ds3NgEtDRYVAxDtbFn1Q+kHLsFBQqhF7B/zgmBUMNc4dyMFYBzg
SG0NVMVwVOZf4lLpk6fWiSreY9e1KHB+uq8ZYU44x1Q4u3DghWy2Bj2/+pP1aXCw24S5T4Wpdea5
poXy2s9yq48kiEAjLF+DT9wXSOrlTTb8CXLGIZNmD8D/dlkx018H+FEAYEdP6mtnYF9G54V0A9SN
VTkMpg3N52zUwclC3NI7y5D+kbXwy7++v9pIf15MIJYLIRQPoXWwQnpYf5NcRuxmdHgZm9FWpTye
ooaaQ7E3Mx2RkpP90c4k1aDiMza4rwURsO/2OupgsW/Yx1BvrnvlJJVR19/vYUC76OTtiugETfR7
yD1HJSmxcD+qqPYN0sWdi0vSfJuUJsUAsTNzPMrxMn5wq0Ttchgm/rgRxCqsv4cTpdWHAYU5O5zU
101BGyrvsRnedL0xNUcveY8otKQj5Gw8tbJ58dDEOnuTK5WkdCjFlJxF8DCCh/pzAzMvA2gMSlIE
D15jkd2upr7aoWUmYAsn4afF0KJNoxSC1404Hw5LD8y0+JnnTQCNVcbO9Hlbwziadj6SpN/aoy0W
KI5iRIHcK1WTqvcYzPvuj0ixa2onB5evh0R/4TXFsPSAEKU7yZaFVevW+bhczcaSsoKAktX+1aAi
SugJ41OLJLtK4r/F/VhHGu1M5abbq4sear6wYOJNxEGnM4lBeeFk1Z9n5HeaY6Po9ZlJZmXXNauQ
JmMP640045XybHSMJLAtnQQwIx2vXWhMdlHf+qnf2pWeuOUJoQ/sTRzDDk3Eum96kyiMvMlc9scq
9RxJzMM8wZkGnXP0eXaSsdNuDKPJ+W14AtUcQHHm4yOdiVfyWZgQW4EoF1Dsh0cn0AygzKd20C7e
wBdRLanij1ZlWTiksyQiJdcu39PFoE2bTpugVGjL5sznjvcPrKcLrP1+k1TIqN949RFcINmvANYY
f+OB+rKzQ1FNXXT3QUzQqxM4qTxn+n2fGyeFAx24CcmsXCld33LWLhjcyfBl7lPx27HpnFRqkhIU
9jUXbl4pem598bIY0qdugM7/WyUQMQw24gdhMQAL/BGZKajFka5A0HjDtk69rMCsMNE/Hg8kSd17
7acZ7B7zGTCpL5GILuN48GgSdJKMVd4pas8VLOtWEHnNayBeZj2H4H6ToW58LLNPnLcXExCFPFz9
7XH4+NoIlZM35uWVPTlj+sBWPijOmKFAZJNRIOTVS8JlP3u9zMLMt/DaoVzdJb5gv73DI1EJ07IN
WFsQJoY0tlPmn0qRYO0g72MkME5/eLoQeK04nH1wZ7DWg/Yht79x/yMzycHTRuvQeGgYpkqp6rZV
AY2f0daWNiGXKGodre4CJt7BUY48UP33tgybbM+myq29QRdPuQEXHRMR1XFZFEpl0RBU8yEU86L4
++3agptCOu3HfFo1f9/s8NHikWH0FBQ0NpwbBllQK8pvh8GOZ0DweXFm55vTp/3IgGuIZIgvirZk
jZ9UKUIvmXyQrebn5yByE0Sihs3Jwp/HNosZCMd0Hpa6H4qDOfvKkSnT7HEKF4+FYpSo02iQDEPc
vwMZLV7aVSUY8NIQujb3L7uL6T7x/zZRgGD0qcnZdPcvbRffUjYCIPnXDhSVndWOq+wxl8CFghPv
+hixHQ8YCnQMz2eIipeILiFOA3sYnsa0aqu8WnAjqbooed1ObAkd6adcYczyJa6KzqUQ18ZcRYAw
2ZgBMnLIqsxCC/xRfCuvcwhpxKMZujVYxy8mhxckLXkB7CRNdsrdbItR/UfPpMkOqP8/dX8xB/i1
gJRUfSKPgXcjsl82DFy1lnm5HN36GrlXt/XT9I0n7lch+nVrXQU5IqCSAf96a0C1LI485qBljAJc
jbZ7z0iayjdPDsSO4ZGKIT+PqGC59yldNCWTtKKcUDuRPEoPKMYzEmibP7T92gVitWMlzU9/CPvG
seF6MOkAzETAevPc/WS3CMVRRSnttYZvJYi2sUQAc3l8xycfokAFvQ+Uhq7Gp9GkPPus1c8ahOHY
828+8AoIXHQfSVnVPN6vB7JSfIR8lA0ONEAXxmpJECscxn+EqJGky1exWrFm5u5jKD/x2KVWrhzo
ilAtfL2BryArHwZCM1kMIRAs68jz2jkDrtOeu8R2+IaV4j7hnwwLTLbrDf7++k/g6rNk2+5yFbP6
4nBEL4OEUYZFMQcyEuzl0zceACPVuHJnNMK1iBsex3xp7CVUKXeAZrUk9ZQea9baCQHwGzh9LAgH
7EjWUUJCJbPwrL7chzBtORpDjpcI4G1focv6Gi+H/CkZj6FnbgiVKJhH6ESawADbQj/eRxG5ieX/
teINlHSoGOUgI29Ri1GU3adwDEMbNzRx8EY17wTkWcviu+tkIwOaRBsJvAQ7HECToeWxT4yGznUq
G3c64bCDaGlPtD2hbDrKhaIp9hDbmr80tNjds88mcocW/QC8QxmxTXUXyVwKF8yZRUvyCGakCmFT
b/6Csoqdr1sEJK4ChL0ELkNdEaDS3z0/b/UJHEdTC9QBYjirU517r8aUBH7N+d0knfihrEmWHZrn
b+QRCdTxLFoLbXaek3439lTmpz73PfFkvqAyzIomoPGHgXzVpej+OH6yB+ua5ERfG3UeVKoBgYlT
vIwjg9pU7x5uWgRuzKGvYGkViL/VikYFmz5wqzxOQ6e8zHXPRboqM86joROMWMVdyiWudohyU8Yg
Eacgi4D/d4AeJ1XX1IK3vu014bWpLGaqK1t2BmLwGCy6SyiHEx8hzDGKOzSVlTISzosr9iOlLgzl
WmilMPNzTyK6OIjbfNarR/kvLOHePy10FSlt/FDZ9zx6Qlc4Ohtr5+/HJgNbUeiOpmg6ewcMFcGe
FReA9H7d4AwLINQl2mbsvF3sDo+pNHzAKmS4sIODv616yGy2p6Fw0lJ8EPcOJQtBBFRObSyxNac+
h1Ydco2LNi1f8bmr28X6ZE3Qs89XFNmG4fAn2qztRxcF44co6ICqd38lnXhoCATthXia3KucIIJ8
y+dpZU/wqwh94RvIQniBTA0pIEl7N/CDqQydylp1y+gtGzLyhnjvyt4hFqyiUINd+0XAnQ8e/trN
bW1zBkWcAX3gwu+i9QR1eIrFegzczdS+q3CiWLBmA6cBUF+7eKAgezJ7yxaIwq999eAcyWl4mzHm
1eW6+Om7CkrGoJh1F+zNkMBJ8lUeXGfQl76sfm1VYwFYA3tzyjNWVzcfVaa7A9YSOhiK6lvCePTt
GZjbYnqsi4tLDCAkGHco5wLaUy1gCBJzkodbeVBSVuIJuEVF8UkZE1WwRt8qLFx1zmA9S/zSi+Pf
24d+QKw0eMucM2UfeAntct5nbUSnHioYMXz+3DWm64UQAutmHV0N1fFO8n7X1F0jniHMmCO/gT+F
40w6MAvZFFRAb62GgS75o5NF0B6P2PavmjW7Amzzlq/RyQfBB5eCxpuUEFgWwSGmSzXeKE5xZdEc
c+ny7rsLlQ8U7zq3FFrQXGRCLCK3v+5RYFfFNM3hZTEXHlybHrXhaWNQxmoMIl4H/wBcedmuecoN
RWlSDgnoTvHdRVTDiVBUYPWJWStuVER/JG5nwD7nFaWhewu3YbZD4CvuDzDJDLPmvJISH3e0jSPU
G6DGf6BxWh9WAwsvjz0FJO2iW7Qp0ZBEXb5fw10jkOISmVlLOVUkbUGwbQzDV3hGw/az8hHBaFD7
GYSHG0e8F6lqs5QtlGfGOoa93yaKfktevV9sLRb49ZPH7I5EHRZ2x/V1E82lSunzwDCgHVQ1oRzp
potOg3rFu/7Dkk4k9syAhfyMySvPBRPkCjTs6q7OEhagq/U8ZcqrLuaPNwQDxmumNfjzCrT7B2qI
idwXFcy/O17CIWTVjtM70v/FgtNkJi0ye5MUPMW8CD6EmiL/6M+7LHljx3hZmHww63bF4nWvAw1+
tchm0DZZw8hfYpgh7hPFiq99/2TROd3WR3sQH06Iihb+5bohPp+okLWBWbsvwhf0OtYF4+ZJy/oO
OEQBsz2Z+tTVSz5EkfHZvAhVkZ20chG65+lk4PNMUA3CFCM291wOjur9jOXpGXCRouearGbVycc+
TMi/nKzgFZOHXbXyyBp2kz6VI123SsxG4Rv8bV/O+sEk1cm18tmLyhcWR4HYTlxRYsu53YRIhM3P
9BAMk7ulzFdz+VHjpuYHFSRxg964fWk2ECFVPpP6oh8I2ghy0Yg7gU4QrpNWU85irJo4D8uvthxG
Vbz0LdO0BX0C4H+QbFcPninCBQesGvbRUk2aa8hMuCCl6xIVKES3+dWqDW65QIuoNvr/wUDG8QKW
/9VXhzj52Rxsiwa7MRjJ78mPFGG3BpJa8XINfbF2XjTPMlDFiK7mEC29Tur0RtgO7II90ydkEZIu
NvgItl+Kmoy/arZy1t8oP0DxMhHhXYGbaAGNJIhgrDS5eUmX45x8NTkPBS8szvvkTeK1XXSmru9B
CyvxrcBKf/umHGu7bsemGasrRQLizaD2HDCDUuLyXYi5pzUKasQYNweVi0gKJifX7oD8Q1S3ITuT
GfOjSa8z9HK7R1EeO0dMFdvgS+rVj0zh0XR6n/Ovl02C7MUvz8YGwoNVtJmb2leXWKYgbvjDeuB6
bJfxzbfz1TbYyU7MOJoYdVR74O2XRQQusVIpVZoRfIXTKaiDGgl+WSgbQkoelztixTx9KNvT+8b/
Kr5VQOH0fRAeoDNBVgdhAXDI/GQ4rV66P+cs8R2OdkVscMXgejRZblbP4BTKJDdHB0FHecYgS+c5
Y3MWr3/0Zp3PhRbRjUFohzfkwn8tK/kR6nw6llwb8+SvNhvAX4OQ0shJE7vfwrX2PQfF2NAaf0E9
zi8VO8ZXlojtkxySOzkSPd5q/Pf8kPj7/Z2tpNwN8D5rDOCPdaloo6T1fs/eBuupPEpwkMdI0H+e
3ILN+un2yEHokV0ytSUruSH10JMb+UPUssOtDJ++9/3Yrb5T/rmS4rAiCeFh7giffdsVY8gXbfxY
B77Ca7WcXJxLSC+kgTY/1fzRcDpBMXRwX3kFNJQmFZNJDdsXdKzrHUsu3huExzNG3KWuVoFolgdv
L7Ukra67QkyWGCwXKljfCzPcyMl7p0e/3Fc/uWCysSVyVu2yyHKU03WGFLuj2N045tMDq6tHnd6K
Fh5/QtW4Hglj0/0fGUyzsONwMwJOc3zxwWcZmQgkz59uygdHAS/yE6u5Gp52lco4uBxHGdTmrmJx
xB4ybquknFJuzxakRkamdeuPyqNVgdpTDwWnYjwb4+nabG5u34ZlMZRkbo0QY/6KHSl2Gwue3VVN
Yp4BGB4GUDH4iF00aqbGjRiiJZk2mvwiqjhuIYWgSELK9IKYwQ8KhXPbEQofVonFLGwa1Dz/VCRN
xXHdeKr3cCfEFHSRJP0rRqgzMOjq9AZkmGNvFXU3+D/10E67hqCNHoFCtlo+9zoINX5rV5RGMVid
PhwgDjRVR6W5m7Aljv9b2RT8+4yrY3euw48MuMS1N3j2sbonF0ymUxZ9BYD5e7783fey0WZb8Qhx
Q8X7TOGtAcpDnh38n22d26BN4tHDeYccCzR6Q637XJEZ82egqC8aEpeazzaNHyg+7oBipsWZS2D2
DBPWOkU6pmHyr9qfMrvxMoiOsb3BNJQpvblgZIQzriCxIr5WeZCsn8I0L7oVXx/KEv3txKBpn5m7
gcqmGp6JJsI+q44zyRb8r6AYLnP9w68lVz9C/jYpMmwzPCUtj/eCQvWJOrJ3CTjbcWMRi+8LcGwn
Ywmid/DckK0CshxvKt3f79OmsQu+4Mwe7CB8biHkYR4FbtZUvQWCjzIiq+uYXEPf8PhiSasNzfAa
BqstWiTaimx/EYxJtlfEIky6HeFcu3VGL0pplfEFUMvtXYmsv1CONR5UoLdVWfBrhl4lmdyhE5Ia
5nLRT/OBCYH9q+CbSII2PZb3iM4rmId+qEi5JSOR0rfSO16uqpJOKWmK+jNeUiTp8u7xjcKW3XUo
su7cE/SRPuqRsTz6gT3aagfnUrstFHLKQH3Y2ONMlvYPcj4f5FEIBkdTT6DBSHVvdQDOWJ0FyO63
EKqBl46lB7xrjqiVArgHhTgV05ZcCY/CGwxy8luN1RNLPr6C5gqqoDsXFgtLECCrmbj86m2JSGxA
/YxN2KAwomOToDO3hUwtuyVjAsmlRVHAZX5dxbNHRoFH2uSTnwd1voUp1BzJG63Pn6Cuht0T8DCw
esUazY+Yb1Wkz5OTXbhjaf2v6aoWbdpUzp5+yONWdE0dzWILYCSQWVPGFJuB1msIKG3lmnlTavdg
LW61EZVk37NtK1XbxWaiJTlyOpHovSys9YvYpXGTHnkd+u9ApC0u99y+Tt4w0qw0/Tkf+rGwL5al
rHIZtdg0nmoACR/iYhORHhOrq3S9SsjvR6Ydletwyiz+QiFcWu1C/FKFLBGMNrniyfM40rVxqK+Y
x+7SM1dOxfVhMBdHs01bf2Zv0atYHb072tIzqFXL1MEyGsgRZjUSr9RbvzHYiZGvP2jhbPcZv1Ab
aFjeBEhyaba88ch+kOx++qFMf7cmd7hfuGLbuO+5vqVD4yWsZFPf99wmNJHmTCUg+AH4miJBwsIm
U+jdCKFeDkSirz64P6Fku6gwsnFVcdhAmGKZCFQirw7PrTO6EAlXrCPbmm2QGt0ROgA2miSGj8er
iSBN2kSQjc3oP+vwyOno1FpLxMSzBrDXB3yrdz6Fc0Z2kF5R6xThJcOh323CKQXFcPbb0joHPXnA
4S0db3cWqtJugg5YbM+5c2q9yIU2LfQqh1WhhYe3ug2EIAub5qrjChbIsvNMJ7j4gcOOunAmDLSl
swYv5f35/SixLliDCWn/LxEvCikUVpLj4WsB4S2qeBbGe4/JO8Cn22CDqH7PDb0uKVcCYo3otQO5
nCxnzZzpPCBcjBJoaWbAD4l1p6/W8F9yD9TwCQqpvy1mTG8/iJlITd05zw8G5YABDj7nxix/ViwL
kB54qNRGM+jF3NtcRrMRIFYSF1PfdPg0d2NuBG+va8TwPczNOGn1LufwdQTSNUspFm3gwmrYuHWI
f9rFKU96HeB+7dcDzkhbVjuXiXwKk6Zreg9/zRsJdWwoWRRw0jPAvO6GcTMo5+lONAaME4ByhBMN
wrrYQoQrDTCYuyziyyXdvVzHReeToBfoH47yp4G3aH1/xXDykSiwpbM9xD9seDwm9vV6nvVGsOGc
hp8Bgy5oAyFP8bQ6/b0R2J2xg3OLNGzilnO/av46iZ1TPNMeNmGijbLr+f7NF/HYdRGaprn7dTbD
eSaeF49Q8l2Je6pok1LaT47LdyNU/N20GpkZ4FiMXQYM5ub+sDI0SJ1v2CnJYk/fFpNLJS59Kafp
Z/MxdtSMAMHBWXqa/a9h8o0N0upOogVW4HL/LTkZTaXtJXI0OeqGyEaECdca9aJ9k3Ihzl7wsVp2
qOn/46slWy9g/X86rLK6Lg9zdJT5qKn4h2nvf1OEkhxs33Xs4MwjtGoVoC3/aDd/gD23QdEK1b12
SL8C0XNlbciqGZbeX4Nivf67mr75wEH1QGj7aTW9g1JTDZIIRcblo3RtKSS7DrOYqN/552GM7ph8
7ih1Lihry+q1mWA+1xWzQZm8eUMYs/2b/IM4NHLNaE/h5UMofWLUSftBPE/oUodHfyQ/14cxqYYf
MOmmkteaY+bYNsgZhcAKrQb1k6xjyNQ1+LFgK/s5jsGf2np1SlWB0WlEucgqmqDwEwvf2Bn1td4u
CmQywERgElW2bdzhwI2X59xYjESpOVvKgPytClQ6jLxj1FWRAoNrVv5b7WF0CvCFFFuQnYJUwXmd
0kVtnUlCT195SRfDCrv6ig8HCysqTlNiwj1P2oVENYg+jrf7D7I3GSnv1QLK35f7pJ/R9fP8tTgj
qdxb5d/cstyBg5iP0ywiVy3ZtmYpKAPL9mHd58mxNYaDvQz7J6fzGgw9SUzLzLhVBBV7o6g2lUb5
AY+tNU7QsG/gAklJhxYiepnYIURGpwc78bF5IUpxoqFo+YawXeQTACazABl2HiVRRtoevK0g5ZO0
EZBCmCEvVkrgxgI+lL9GiDP0MyOTFKzgRyued7BAV3Rd1RzFCiPhkYjl1CeSzTm7l9nXjgIl5/f7
ccekUN8VjC077eLHVAzXSWNeQaxHNOm5cwrGYpYmf202sVjwXHBx9FMkr/KrGeLLG2qouwKO6tH9
t6JbmQh6lys4jva9Gaqj0sz4/OjUpW4KZdMVRBbSmKdP78ClZ3HvmL6SsM5jXGGpyqf/K9ulApob
OkYvcjAKg+vIgvuJuh5wSAFQ58MYj2rq0D0Ot5gOVW+PB58NrfPnij4FwJHoq9cjyzmQsJ9wlmPD
LTgeZew+KAqKW9REAvksbuZFVq54MDnR2OmBmPlQ3aEQsMRNsDxlgynLpyCAhxbilemeK8vmd55p
znG0pq54A90dpu3SpfFBuYH5jeGcOVk2eHB8Rm3mmmYwXwiXjHhEM1m60R+s1A/Oi0yV8VzuyFr/
ivfzlVzsOc7fVjGXd/hFvAWRI0EV/OMj5b7tfTisgg1yPtPLf2/bb1KQimEbfHs6du7eW9yKqC0K
38jfwAlTmopupI6j19bTzSvUft+ACvjEODLVf4vcLlHRW7VVQ6+/5GBAXyv3D988seLMHlu7nQM1
KtLScGwOhGD/eCTOt6NiaGfrfN7bv/bws48IFLOsX3BnPqQZ8ZkcxUNrmc/yZJc5uaFxhspVyc2N
tggje9+2kIVZUoNFL9Yd+T5hYORPLhY4OWh3zEJpnGbkrUqpUeTpV2xgWCJs72exEOiklHRnNRUf
WUxX/kbtk9Fo2Ic6J5K7B+HPVDpz+Gf7dj0HjnETXXBuUKeTFx5S2/129CRYzIzyQznxuwOPxZI8
4cSVP7tCrv0rUyOEO0hYP3NWDezbPqzKGKZ1HHrmgIQ7+3pkKsGwk0mKRi7qG7buNHzcGGZtIDjU
Hc4y3U6cGIS+Vk0uFYwXLEe4IK+nxflzDQ2fO0x8iYPa5c/YYuoW1J2CvkrDLQWzLVOzCh2zrVtj
bIZbW7wt7XKjrGmyOS2SUL/ArgZ8q37rpZHynRsVnAUddiGNveF2C+2UVhKu5HAt5WaehbZ9CzxU
X0m640Csf0fpAI8urLtPmOTlOjXlqD5TjC1BR1Yr3GXoeeEUflkVZhDeYfW9cVTex9kt7cDfmgKQ
rgLnritBqRTlVQie78cR0oOhJhlDANf+0VQBhQhD6gRguDe/vsDJs+rjKYuN6PD1Wn/gewDynDT5
O6rvr4bcmuti50mtpMdNAHWirfjryy24qCJt9+2ZY8aXREhjtuIT1y+YN9RDLrxDhxxIb/Hgw5BS
l8x5dCkaTSKva4k/iCKSeeKKy9jfqpPyZbXVCsLXRuHga3zV+Nu1IFCJ07pipCmXSi0FnwE2G6a6
zELPU1Ds5gaKC8uNFqXX6qm6JZQNqURabCeAbOu58A2bvraHtFCX0iQQ50ly3+3UcUcZiaGxMfDa
GWCLS4JKHA18zE73l9AK4B3PdZ8C8uBgo7/jXOvtTEnRRyn/s3w1pou1ehqXIGRAvetLT/O2Z1eg
K7CKdmdg24Fpe42ZlphExrlEPamq0jA6ou2CsaupjXBzKwv8MjzdXYm/qzPAngVxy392pwxuy1JX
hr6ul1dSXoPEToiczJyct1IErM0pUWfUXVjSsALCD/jUaz28hoOk7OcN1gJWeJdmu+zMkb/ad/qS
kdicog3x/P7dY1Bky0ETv2zI+V8f2yl/O8xLxGqGT7Kx4lCWWaJ8f93cwVPVL+Mu07kG71kmMkjI
wo1sTVEvPuD4vM6l4hmHhjJ2jkZTHJMn/I97jtifawlMoQTUnY/5aPZkeuGlTHGhhgvncBxTU6VI
+Kz+cBlbMU93usc0h1vwZ80IfryKRJCRqFSkTXqPVaWQwgZ+tNQtI2craLhWN30R+78EovFPAjqI
Lz45dDdPo6NWdUIJXC3gOtTBfCS6vnENiXjVX09fWFI++En8WCL7NuTdkrSBvfXMopGc3EaPEXm3
VsaB1LZbNTZw43HYU149/sH1qitFaxshae/jlmoIoVhZC+W4Q466mWZl/dxZ6PN/et5FjvfYG39T
P6mfMOTfywZKWdwQI8nc/Yv0rBX2hgzpSEYofKTllnXOd3/C1JRFRylyWx8+J3wiuErZ7KsTdwhb
Zebl5n9jdbbcXilOQnrMdgQhQn7+XLfftmrVCJyWg7dO9Fv5XLy3/E1Rf7JB57FNPzJWGR8Edxlf
eWJpwiJpWVHwFCYTYSCAV8eyOJxyWc1iVI50Y31tV/e1jaNiK31ASmrjH2W4aHEkkL5S78GlQjTQ
g3BYLE8EfhwZ1fjleyg0AdSf47mquK8JW8XH+N6bRe1e5MgGlNd4Iqy9WGKSlFZZ2rMp5dyJmxfW
85iQAjREjBWX/2PTYzm8vk/xHiob37DWAgk+nkgasvtlvtsb7v6l6fHJy06EyKP/pmUkpZfCnYnk
KCmhYNKnI2jkGA2OTWYsnBQMC2Octm7GQacTCyBLkkKdR62GpJRjC143NCHQrSvzL6rF+88LQdWw
Xy5BzQsNJEBmgvOqY3jM0r8Ar+TlSvOG2g7+D2wtUNB/+gHTkeim+wIkiz69Q7A1xbBSjjG97djv
pVlFw/v2ETq0FhOIIAztLLZr2Qf6zF0WjCuTgoIXF+YC1HMKAtkrnNAHcl6fFIDqCaRg4L7epuS4
H1cFdxtLHaASExHkQLqs6T7GvgM2SmCbl38kigE5hbkAtvtOTmOYgSdg5k7Z1ijY2/CYkvlsJulF
xKQcVZKQiDk2rMP+9O2gb10tUPKnifGKDcizMiFzr3jTScctpGgnxg5gHQxelzEUZKhKx7bmVttg
r6ajQrBVqvM61HHsabySY8qqsOfY/rTa5jXDZ5iDZI72P5iuCI8YaaHIVwalUBe6SOusHiYBBVqo
0wria3p/67D8n83kYKJWEkNrXxusGIYwCR74IbdbKbH4G8m+8Kzq9IltBPxLYb9mjnAYWYyudmrN
m8+97l69TRSyp7hwuPukjSlUql7NrNIoZOvPwbKRG1e2Ag8IV5ltXE0Ll4G9gAvlhiX5ZAHW/x9O
KP28ipNuZkvoeZAceofessmLEZ3NrH1Z8AsS92EfhSYcu4dwQ2bwTrEocHrZ4dardMP4KM3p6BEI
ik7oaOQPoK5/NQ5IrozpBLjiv8N9By1vb55TMUMpXL0hftBL/bELO3vM0jk80bHDugcyoXbELYI2
k+UVp8A4N0DH9+blIoTxJZwklOWGiEUP06HU7kzHtXeQB1VnD4ibQfEe1eOeD/ndyEVkARDuGrn3
geKbBtn0WapS1gXDF7NVqsHTxWEBp37i7bSx71edYlnO7adNds2gJ0fRcIbzAdX268YVS2JGRP01
SItwtYG0m6ob4SY1rQV9DISzbjIR9Q72k/Eps/BygbtF8ZkJLtMj8mx2dyq+HDs1kGvWOS81A4WR
rmBI5Yqz5qSug3QTCs86DSD62I3f+Sdj/dJmvwjNFZxYS+FJ2v2rdcTaRjSX3OfbAm//IkDnuHeJ
OFrUJzcMNmT4n5VWsero3zcbjT0TlBRm5B/EwLI9u6AhffMD+Zx1cGTtsFh0DuynK7eylbV4jxXq
CEm0teNj4NEdPb9emwgKOvWK12+cZPe44ZJibNyffsVHKN+zimoggK04RRuWP7Drbg9Por+xX2md
PG5Kf3f6aXjRjg2Be3yZDjB3QJnPeLigWrztBFroMLEBMQoh7ykCOGhxmVgm5c/QhVOoqvtkIgqp
9b7KgIQRmGRGjfnieTcdQ/lDaTYx8L3dyDuXfaYqqISz6q3XZ5ywbBJuI1fWJTioWzGaf3SvdC1r
QEd2F8zgMfKs6dSjW8OJ33R5huWo4eMaCLRtWoE93M3YMlyyXG/SICSB0RjjhNpMM8GoQ5JLFNb5
NRibpCs6kpIbApCe1rlXoTIg1CMot5hlN4Sfxktq3w6c0hNlxs4w/D7o3UnKbCqiIhhVbx4vnSbx
aKNVaYFXS9HGr5oG86bsiFcYQUvAS+tNawFG6V69JYoZpIU457haiVA70c4yLRcvq88585UrqV2t
Z/mq6mlt9zAkjl/bnqijhwPErd5DDdGMEnzsXENzdjWzS5OH6cMxna0oNfzRUI9FUXpaNgNexUcC
V+XtPZDNXECYng3Nsri+Xoaqn20zukCz4bwPpYXlpT6d6lTAv3bIYU9O8oHRbEBjGcbvGlWrIvax
97RBtez24zXkLOdrmXFsi8nAlFF04RYBWXR8fRp0rufJmYFao61UhjIwbKO1DFHQvM5D2hCIQEwg
g86BiJO4c4qrOkOAi3+K1I155HwQdPL4vwzPZaaihXLa41V1xOlOIfwr9WrTqazPV7B+cO6iSxUh
3VO9K533Q+TGX7vkqB2FQDxHNS6MvzAgpx3Hep0tlLKVVj7qP2Mlk2F4zX6cInfxSAL6CKaCDOXC
Ekg2JDqI4CNxTFe2ixo6dxfffIeOLAQIcVLzBt3bQ6ztayOJgenbhgLbYSMCj7HOxW/YTZDbtg+S
KGX5PSxkuhniPiEoQJpG02mL/HR19EdAetmaKkbdxlg8u5fyPoNWce3lHeb6JU74Ib2yArZE0tjc
ruCvwLiND9OlULWZJDClkmUFmgiL5GK7eHs7DSD7kx1dd1LldUKdLCFbbkWSbnON04lYMBpGmhb4
KnwWbahbqVdxmYSL8K7jCn84EcIuLt2BoW8m+fAKW1HGKwAtfpwbiFhAz+jMuJ0xi/tJ40jTWlJm
PnQsM0D2yl2eFg+4a89zGzVrchAuTUESR9RkD0S6wYd+whu9xxk9anz6jwGrijt5fPdcJPO/gOP3
l5hGj0D3Z10r1IA6hru9/Rh/CeQkwudDMToWM0IAGw5pLLV0ZuLg7uwxWTw4V2QD8TtYC6j+RD7q
vu+nkKKdkH07yUm9n4fYfkc2Nhzcs8bKk7mSbbpohUZktwsPIeLRmMQJIDa56o1Fb9FK+0VIiNUD
iYTUfTVD1HFn9mZXyludZm0Dvz7oENg/PvkDPFOocxlg5GY6KCEDDEf83YC6U1z39z1FU2VoLY7x
6M8miiDp35njk63gaTA27StYYjlVQfAY3Qn/PuX8gJ65ZsLJ/3/mZZLy+pAMP084hvbytgbo9IzC
hAitagrbCjxCMMTMMVBpmyxCOtndqFfOJeI2CKQpmrESu/zl8lpt1Pk94E2GqFq0JtStlo5KWjKl
UphdpT0DdkMtN1mfd6CCoC5deqHRV2C3ZEBK+0g9Kc0Bmo7htolTVb5Eg9AYPhdNCIZ8+5QHzksK
76j3ZsEL/3NXURgmsKaApG1CXyy2l3a9xbCGrOr/1bP6A3jMp0eMl1VHZEMVlhEfdAZ+lE1jXX5o
V/Um735At5dkxwc97xhrA2kp3FXjoAdzasntc73jIZtFh8dJssXV46G7E1tb6CFgfqU7AKPyQxzB
+MtociWN4RmskuTYX2l+4O1/T4tLk/8PPVuaFgEHGqZmSS0keNl8SqCcpviAae8u3oj2BSIUJ+vE
C4XVYASwXMrjFB3E4Be0r/EikH/V2OJgx/I5LyBDkXrJpq4hAk8vQOwjzn9pXeHpc8f8EfgOFkxx
CYniHyxemhCdcJ8QrF6Qx2vKn8L4YjM64jNPduxTLyH02vQ0j/wDceYlJVGvIQm0urqRMyXpTVMp
OVonZOiV1KpiOrKluKqtT1hkYAY1n3wPfyur8XMxUbYlHWfwmgSEzm2C6RGGyeAaiosc0tsCeGL1
0QXrHM8BxMKKHNecTJ2EwFjwIBHkmqhoL9EeDnUn35WSRDbRktTZ14fm8cuR9gE9VUOzNxltq1Q7
pozD9tOdt/bobrn+Iibhj8Ov82KUJd9YJJ/MxwRDoxc2mbtzLmOu7sBmvgJf25G7ZQ+OudKpN9PR
oIZRDMWqaYDBHyNkYyNSK7Ae0iVYbTtuWqgBgzxfx0Cs0BeRT1juQa9xXvy54VemJHbXVmB1tOAN
K8S7DfQwbq11dQdppn98FVFqpeutJgk0QY+ax4haN3Ch3MPfsBDTDrEUYbOV8fyYX3n35CUweV2Q
wBcbUQvNhBd1Dx94jOIbzOygcCg1ECfBtUQY70U8U6tW3cJ++H5klai/pcM1SIQlG1L1lAL9N+c+
wRH9+rvRh86HX1cOuYj5mSFo+5A/HWygQMQVD7GEsTbJhpD28pqjrNQo1mSKzhPTw+Vi8pkaEIlE
yasGx0wyseAb9u5cWDNIQuaxnMHVzp+AxYNkVIuGs8p92jjvjCK/jDsCbHXVtBEwjLwJ/dOLm/9R
kMIpKrBmmxBOE8bIGCMu6/q4g00ERJ68bSiZC2lJvk6j+napPS+yo+LZKNr0lRHrTzpDPG/GkTIt
pb6haCnsH/5JDd08ElMSIZv75TEJUGV7PUOuCDiLxs2TWWcNjqJzNMfU5J927kVFzkmQ2O3UfdHG
xhkvzWo7R3FrR8BGbBJl34B+Xw10hAM5N/4/3Mc4PtPHPf0s8j1toL0z0U6nNA2FCI4zv7BvAkEA
S8i/zA+YJ0hXYVTWWH4FYNG5wDx8iPbp/YyaBNYe83sVQbzKLQzHgS/AGjPg66VSBtQo5o8fpZ4J
N7kRw7JcCx/bb6C7DLXvraCKgevg45drHDpqkxhdBeBS6kMi8jcuSMRbnY6h1+XeUYOOw9lvZ2WB
PLxzsLIUhf9YrzvmdTR4kLY4jzAsne1SZ7VILpTrxb323hvT+pNw7bEhJePMkfIkUuaAfd/qfJZ/
IU2gzXtmMx/XG/S8inzLS/4KKdvzrqyhcY1iXncNuEDm47IuiJXcTpbzrna0rjOMMSYUBcjybxvV
B9W1lj46dCmOxEKRQBexic6cHftDGFfQFIgvPh5Kh9l24iyhDSLVu6Tn6dp3IdjavgcVE7NGShEE
pLaTAnIwmvVMwt75Z8eDtegGqfxP9pF2NhX9QEBpByd3yMii6rwSXeadp0Jx4jheSV5lcTZFPaOY
JXHc1Yfff+A8y8GfH295+bz2tcfS2yG9RIEG94vNcQxPoF/RM9m3g49mUasF2dcFGBKuNws+kmnj
7Pn7hsb7WdBtrLN9kQ+qSngQGP4XhmJBbSKp9wvruJ3sljd7O8HXvykvMWfngjjgtkjUOyG4otcU
YdS9jdgeW5uiGFsEgju6aCPt3n4Gnlyv4agEEwmBwvLQhJYJWWOi/09H4ExCjTxiuyTegkrMs9s8
qHbt6X4rctnX/0owXiAlYSUM0+LEurE55HIZjhLZz/LzqQ1N3A5dQcE6rBpVl2GkmZEVBpLlqSVD
Ard4nmCII5zwrRIxJkNviX+FbUHb9MPUxz7ZjrbgyApNm3uZUfJymZ7d87waEnU/epIukzuI0yMb
DBpTBrzsO0OFSIsrAVeKlxgrFezgLxuXphlinaw8xwhyasNeX0w4jXaY9wquBL5MCh/K4AVHuTMQ
2yarSSwtfQXc8MRngUfhRcLzc/98WkDAclKCNt6igR3j44KUwp3M12z3g5EjWXQSNWrfeJ3LPBN3
APMyZwWU5j9Voy1M0Zz1fV9YgvEg7f9nybk2s4QMGq31fOF1pIs2XFJ8nkT+1eYbRRJhd33MCdg9
r/p0jLAaPaxbvll2thT1Qr58u8YsurY1MxGeWLqX3Iegv9FKiszAhHqqsFkyEazOkbUC8TJp+9ct
xph/EITZew2sQ1iFUcO6TlUWl2+T75oQScABHbqXO/e4ECguxpGiFyvdgJcpbKIobP2oENeVFkdh
uJfPXB2B2Svho+si9WqR1ytRDjyYv4/7ZqtXbbC+pKlZOObMXP8mTlPRUpQ02SzofOOtvQJ4yww7
Ax1Qhf/Dg5HyzfnQcq8nwQYS0ykUitOjbbEi+D9rZ39i3AC4khw2xGxKNDRDDXekO+DeowtuIEs2
FpD2qYn/ohyeNZuEyCTH9zZsbGkapwWBFHenjj8p69kQOLOl/ltxHqeeyQO9c2eI8mTjBllGNWAE
bPr3RfqgQV9HpSldRdlS+PKnU3cyMvVPR3HmQVpxqHAy8f2bjNIlmoTb+d6vfjBDRFn3bxeq9jWG
lqES7UpX0vIj9bse+/jymga9W5mdRXGe/rbWBgaixCimdQU0lW1SGJHZqaqHgCGEuLFJXZ5bDoLO
hJ0lxpxmNT55Einw7d9PIzxps4+FnZOpmLPaH6NSm3nhypkHxZ1p9LvL/zor9IXnTJfDNxDTm2E+
RRlV9Tri5xGaKNUjeNv/U9vKAfply8eYaF3uXbVZQbVeJamVca1oER7Xev+cCs5V7paYJcSDOp5v
LApQIW3/GA3pnOoO26diL/i4h2Lfd83xU/uteSKwXw8VZm7BD6y60ztgExzXgHTBzHuxseP3PmEB
+g0gj4Lv26GHXhb48kpATCLJt0VFpDPWsCTVRt7m5MQw9RhT9UrccPpMoVsbeCkACpEY+GyXBYaR
BBRkpEx3qnKDsYDRvw1JEX9VksT5jpWHY0Xq1qfgpnNkrVLCq2pO9jDdSKODWVXuvA3QVIHfj86/
ao8bP1Xw/fNixg0BrBQ52tMuFIyuGFkyvNGofTFGbk1Ob1EJazVX1MAs5rvDA4SgJlZjgmevpm2a
z330yshjemtfyQJVT3K4MZT+FdlEk8FAW1Aa8268VtE8ne9d58TQUXXsN/GG40ugzOlTOz76PuEv
Ucb38aW+r5y27PKQ86Z2NKr8wTgKxOkZSZ0nnsdGZPcq3/ekcACFFqCk7bBbVwVt+tsXCCEq033u
rUekNZjIBnGjTjrFjVwm77UAe5DZw6iRX/WZmPlo4pXnxBW3qxcikHfJ62gftwJtk+XT7RVyKFDX
LWkIChf7ZWkC45RGKA8AdxGAZJu4xT3zR/ukTgKeFUnmqzKmmwqsiZSq2fCc6ZlE0ls2Xo8rh+HT
h7ap+972i9392HeAKASRBSWcb+l9DqqzaBjfopb99dpFX+Qk1oQyiaPQDued6EHcD0tNL5FtktyZ
q2DqCATjWzlkzmzMIvb7Eztw2D6ClLVfV4gbyOnWBmXQEeZBMNaRpp1TBzG9B7nc7KhGSwj6tRwj
CRLx6CnHQPq0PB7wiCvkf4L6rm87yIhJaHz0zrIyPhjXcGI2u+JpW4KpgdE3KSZMUjTzpINZ8yvF
9oBSQV0ATZNlZCkarIbh0qxm1EOU6yOlb/ZTOl1tYXRQraeVJH+2pT3gD0EVfhDrwRBMGqRTZxGO
vYzzs91YVy0dtfuYJSNo1QABxBm4L1QMNYEqjQ0dlPNOROJ3wj7M7A10uZEjHekld4s6ZpRAyzza
7zhDuBrTDQtT+N6YRn5xiYTFwXNMaHRgK7jBCcXMeQZCT3tgQ4KxlKnejGss2V4k9W6SXUroS7wi
mpxNBcxNH9pVkJX/zitaFCrYfGKM3NwHh9KRxoOu6OZHd4LzbLAnJSxRDkZCffZ7Tq2Znz5EAtxK
xkqvGwiP4qY6bwSmFiufoFwVUBBFCgk3XTUvkUU4Y5EwYW15PxMgaBbWmE2PTgFwgi+/Nrz9Z7Tc
Qq185Bif1LJ8vNNznng0QDiRCDsj1I1bgWkAFL5/VZUxnArh3LRewMvS5blMANrriw97YBatNBeO
lPxJ96rtV6825xMkyqzXi3xTlIo1ob6rVHyU2972rCdlwVXvC00LkdIIzl5tRIfXynZHYkGOkvf2
T8S+7iX831QtpF8VOZDfMhS7YLcs0oSxvRamhoVB9FvNKJO935LusQxwN1AeQjJo0O19SQ1tCL9s
MU3/6kNde0ANEDqVQEpD4nLHfK4NPlr1EdlKNLECAtnzkZzBe5m06qUABl3pShPWEFNCIG3onLF5
/DABmMtPcXqVM6BAVkzuLQDX6hMKHgNUrvOvA5dp5t0oRlvGzZtvd3W1/9XFq3B6q9my4PE8uiBY
reVUropSXvtRxrPuK8IK29K4YH9jwV9x4VbmUXnN4yXiBPPdsVGv0epPmVlyFKLDttbR91TwgMQm
qI46VZTxzC25wFWNh0qelUNlMvHXFkEtyflR3aioloS7UE9HSwVZUyvIGcPCkmne2xkxtj5sKZv3
V/H3UPQ17EdlWYFUdMukLkFhXuMO6xZgsfTS1DYi+X0aWkzlwVQqhLV326Bf1Ygj2FE32rjAA+ON
SIJi97ivdZqSViuvOKAkArlwOYgiYypzMhixjj20XqufMlqkGTzqgSAYphBKPXYOTnBoBEAvPIpb
4wicxi5DXWTR1X3ZVTE2xo5XknPgpinjiJWY+8wIAQicNCdsW1z3OqTOGDHR4xQVjvAE1lNPdK3O
RgL5kOeRe7K5q+n+/LmTGmQOMgMlQyw5Qz98geiZxXE0m/vXeqUlyUHOupI9zNYjyGIecW6cFI+v
og3+sM7Ry92/Z5zTJ79yJt9PbNh60TBQJEw2QKRGJdQgkdejhQxSJK8gezhlMnvCHH8VQ0MOgF0A
xfQO7PNB0GM0ekL8uhcsbGecHUsW1yiJa871IrgUiIM4Bc+Xrc/+T8CJWOaCh9KLDuW8Vg7zTLt0
/h/8kXOe2bqoeX33zvxfsURvGTKK9e/OyOBLkPaDydepbrW93MlgbK81DqVVQmjUrMQKIyRIA/+a
27JWZSYVMSqk7ODv3vyb1bSrRGwY6OHA6kKtxb5fu4qqii+NcW28bYsXls9bd6aCIpy8M7/HHTWu
zvCHswCzHdmLuXO5g56tfbaBgs1NbqsQrXzLFCmiDaU1I00oBRVVvK7iCjvX6P49vXqSqTlg+hAJ
0MKmeYuI1WEDrMbjrcnPahu1kiCjXTlMimNsr4pouBhIV6ahr5E9uQ4dhZegMTMbvYsO1boochJG
+Vzp5HcVKErAKfY4c2mGlQdQsUz/3ktxmYi9XV5pNBghK5ZEmJ+FK/BIPxYNbZq62fuo7QMBSUlB
ZafWD2jXOYRi3nsZFH0SnYJb7LfEUW4A+utUpc4+gz6MKEJsw4RpVCXzjdwOZFrYzI9nA5mh3l3Z
W6ZF5tcLw2iNM1J+melHwchFnUGbMqFS2S7SsskmJ4IYXjrDuwWg2w8AHj0OLQOATAV3MbJLyKE/
yF0RoO5qKSEhWfX2mzTDnYytcFmz2cC3WdDnzvo+84kJ+Nl+JGRRQdB51YVgRuiPJKlxLgC7/bHQ
PT4IidZ43sgMDt0XUhq8Oy37Re0Grk3BTo1HiI7bFigV27J5ThO5OII2R92i2WgB/1sEOADg5sBc
Elxjs7p2zXomiiG+G61CvomU0S26U0FUN3tW7ZFzy5Q1fJuNNKJ5a2x6hJMVD/uq+XUEzmZ0jt2L
/7am03U3xl7OSB+1BkNHw8ALncXJGgHn+482TpxgPiKz8+kDBgzj5Tp1/rHktW8JgxqyyRo4ya+A
1Qo3UXX66tgp0+sdTdyhPE15cYdFAD0ra2J11DwQRrGNtbqRmVY0wn8EKtDTZbPiK/LInyXzeQZD
zpaqdebruRMLNcWUtqJS9EWUuUijNdOqOeY+/Lz2s7pwfyNN0fp1UEy1gDd8Oc4A45ukJeBcvMDO
b1EwSW3L3pPknuVhs8AyOr+zBVLmqGZLWN9E26FRO6o5lV424/VuQBrHpkS+TIEvBHSzyKka+FnR
ufEVIpkD/PLqK/PUz38XxR4t3AU1JkuzmvOPFI0sNbSl7cUmmqX+ZZNrzvrcwrjo0r6VWXH3IGU0
ifavteX1SnPK7tkme76zZGYwPUDdDOWNELrIe3F2xNDXZRNel89VrScYUdLz6EIkYXtaJnqdwMM3
3zK4zl+NAJfKrilKU89r1fuDmwchs0P7ySm2xlxCBL5/Jf1qip7qDlj6ZMGtvrMwUomA/fxSezqo
H9Ae3nEziwZ2n+W6g6SzArYoiUJ+Wy3nbLGp0RW5/QYIgEbyhjX6AyAAfzpBFl1zgWQvMGRyc0u+
eVkw7CX2TUwmNpkPcpzurSCPbznlT7cIkrvjjs7HV1uCCpNavzChsmbkx7+gNn9kpgi112HTraG4
cZHyCdCu/zd6pdmSDDSzIwkyMi7UXD1+0U3O0KwlIz39Ysr8oGSxKA41tArIgW9aqhF21pL01zk9
WhBUT/qLaSslWuYl+SrZ9w6EhxNOFqWoLAyib7WWJMiDjioKrPixEY0lCqG3ObX4Vabz6oA5ZRk7
Gu389pdLVSALg/t95R2fJmHw1hlYUirZztovkAM05KZ3yOKJnK8qXZs3+YwFkz/Zwv4bhELjt0CQ
BnnSalBCBaTb+eGdr5ySymkOVJcw9j2TGO6xfiSfVM/idoIEsGq9r7WcSERZfQOGuffphpN3WyF4
DM4J6HPYt6vKIrrJiMCGZTqG4m43gy3OtWboEiOhu5gQX5H7DgfTxOS3Y+2nwj0zfdmQBnk9E+Il
0FoqKhmeb4eYoVznZb8MX5lBY4Dpt1yw+rT2e6vvYaO/Kdv7vr+d2zBXYpK/Z2jUFUC0luZK4z7Z
3EgpEidi3AcFkJ6BBjXe0WZ0szkL8bGot6KMhBMvCasmtv4Dll781HWla7OQZPE2JqHDf17jRdbs
YZq7PVMOqj1XHR8XbuwG7i8VuS7pCjrmpwlUdAVoALfkongVt8yJQY3AFHGPETbs4ckstM5KyfKk
wHiczXH2h+czyyz//15g6V+LELgQBLtnMlqtiAPSjQGCYPBAPW11rUCDlnsaKtWaBPQHOwO1yDnQ
/LdC/LjyzaZlGpuLCmzsJpzvcV0POIrfUq4ncmaza2LSfAOJ0cLjN6l0wPzV+5fwVWteITfPCcjX
hYt6KhQnslJjyLrLToHQFN2ULBQNbXXDWOm5XO8CfPM5PT2bdehF1ux9brG/SJ8JBXYtYG2wIwWf
slpk9/2WTlkqy09MF65XrI6l/zyuKtbxBPPsaR7Zt6wALBQ5z8ln3my96KSr0YjkuGdmOKDLDeO5
p8Tgv1VUOXiFKOdsn4kEFSWzHNYF9HgSIs5BJaq8SA0ymO77snrMCYIx76y9LT93Vx0k4q8uathc
HJBa2k6Jk2IU4YJRpzXYhB85XfnkiGT2s2CzCnuGHqzVz/SwySgbbznTmoZZ0KbYgh4YA7fa5mdw
0VqDTnHbw4FOnUudqz8udgbSiemVnhx64gP/2XDzC1ExyiXwQut0H45jQ7458aNhW1su2DP1MKrM
H0b0Sn7CLMq6IOL/XFESz5GGRam/QKI68pBNO20tr8m5nTYc6lA3ZzT2audfGinF05eIUWLKWkI4
yjmHZmQpviG2L0wJVcwD80DIqMF1RIR+J4j1cGOTH5FjrzMj2WehJfPNj8/xZvhRvcWMnpmB6VwZ
A1Gcq4RRWA4vC6h9n5Jgr6NxJN60rckb5nYpFrhmqqREp1zB+oIXCCqV4DbaQEf8cStsfreEP9Hu
DQu2RjR/bgTqVXSBS1K1gP/JJag75Nsrqp7DYOSDd9VoUua2tj+sctJ2nJXFDU03awKAMMi6irQT
pq11Ns09y69P03Y0BzKcKCba91hApK3RsbcLi3jeUDUJAFqm2ZapmEyrgt6uCqndkIJ2tmE8WmIA
Ytmwuj18nFKEX1759e6FfTu3ZuhB31MrN+7TFt3pf4fKf4GEfPVwOsOhhirH1A2WfsStfNVg0zmj
hjLiorFvQpGZaX1JFA6mU66vHB5j0qoSE3Q3y/iLhKNKo2D0y8jkBiSAGUC3xcVamgEPF0NLqaeH
+eg2frDBDNMTrONyJu+9DmDbZWDi98WuEeYWh5KPXwRVDsTHTOw6OEmZI+xiG60eaEo1HW7qsAXA
cZVRGFZU1oSVtQbCLBlc9C1yFDeyXZyRl1ze3HOPD79/PzT/46Wck0rzKT8xoZHa/gKja8tbV0B+
7YxhICjweq6MxUTHZbvsQiUk3rnMILLbWNrvGof0aesXaeUw3htfg8o+SMfbnnwUPm8xXRBKdQo3
3sZgxX3UEtAD0AZPg0zhq5CV/xpJjGSixa4hkYP3xq+J4MGet2VSF9dVOWvVuMVsx/AsJmkPntX5
5AwjIi34eIP9ry8V8dF03qv9VbA+fVyoSQstO6Df6/GvBWz4aBmfPnCT6UkXMLdVmOGT4XyJFC0F
bBVa7pVOgEhZ7lj/8f4tbCy/RibqLD1RHKm5z9ix+lJdPyvtukp6J6Rjr4X7/ldEsPiA1XK+Dqlp
VyNDzjalevHvmRTdo13V0khre5zyERHuab/AS1VqWdn0cvJn3ifVvUlZre6g+RAaX1F31mrojCLZ
+9XFz/rZoofPQUwBf5KTMW+m7UVoG28KvRELhqJro+Pq69/xP/GTrJURp9K2yWXr5WobPTdYdt2L
NGZ+L8XO+xcKUWoLZchHFtk3sigWzPm0O+2xAzz6jLgeW4ImaY3nTVsJ+f8mBXrJfNzQTDvSxq2X
NbjttwRIIRm87ndDY9VU2LYgkQRm4TjW6/I/wAkXL8aCqyJ7YFOIpijXSvK7CKeCfQTUbdwapdyk
5gJ75gk85bxys5qy8lFQ8uYgWeuZ3UWTTpzN2sO5ClGnyPvSh/o5urvk9tNeTc4ET16+YuGruG8v
91fpCPcc7LrhTzscQKpHfyMEiRemmy9qwkEWD2tRApeVAaSRevMoPQoiDfKF6ixAn+eMm3d5i3sI
/Rdm3/374gkkHBGoLMR7zT3rLy3unG/cEPRmrQm+CC6WtyaZDzVIFFdfn57KQ93KTCU5LLuGpkzu
S1WM2eO5/1FBpbnR+QZKzmGqVoep9S3fkDqpis8gsxm91LyZ91ZlBytGsmonU3PT7hx9lysTu+6p
boCHBTi6Qj3imUP6ZtP3lm3PARZcPN45wABWy3dBUpUc/BvJzxx04dQc5s7PfqBROr5aWGE8ew71
AJo1NIOixUhiGkUzH1n1ZY5lm8iXN+MGW+N+Sl3oy2QGkL46k8cH8oL0k4uYSL8MLBxOuYJKmx8s
cjdWei5/NmogzuGvD2GSkSX6VhEYL4ds3UXg3l5KXDCdQ6+OErkHALxFSt4uvdSyJpmHOxRgEoLl
X3ATcTgSDM+++9SV1lVSzia4wpHZBUbgt8qjP1iNX0J7Mm3KXLo2LTgMA5Y1GXq4+OUwTbpL8vgP
OUeLYbMmrMUNgwS9lRsaTEDBxSNJ6V/+yVq+xjU55Wg5MpL3OhM7YuLGEgXD9uG2e8yQ5gr0uP5J
7vluvPotgE3Y4Dl8ykIgBIopXYMJ405Rf+yBVbTOAowwWR94SoZzl23RPts/84LuCdLj2/ZFjwWa
D2cPyHrTQAANPLk6dnxqbjSWwbeci0QKtcCLNaW5n9c6W3wc///NVWL6a6ux9nvW46cvahKVj92a
zHtJf+h8/Qn7pL0fkmQwSntQhlDwx6+LHWSDNLkAzmhwjB6cheGJrPjhQ5h5n74MUpkInnbotxBN
12hTpB+/4qekTu3MwEI7drX+cAz96Ek3PLRULcxOR9b4JhEh0A2Hu228swPKNnZDyObhlM7IVVhU
xcrYXrw3zjAs81zhr/dwJWYJuxLGLXucAGgU9SlzQVdyHaIwiumrp1qaEbC4/lHQSyZnsqp0Gv/S
5/AwTXcmVjGvRZp4BWNrMQ7S3BNVTuB2GQe2KJ8ZZaNlflO8OYKP70WWbwylNUk5bYXMuOfWmYdV
lGdSlNgnMKMvVjMIZ2qT4EzoZsGT2BW8SXjUFVi8UScly8rP1xcESOB1mG4BZVPPnMo4q7YDn3Nq
xzJ90Wt5nBoGNixDL/jlt6IxfiH7V8hRwTMxDg9CVt/ozMBtughRy58erAo3LhqnLdTopS0lA/Qn
JvX9aEhajK9o6wHz9JGETSyzzocCGSn6fqMIVhwrjfijo3mCh8chDBZ0KB/u/x14S+CeN+0740VI
s/GV1aQBjvbBJqsSXGBTqlA9sEopfgQRiHMfdINs45vZ64kbKA0x+Y7dyZBnsPF6MeDUOJQshDgt
dv5D635uxkgnY+b/qbOiMfjOT7FGr2hhC87Rd6BssQEmxKvqX/9wuK/uEjEshPCZ3ZJJ1bL699hN
Cqtve7mXRr7LC9LWFPp9U+KMf2yIXurXuiR6E2h0NcXh4wQWWqtFun0vvwaTt7JJoj5UIh5OaN6o
3Tr7R5xIFr8JPXyK0othDmsEBEAI0ztq2iYHcVkV3tC+L+jrzY7QHP1WlU/VESXczfttorFSbZMi
2iZLDkI1mAgM+ErqFVk+a2WxhPqWQg/aWmbauIvDCc0sOI+yf490JlqoW6WRnaS5ejyeMZFKTyJV
N7Ti1miuhhTWzB2D3tl/cc9tkGQMhkFWA7auVZlkW5zTyVQ028ACdEadghyqZ1WQwmZhxrmFeT4c
akRqXoMoOGYCkVbAuuP5LPbTspESGjkBX5F8RnEigTLB4AXkZVeWSiScT0J/Zri+ti6krdH56bh1
KmE3WNjg6VWF0J0yoWh201B9aM9qZHOgeGSTre/ELXGFdHgn2TdNi7xpNM9hEsYsFCD+WIrs6MMn
jvVmBtLA2e1ghoRrHFFxGRdrgZ52zt2EpttuI6tODUIQyskVy0bLZkWx3YiXrSPE28WKosz+nppQ
7r65S53clk5u93FrYMzzI2AAiSu+o3EcdxcF3rQ+fgA0viztTszXCD5LI+pLYgtSP40PR6cOXg8P
fsnhg6uSCP7x45xtYEeuStx2OBoqwWLNJ146vpE+Ql4flUlJ1A///zLneZGbwj3y3edOK1lCxXHs
JwpyhNljceGNR49fyVjuOLKkCXvr/be9AuCQg3tZ6lfcYz9iEzJo9/Fw9ITiDXsT4cYfI/Vda6Qn
pjP95oYeFW/NAxZ3QnCSp6fqP8qYs0DWRks5ZYBAcv10MQEs9L/7KDSs5qMtAILT245aJrICZpRc
AMlUXNinMrpmAamEWs0a2zUCiJygJJMaqo1DoJSc/zikvsMi3u9xhBLQ5Z+xLbuTFeCWA9RcMCll
RKM1SiWdxmRmx/qPuo3amDss4QpiaO8jLwfEF+ZG6cuwasRT0MobT6KWXSXAfJPzlNvOiQnX+1kG
OoU9HX3y9SkX0M90z2R+t07taZNQmCRadV6ToBpVVz9o+ML6bQLHByCPGVPYzVn7rSIiMS5zRqXO
1bQYD+3Wfo8T3IzYOYBUHjgQQPG/l+3A26OVwyyFLg6VYPFhBIade3TV0qsuG6zwyKC9xNVaCo2s
HzYoPlBFGs4yKEWe+NWhTgdDQwAq14Xs0T7y2J/8+Ccwjc1b2W/QDhPctUTEMdZXt1XnAGA4lwwk
/dVD6LE5DqklDu5LgF8vpS5awnpYfWIPFENMyQegESkNlHnl3MSVX2ncOq+QZxWYHOcYAxtfnmiU
aNNcbgXbtTO2StF4jggzliODtGaRuJMuIyD9JW4VbgE5O+6FWu8UqPTT+9O8/AzGLp0NZ/BwkZnr
fprnzqU9lZAAPbx+u77wzq2ssQZybN6xGGK6rLFmVDLuSqR8CvUFbbo0sX0/WOYMPjpkGFjEkoNI
pvUj1UkMnX+cpmweBOFEBuANF8yUah8ubBVChXa+kcZko7AxlhdnGIlWJEziTKQuSH0edO7HpLnD
Zth9kE+3OfoE0USqONyEHeNtsQosLC4L5+LyL/2p1Hyt0m8LrPrd506Y6R0i7Yuu7zq5phOs1PxC
St/B3YED6mFcfP3hcADWwnxi7UtdgGctbwVLAxOToYFBD/ABkqrX9oPUmttDJgvhGGWy/+rRXq7a
NU6d2bZoNOo3Yo71zTeh+sYTV8ln0wRLWDzCuVgsweeiZkI1RYV5fw7dRmKoBTXir+AHos+bVYZ8
qV2RYiM/V4rqTVhHwD5+KhmzbeAdKmdBwaLPo/6EkyqyoEz80Lqz3x94817YBM5zBD1THrVKj0S1
YAWoRkoPwsK+mWC4sH4Hda2YDf2zr5S412MbwMMLn8mX4kXjXSCK54sPgxft5sSodJDM9A6zDpqF
2MN7sGm6Rxwrr8ZiYcySBWnJoEdxjAyipdPc8L8xAiAk/XavXwHz9aA3x4HuXorO+TZj78clKIhS
trbtQu/X8Zwjl8j5IMR2aucbqIm9KePRbHWkDIxFG87ulSAMokDCgSgylNGGlwvIY4/Jcs4/FWpF
NNWkhLXX1BehWvajadCsQ4P8QuMw102iVOdH/Mr9i1XyKiUihoS2ItNpzQiVz/3oZ+F361/r2g0i
PflY96Y927VY1bEbVc3HILOOTm4C5Zp5vEpJ9v/u9ySnPLUA0dlWC2jiVUQ7vQHp/jrmCfAazi/l
XNvUAdPhFBrtHB+YKxnSPBpwWh2V5kGn79eyGGU5Jp7SR9B+qlW2mCRQVfvSmBvtY7Dp7e7YHAch
/dNZE/p3VH9t0I7acf9ufI3ZHktp3pSeWsYYChZMEbQMkIVAWaIsUI7CG+nrF/PxxZ9/K/TXu1GY
1gtE/5jb3Iz7Pq8mr7VGu3wWyWKa1q/rrA700zA+Q1MAuqfPN6lyFDi3daE7S9NmQo++D/MiJ374
fn1X+bCrqG+W3vGJCS59H18p45RVLVypimvkTyiiWyL88RSRhoHn1cDJfVZMp9ax22xprFdNwXex
w+VDC6VSb7k3heuQnMwmfDMr//BBvdecFwelIMjY3QMJk7EZGpytiXYzXkgYY1oh55XLoOy+I+Rx
cMGjM/I3jaeBy+pu3Kz0NeiL2LEP7EFk8ryKp/gZ+wqhhw2h0M7kZgduRtqiqj5rT47k3YEJZghU
3cGPB37tPuuNxzE5l83pGhK0O07wy4fHK0nAR/1qP9178AJ4CwbjSHtqfPbj12YXmutHHtedKJPO
LNSTDlXp51PGEufMxGaJTrQEEumyxqOgyDohENVlqixozkbGQwQXGypOtKs7HyiyNRbp+kol0c/i
ULedKCHiReHOo0Qlq+WTLk8BOnVR+LBUmIGRwYMOVA7JbnpdEfueSykN2CH7bKvnYALvKkX0fSCG
kz70/OJ5uAQrFJtWfO8OsP6Cg+1h++zJHHGQk4W9Df9fb4spEZECNWvuXPeSYTj7PE6Pa9RMyx/s
2Eo1cn0DfZKZSkSzWnldznUe4/yk023RAptDgxnY3oODOT9r/8hnpdWbkPPEp8xc15/1U6ZnLoKn
ENT9s5V/eyIQrELY7aOAGU/aDoG1Uu6ZJOOYzcEYrd/QmueZ2vRp3r99TtVe9+tKslR1ihW/Sv9l
djap5aRG3EN4m9nayY/Nq5gnP5lXPGLoH1nhLeB+lruWnbu9ELtCQvpwdXIJjqZc7yVe9XFzSmnY
P9C2uDj8vIrOmHmBu+Lbr1CJRsOeHUenEncmvYSY6juvZg0TkiWG9tZeJ/JfVTUcPERMA5eBWS6c
hRTnYabZhGY1/H+/oxhfg0sEIwMsQsWzeKEGjnvPlzID+zRbrVLgkA/iPH6y6M3AFtu/BwAfCRRw
5QPnSTHrR1+2TgBxMylX15YDwJipNRpNQ9pd0c0eb0H++WBgorVh3SAlKB/HslF8qGxQF2fFNnty
khAw+vEtrpdBkpbiNb/PQfMdeKeayQ/Kk2rQfvj5sRRcdrVaXjBRGm0Z1Ju7p/gUVXD6ky3STOC/
VIX9lKEC4SvxqKPMTuF+eal/2o+IP5UJkV9Kl3HbG4E+isd9PiqGmD7jH1ZrNXtwti4haTOhOtFd
6jExdgguDLfR756gv4kXsW7nmyNPFcUj8DYaEFllw2HcZlXMGorV9kIb61i6G88QnO8Gcj+0mWb6
rHs6d5OUxox0LZ4msn05uWBPewX4NAdF88oGJCmPl5knYxEGr++ZPhd7lBqqK8bb6Aity0/n9mtq
towFnPRGKn+KC2/30vrrrGlx5LIGUwsE7TB22yyX9I2i5aY56cUR9WWRomV6fWpWZz27cUSA42IO
Vg3Ip3mu+34MWiBaoGY304SiO/JdIeTg2p1tEJT5XzwvwDcerRhNa7JHUhq5iqeKaOiSFHOgPhSa
+V0Le4/rLVx2d6DwyJ3stISJozLM3G2EgBis+5lVZN5feG5Om1SO2yLeIzblkzLSF5N9wJeVt3PF
Hmaa9TAhwPBcbCh0tcSETDdV4qKooU22x6VhT/FjFx4bdIouDhNPzGTVyikKP18t9XDHn80uaTvj
OeDsU+UzI3RdXRnzHHgmcyFLGz8jKPk4mdI/MDZaIzsToKFo8rLm41o2ofW6pCQkl1n9ugT8LD6N
Dq9kvL/v8dR9E8uxGvGxlZIfQUWm4v7SgMtbOcFYdkLwL6SSADb3KQ1E+ENfjxRL7dxhnNwPtBCh
hJ9K+ED5M4m6OwGGrCLlqEBYl8aFxVhMrLqwLHHPoGTCXoTjL6K/25Yaybh0TjgzOFUnlJXxNLZt
rZ3P91PODnRqdVdz3p5oLxB+r2L13O1b44vK2cbz6cZ9xufF716MPK/h83cMoznQEdFMExUZkmV5
z5jH5bowEID31bfby7Y2UkQ448B/prTRXG16zU/rlA+4jvIZZ4f4ipUXR7GeBv48UgYoOQaT4b8+
Cij2u4kDk9VdbolODcI0qFV005wtTe3rXDsZm01CaGu8bhuhFESBZIvo/H66QfY0lmnQfPvnKF5s
Pxt266Aa0xcntZ5oGuCnJAA/eQ07yIX8SoF9Sy8fX6M/4m0XHe4yJ8PQIE4+J2TkdTUUTqlQS+q2
JY7UwzWi3XRuiiqCz3of6vHbf5YhX5D/kfo76mZR0Z1UbLEEcwE21qmD16pbSX918WjaelN9L7X3
F/36lZWKVCAl+RM+m/BrPGlbHuFIK25EBFmhuJ0zurku6fq9zmRnabo0NX5uQCgYzmYUCrR7YIKb
byWzbxpLXPMEqg3WZH6tHylgcJh+e4vfveKXkDy/TCYwT0Uxez7UG26meDa1xgpaLLrLTURFGbEi
sfUnx15V/Cr7Vs5P9Z8UwXEadzv+bnjGBSUot52fmAaCU9k+K4q5FHe32VkTaUTzClfr4CU1s0N0
Rp1BOMvKDlYVVcACb+yxzLjmoS+/6WBvpL6uJm8sXxqZS6UP9jYZ9aX55uf7EpRaVcJXgDMiCtSg
1eIWOMQbkBsH+JuKNMoZUAbeJNsXaqQ42Ty2NxCaiIGz/ZEVwSiPeGL1XUUaH9/sSEKvdzjPomio
v6CqmweS0QK//Y0+Qmdoi9/5pJnxrLpitPNq7cM70wrhtD8+mhi/wg3aOenUrofYPjYSaqq8JoQG
W3XFNw9h6A3IiTnroqLwW3GTXUPwL2Erg4aHMnciV3u4EKvYJ9f8sbmTOvl4mhxTi7h3cIhLm59q
+zx20HI7mr2glfhgMnZoua3sdM8G6l1N5Cn/lxAMFNsTEGxzYXLPNrFLnlvhj3OoyKhs2LpFHeLz
kr6k2MVzh71b8AL8GebAPDyzTm88U3Xt1JXLqHtr2lTHQq+LIYFIFotY9XPwxwE5k01JTIsc2oIz
WSCd77BzmnofMGQO+pfzqrfK9TWAI7aW6gI8FtdFtPu6aawTL3By9c2JBFzvWawJbww/hUY2oTFC
eKu7sAYpu32wX3Kux/CxHGU6M2to2Cl8MycE7jqfqJqs6xnLMTjDvtBz+3hbYU3UEuA3o2x+ydfS
XaC/LjGVOa8HgJdKEHnKW9tvUkvevejZwQncOTHPIUwnRITpYZkq+pJWBq+vd47GUo8upIcJe2HK
pNZkAO8D9/d0/wVP/IaMxOxhDGVpL0q1bCQMQCOzS4HvB7YPqrCPbxkq0YSAJ36Aq8rjHdPy2b7X
ZmX1yLMekugyWaIXIRSOIuTztIHS8XwMX9pxaAycDTUcTvmGQSRvaPFYLF2eHJgkwx6T1tIAepxy
L9Lrt3XcvGvs5+LpjgLTccMcQBVdwDAbEihfNZdU6N0hHpleSyH1dgsH8RUyPrHwg0BB+/lnmnpq
+66FL4kvyIFLAJ9cfcHWBG+sswzTfy09yt7ASp5W0lwCK95GGatBJN73Rc3fVYf/2P81G2r9IyCs
Fpvua1Ai82c81c4hL8IbTL5oEs4AaKeRmVeQrAUtb9l+JVjMTOe+bnVI7WVEoBgUGGBojGafjKPc
PkU2VsrJjhIkb9qCLgbuPgVZHHyqQ8prkMI3/y+rTwoZS/NHEAuC2zM2vJKOIc9rNFrbIiAlDaMl
97VzC+EW506fRgbtXb7YSBkSuikH/T1g8pi1LZIRvz+lDRxqHPBRa3ZXqvOEAptUE5N4pMMfyEhJ
ytAPRM0FEZobtm7MNhd9r6fBVw/9ERWVj+926WGMKN+6gnNXMUaG54QEDQ/0lWmccPQIYrGLw4XH
sqUeRWcyFNb9VFlN1585mlrh0f+NG2rnuSes/FGCPn9EpCYgVli9nt53+ltpjwsmZJJW/5FWUF13
Ibxo5LbRwoVViZbqBuBr0bsgZuixzS+/IV3t9jBOfz/tkicyAQsveVH2R1uXx+G/jwXYw70LiuDo
c987JxJSE2zZTQU/VHjm4gcHXLy/d3kOg5Xfh2so1dsgjS+xXRur/Z4qg4ZUyF/SkRU2fgB2yfes
Ex6+VkQXMmVNiQ2Y+PQYy/dacoHkVDTSEZbQbHuisU5i7V8eHznkU29Fx/ONnh6QEAc4nhdDlfCO
pZ83z8Sw+/hI69xhU2dFiwFefnE7RyEqfvdhXH0pj3kFT1IXJpxsOzZroekypupzcb88Ib6HILQQ
i7jZCNFm7sVzYqHkRvHYSaq4VQG0xk1tFJG82dmqcy6S8YzQVFrsPHX87253QqLJta5imvAfHiC0
hh8tBOtkEOECczuBO5fMYQgoPDGtnHGmJJ433pw7EUnDDCp7luB5h2i02tdZFGMGOLQ7w0s51Nyz
94e7Uo1Ykr+sig8SmXNpgOZ9cnQkzMILqeXbdjsHXwq/pVjAS+K4+po/zNx9wQBTIhMAxK9wVwM8
WeYRK0uaEXXz9my9rF/nrLle2pvSZ+CiqZMqc8YLqdggwDfRB0S17XvAfmVimuU9abczPEXJCnyF
CFIMFImKDz7sIaQJzQdnXEcu9FKWG1gXT7cIwCT+PrpfHjiKjqU1WNwPstPCG10I3lQFluNr2B98
5Fde8db8sSOUXolDN5vcvh4WyqPeqe9k214BnrMOoOIyTy8asLyRxCceled8tOdazP3Fc+y7+U7S
VufRKrQpWrxVKi79dBgYXADHG7Ssq1Y0OqLIYu20FMmQzWqyrPvaO7pGMozzoNrPx6i0+L3lFX5y
vuvoLeQMIHyUJpsoP33alkJwfU6urSIOa6yOlG0t4JtH8Sfy0lmm4bvGBsCSyF1Ms1jBaDkPD1CE
GCM2Dv1wmJqrA60danZiaPI2unQ/Y6OetZMJf2gbIJEGDOUIVwcC+czxYdst7gslz8tcEdGMx7cS
VCVwSR6jRxEi+k2heXKopLPQHYaO3uWgidz/CYSyLqH14HXzVdaSMIjG4tkyW91EW+KzNqhRpYXc
Gc8ZSCgKqV0nv5VTZ/ApjxIcH6wwpf3TU8WyzfXRagUrMaENvuU5uIj9M1NsBTWHCKCB26KwWuFp
evvE89K4TgNgebESyzXEurh+gRsh0VaqvYnzpXyo7e+ukuHSCVWQm8l9XAdHoOQlHt1ret6fmvs0
IodFRsPBXtDilJncYKKiT+lR3cfmZJ0NrwGSVoucRYKIQbVcfWmtjuoHlYzrwem72sk6p1ZNQOlV
n+1il5L5MkBuyQikKEBr7tC0zT2qeRNnX191NWaUXMuadSRmbsbPyBeA3SuMUdHZQ3RGEC48C74J
MVLU6TSUMk2bQhl/vosh1TjTXHMPia7eQsmzH5XJVt3bV1VxVrtP3deHVM5IEu3C0ckaUKBBV+YG
WqPTRnP9lTVwaKO4JVR701XPMTtlplyzv6GjD7WHWBhwlDArkX5cFrgaQG2X2XlbHkv9j4rdaTsQ
nzBif3VoWSH++3TNaNI6/lEh5mey5sZ0PxNl6drZBlbBtWBKTN3S2NqgSDTxUb5FhS2Y9A098OAb
+qihY5gVLrIEMHWcaeNyv0yleEMInbReNm+Kfb2S+/BTzzaT/Rk/v3j8D13aP/yEgPkq9T4VEi0B
k7xqHqxPE1QuIgm7yPlj6QmtOCPGs+xrslJhMYXuuOsocZ4X0tGmzZVpdh0xFVE10lA1OFqURrH6
IbizwX9+ObZYF66/Wx5iaI9odEGijkt9QUbX2pyHB9OE4gIj+iwgSZ/c04+HF2unsFcAH9gNRi2x
f6enmCjcJYwszj2s/QN3si1J5GGDu5RmIt6WZ4JjLnVFFPhlEiYO69tTzD8X0IEbW8KfjidQ9P3G
uRLWMp413Ai4Kexwo1Z925T0N0NRyJWpaXF/Pb7RpipQCYmYSQ7JJ0bjzHZjkrTz/3VzPw+n5yph
nrNuPlwyXiVx+jm4dynXLlKRNfgto+oDzsPIrGqLrdP3GqnLuA8Kq3MeVrg5fwZKDZPTW3JemXFL
CToyCfOUXcCgR7sbN67BV/oorJJz5Za4C7M6G0Qs9sWeWWaCGmKs3i3/bjLSU0EBZMbT9miUO4pv
Q7qm11n/DeTUu7ZI5edutC7EcVnZBBdWwGUBEPoJWTNbiKWOZhaNvfSatQdXI4CWEAzXrr2pXHr2
H1wqGvo/3HgogYp6i6gj07Hd9KppNze+T4zQ79BSZ7rS7bjOKHG7VfByfC7rJmJQXp9OgwaTdpSB
gG/sTHS6FiGn/CCZh1VCspGLd4yKRZEv2KleP9BRO++I8hLSfc3jkLeCdTtvEbv91DRq54y/GoML
WJjNzQ9KgB6bwyIcuzuEj9yjSwJQBvW6eezX26fpi8A4X7FbqtURM8HcrdD4rHchzPXbNjpKlCv8
oNrvUhlmUfKrhg7IHkQXFk7uzJ19LZF5mJ9eMXN9w4gXgMUfSH/u48fzYzjkHshCEZYkSpfRb0St
tM06+hkiV7r1Q32XA0loHKySQMxLlgd91y1GwM541IJ3w0X3TjRZpMX1fle6Oy9X7DVVFl8JSN2g
9V2/4gvLDn77mUiqizwmqNAlJX6od8ZBdhee8MPlMaXCk2piwxKb0DodlpMjjpb+2GUmdhm+A9BF
qm5eMjoU4Rv0STvR6/CiS/57PG+Dw82uglaNhh6rl7CuRh5nde8Ld/jPCCJj05YIjbItY0vGWDyU
7JJ7bNMUFJNkd03s7NziDbq78Hc2gq3mf+J9LTWHhbTRhFVUxvf3biD5HfmkysNxWPoW2AvBdfYo
QQCvI+8DS8Nn6ySaYXu5T2AtLopO3/JuBjrYSRlOdv2LHkuldl/qoqd69NykcpOjt1Tqpx+F0Rtj
ehmHb0N6vulAfZW7Fdf2I1dyqSdN8Jsw6vVpfetyax5H2Bg9hAPiWy5GYaxcVnVhplJIRFAxsjuf
R+9/JHAwBoxNSbacg50ELMgrPOpspWsEZUejZvJoFGadMNRYZYSck0khlWN3I3kJfDHKU/2/AuhO
Oxi2B9h50PgvWKTCUNS26RcM+sN4Co4+8oBR9+bIFqlPTFgm3yOfUzkamBZTuXGnQfwtMA4cvfrD
tr/unFMFz5vQtber3UBSNrjfwU7UC934jAOuxNCvYuZP02Ii5B6UIbuioITzcUvDbG4k+cfxlF9F
KfmvyFGviCkjKtuiz6xz4QcntdsBRphvxNNxKycC0XFpH5YpUSleGzsx+/h3f0z6OP/UY7hznhIr
egPi4Jjb7qY/0iXUUs1ZTe1cn4THtHiQCNsIGCrrxBs8qnM7lb4RuK9XgAWEWuIyom5azyAeJ+z9
fx+keOuRoISfcI8puAYny2/PP/YBdWnQe9YY7dm1hCGgCT9XkLsLhF1XW8EB65p2zP30X1odZWzX
Gu7An3IFQMZITMGYueZxghpCyEWByKn64FTnTSOPZZXXfsUFt/t2HAolsPSBjO0eLtu5slwUbM6o
hWHpQcxTLIFDhdaV+Q45PexhIKDy41tqQV4elHKbq6WezKaB9a2bneEPTGbED3j6C+bd5MyP3GHc
jxoYxFL0m8SIlnXjpRpNjWcErcQz2bXcBPdwh8v76x5A8hRr7JAbG4jOii38ABspofn5yzUs0GVS
AsqDQoFLNcM5w5K6zzB0K8hOow09OkSNSz9rBpHRLm4wHudazWuOJr9pJvz3v4ybKz2dTvJ1TXY6
Q7OxGCnfMLcBIHy6GweNykwXI8yJ6QgiTbchIvpCj4uCvN1e7LeeTQ+9FpaFdlsDLaUrKYtd8hjM
iGJB8c9rzBpahcDXpZKRijMBJ9k0mCDCxMF0lDhWp7ChjHX5vX0fEJDQlrHPwejm8o9q9iV+lr0/
7dMdqJ1QGSI6EuNbnvERhtv9ByRKmQqNQ1rTtcJCZptIOy5NENEC824j4UUVSr/vZOcvGs1xNvPV
zCOfkQM6plgdUUfFfJR3HsSPIBhsS5D/T379NDmjWaGBkgMj42keOS2sA7f5hH/yIqNmBpzmHz6R
ibcMS//vXrRd0QlvbkCx0uy4U0jOWzwziZXHb+U5+E/kbRVbFKgr8d2MQXQ3DVn7V7mNAcicpKrX
/eX+eY//87fr/22KAPmgorHIdqh7ADdciB12nvOEEJmXJNVO7anxWDdiop1NBUhLTg1f/3WHoRlb
i9VtJLsZQpAaToNIYC8YKv58tRMLTUOd0GvvdJAQyd8oZonj5kd36nZ34C9+cEdi9PQeVg7sL3ji
19odv9QwUxWeqzsvk2a0FD1sNghzdZ4zKJVzjLCbt02+BwZV6XrPS3UDI7FCrDu5VhQBEk8hFNR8
Gm7sM2ErcGNfjmAIsHBqQP90RZhR2u4tDRdgG1eBNFn0WaZ+65l1LkBBTptJijbFnAMdwEVS3FkH
TvJ78ar87xUvja48B7nAh8YEq7x1T8qP5tSU3cic+nRG6UPoF4NOBlfvvg+bQnvjpSIQBvBeWA6p
Htzmcg61nLr7muFUamg8h6gdYde01qJOr0J0azdf72IROHaH5uHQFGnficsUv/MXU22hrGOSuF/Q
/3ghAy0S87FPr95Fxs9/sd7k7bFvO2IFLV60bJVEuWu9UyPJKiqMFBpywFWHhxh0Il8ISSGHl+dQ
BKtZ/kwFRPbNP1miQjcql59E6dDbUkcGlBX9HNBbmteLwaqSiGpL/6Lno6OTHH4/CD6RA/GL7nTt
wzpKxkKM6Ikopoedfkd4vd0rUAAo9e6MAt970uB5qelKBDm+lCdJtZL9IgFzV2MONc4VY44fMs4n
er62HQe121DctZ+XGDBYM6wQJJQuL4PC+WZEsRYrk2HLj9eB5ZVNVHBiazv73jOfvoYbgLYhVn/K
UxLKkkGfm5JCto0OblF2iHLOWgjHeGuN/S39/rAM2XqvSHakQWtOdA5dvIM16sjt4Vkhib+HVjVg
jnSkIvye8bdrr5N/0/zYRle1ztc7XTbFG2SDri/ajyCHt1gcPsu+4voWOl+RgklpMLkKfNG2UBuz
2eq//SOWfZcpx0Gvzv9q/RdS8HErDDoVfjeHeStqVmWj14cxGene9D5gwjuO9GpvD3iMxNQplxcu
jHMgKh4LlNp/V1IZqMbY8ElJnRvG2c/pBvJmbr61eDd5WMqu9EEJlzwmfuk2kqkz1f1zMv5pbPjO
pkN+vQO80iC5olfyqp2w81fO/MQycZixM6lhbE55JnQtrSu0NITxfBntdjCVmeNXvMNNlRsa14iu
IqokE1VbLLZ8UCwYDHNSoAHToL8sYKq0RTdH9FqNqB6z30ExyHMgKkz+syDA/hPg1jnShgyWarqG
Af5qbpR+h8hCFwkTcjPSWn63x8BPSrOFvoQ/kCQhW9ES2GQUrBPbgH8O5QPLLjIFxs1eNzwPQHkA
bWdWgg42AK5QVNqVORB1Eg4HSr8GGWsb9PpB3kV/gCKVZr9M+oEsxroArwxET4LdYtM585igQ/bK
97D5waHwxxHQ8f4G6AAHzPM9tjtEyVx5365+YobqtrPWIcF3EDEaIDHs4gjxHN2qDwmZDsiZt7eB
FKBXNEJQSXppOoxJQJKdTW3ao/3Z3tSs9rpqoNpaKlHa3YPj/sUvTXyjTSO3DJbP6C8RWS1gindj
9rLmZ+pqStgXymgWKXYh4ZB4l6NhiG/4BD+lf/AbZis1V6DcSuebTHkCne078bLfVnWLdN8D/08d
Cgl3vJ+DlokGaZEuHOoCXKwoMVpfCP3ETAu8b8ErxaQQbmL5oMlQwuMGKbayRHsPT/vs7nCyiVhy
GEGp8h1lMKHsh/8lQGQKbNhW3Y2e/mhZEkFnfLff9N8q00u/hyeKsIyqEDP3McOBC5PludjGwp99
JDbcgGr3frZBVIVUeT5YQRBtsSpr4OUYq8EK6CoITYhaIhmFlUelAYkqmlSlKHBrZPYqpbmZ0o1C
htbEXezJoT67rFNAjZprsFntRvtrx0ojyzEmbVSw76e6fLIO5V+vtlmIsRr50dFb1iT5voeqhWCA
wux2c2jORhIUD7A7scOW3Dmbi1vhwuB/ivXFXNzgE26KsW4qgr8jSQpOD+howLE/zLxwtcWS1uxx
NWBt3xJQ3oOM8VCWxdyPN/yRwbVIBv6xAlCk4xtWODITZ5On3OfO4zVCL/Pqwib0+zV9UKyqihre
EI41Ji+1CRV2BkgCf7DtC1LrzPCcWrR5TV103RzOBH+d5q9LQ7HmFy9qShXWMllsJ3cMIOJnwqZI
9L7Vui2zR5hwbPgdBxyRr1NdVHkjrsJsV3R7S4blvITw/tlibpWo2N8rUjgvcJHbIdBXQbiUpMH0
Qvg0E6caUMpiAY/sA76E5MGTFl5E/Sz9K5hCN+r4tudIKuuXFoChNQ3bPafk4BWAY6mcxvbOWwrx
wLWbc7139Ds8+4aQ4h6o2aSeZUOEu7ON40cWlUmHa4yMiIUrx/n5+HyrkJKFCvZQV2MVJE6CHT31
ZH1KGPND5gLT429UwBcgHoj0gLeSFkMnyqwG3pW0XaELqmLsNy3xctbXMIAZ3pqyZ0ZPpDA2E+bE
Yq47lb/dPKcdnPHca8AelCYLzwUZANoc3C2oO1zLb9M5XXioczaDpB8fv+JHjahqA/GqEDmrMHLn
Y8OeA5yLMsKpS8WwrvXM4GySGbq5NX5wzhLx7QytuumFaKEeo5XTjyyTGCbDAIvZstBD3WvkSAQO
lw592ydH+hhFl/fxtJWh3YPle241lkp6Ya0d409/k2pqDXp/d7leja0/8gxqg9dLAiOOC1quIQU3
Sf2+gWiMyUJKzbsrHaJdsKF18SNIy+0qocG4lZ4y6JDFBf5jBtAb/GOZ/vXDJkAZsOQcDXXn5hsP
vwCi1Fw1E4j4PBxr1qMen+KotibZW+7ihTsruNc3ZI810u6AwwYbDeD7bsgjumEnlAJ+EXY2tMUY
+rFKsk3UJh/nWGivTkR1KjJOD+jsCPJX+fsbl6nxXQcHd474eaR5Rup9aC27jttd4To7SSnsHdym
JVuu5kR5uqZs2Zla+qEnBPzMMhG1KhH8pkIK72wz/0HVbss4CCOOVGhoEp0a/UXgD81CACh80c1o
INJ0L8U5zPybAi3yjqhtFEpfQZAFOUHVTBnWRLEE/J+H+aql95qjyI4d8hXuR6kA/qX2d6Vyyesh
2cQqIS8Rv6ijhVNjO5MnCw95aY80x5cWGZ+47kxwvDY7QVuGMwe5Mcp96OpUzZ+jCZq2NrMeSUnJ
kxWT1cy7r+IZmDoEhPLo6BH0Pa/6BnrfCmQAkg7qekUh/Jrble8BynD79459AXC4k+068fnaw9wV
D3utzekzT1IVoq84X5/wITln0qgsCmiDhyLMgzGwBR1X/eVVdQSGSYAfnchOWdqO//sd8NWu6dlC
K6CTWOQ3YKpMjLQXbtd+D/cPnZd7ZUmJ2XxFd4JYGbAGmnfvbLM0/zJeuPsHVHc+ReO29ikwGk8u
V4kTzh4AUfhqWsaT1dv5yJezgsbvdwjA04HJ6eHiQgxyWPGaAQb1VjAMBYAPsyRhMWxbMw7ugrXE
9mOE1qMJoZeQM1jeVckiMNZS9yI9fl1Z5yJHhtcpmcaADxRGjlCWMub8JIlwnIn+mjU4DOQv4Uy7
K8lloODwqgtV2q/t+EoXLpFDcWs/vkSU59GUh7pt1z2qoqHiK1XIbwik92Uxx+vESaQ+Yx0t+UXF
QQheJingLt2YwjIt5cV3ym5Vt6pyZW72pWgPjCkPJEX6tHfh6HJd2X+KChF8lq7l+0Gn935iyKLY
JHUSaslCUvKxUIk1FEyAy7PYdr6la5LAdE0BpHWjGgUTWcHRKQKP7B/bXQSs4PSlHndiZ8hV/iEx
gJtWSCKPOh6aNwpliyKGsiW49psHxugpDYhqQ7a7tZdlPgMGWduzrhFZbX92JAAgZysaVCnBCk1p
rZAaHjevGP9xiKYGAN+eRIDpzglkFYohG/tOtL49dxfMpF3Eh1WjB1KWoVCtjdGBmkEhJ97r4pXv
t0vJye2O0kTF7pv/eT1Gary54MtMBYGm044kGdfneFrxFhDHkqT/rbhTO8gntiwQXRNs0/nww+Ik
AyXq+/2mVqRUVMV95CaHEjRUOqPO2aK+xhfIhLC+3tvWJvzzFkPbA9o8Si/iArgzc6Ozhok/Y6lg
R1A/4uuLrPQFQWjgYQguF6ILo/CxxtsYzY1rGun7RaySjlR2hoAdNiqVwiXumA0hvr/TAR803Oti
ZFmCDXMLTER7oMSAeR2cYp4/5y7DS6DJYC/1m6tisSqu4K0tGNLsOuseFHhY5qTodQ7+FvNwKBGZ
9oh0v6GmLd+6e5JGpWpAmvSGHP8Dkd1WHK5AkxRc+9d2dVeKNdp4z0FDtIzHDaI7NLvD1hfZ3ovd
2uGrZAbfqMQTQf+is9RTCUPtdb/T3EAJl2lBGKhp278cdRbKxKZI+GwqeLI2V/e2XVRbpfhjxhdw
UPZ0GsXPpGd+6nOVgjG96sJoVCImt1ouf89UgtnviDVlPDbRO2RCMX6Jxc9NR9eBb0r+O/TLIug4
VuwgwwJKB2pQIQK49o4tCLJQVqxityrWbrwyN0WOtUVEGWW7LAgWrL2IYxCrx8S/wkZQ8IDYg9nU
ydcDcajpHVl3vNKjo/U5++6qR1AQi0eFvxxsTfX0A1aYuZKIKuPc1svRlmz9kXBVZygXh7c6vmZM
s08rYghM1mUvesFIp/yORrux206E/sVUfEkr71fqdYFrOiZ3zu0Xe0F4r3pG4J6AXv19cw1va1/L
GEU4xQjMHbrDyDXvuxoTeKaqv/4l5+4bcdLul9Kt1fZP4cgNgcviJPZcDsarFetoVpU3ryRYVw5T
B+uCQ48Dr6DojB32Zhy2rcV+gK0uUkOaB4KVuANGr+sW8xhOypIypFlAabVjqvG6AAtLFToqdNCc
K4U9acfZ6eOgpgCn8aq6lEvvATZm07Ifr5KjjLQJjP5X4HhWb4SLbtdtudYVC3Ip4ieQKsd0b9dG
U9s1cIMLFefkCfNGJoQvBeYQoMvZRv0xGRW2uTjrL4C9j2V359NNhL8bfi49wTBPf5spXCKhkMJB
ZCjZNgP1eup1UK8hVKFStgXRZLBRWNaqjtLkF05WVPANo4RAxLa6JUfEVogry0NE3/AJsHXUBukT
5XxyNLk29LQfByLsnPm+nJPc/rwc4lgLVDZCLoAPFFZ/98+zo/5y5DrLSK2yty5pBYKWg9hOXOT0
ztJUWMUxfa3gTa3SFNGIejt4x/JNh8ZzJtkqeQnyuTf6I9H+cvkPobwHwy8IMwwJo19p/Gl/5MEA
JMWQsmUSTB2eJ9gTlWiqq17+Y2N9HeRPtS5zzhj8nMci05jaVJiJjGUT6V0nBswbNcyGSRg3gZ/M
UTY/www9yJA2KEABhdbcjZ8Dml4s/pgsYEY36BGBPxivcULjgOirX2MCl0GbFHJbWkPG0kIIAnON
C51dty81p7A8r8HpXn1cA2UpLyUe5ZNCvmJj2wU/onBD1sPMLKmR9OZtJ8XglISwLY2SeOkVVsSG
CQL3z7N69mEeM7h06TvMZ/ZJcfcj8LcOYKfpkuAuFJMizKj4l+R/yp3TrwVBfD+RBcvumLNzydUr
QuVkf2BPf3tZXtsrLcNVzMPWeUyg2KHQFUnyFVF3VqmZO2Ooy9nkW02LZQNdKYnSPCWEs4QDbgI7
dctQuIgLXuy2w6Bt0P7tUO4IMIqxtEi0WI3VTD7cPJMqcKUBwwrGABoIECqnVAnHaGTib3uNV4v0
fqE/Un7r47E6DKQZQuT+FCAijJW+I4jSAzBfrio85XjkMT6nFLeX4ASYs+Aeft0C60bqAAwE4kpk
+7OPjkHuHnUcXujxFXGtWNpRGYAFgW1LyY1lPDrtrp616ifiuCzr3W8RFEbOPKgZD2p+7i9gNHjB
Tevi5YzCbvN0Eotmlt1HW1ds+U5vuximmIuiF6w6mxpaLoifrJhZcSb0sD4lQdmnZaz/d+/pk/3C
z/amg/ZMICJ4cTVUUfcJ9oROsnWcoR48PmHzy1hu7XzlJzUGHUexnGGJrOd1EE2Jk6KCk7KlO5pz
wzVoAoVYRWrYF2hXj6ZOEzlQ3BuX16NrXlpXRZ9RNb1FtumwstE2jkFUnioBqYvF7porVfPMr+Xx
cbIDMDLbTxXeu/LIrtVdXke412txXVjzFarNj5cF6DyeKhxlyt8w7eikWhIL5/ADGdlUvr5mkWw9
jIjQm4vEjk6PnnGZig0gIBZV+MlAxuWyqUMGVevvw5MhWr55SVwWnGlfTL/4iTTQKKzlv0dIEalU
wQS8caa7oXBz6yOr+FAKEELM0RTuHVd2ywhx4J9kxXbVavfjONQ2nirfOJLxsa6BAWpG66SuYvdb
8iT4fWhdymgnJnL6Ro60eFk6B/GnKRZ+s1d+TZ/IoYXi5DeK6HwN5+ca1YjhsN0DUV9dEZ51CVNH
Dr7ufWDq2KVSQZiZlkSWubFtB9OC8kvLs63yv6LDnwndfsXxOkT9rsWtkU8YB7HERpgMrhA484Qp
XGoPV2cul7NFfAUks5d+ivj2BecfYB04EoUrB8sVv9kHUwGbgPtnU9QOq4NKJ0zdrV12KRAlZn8a
0BfCDgWqaqhuqrF9sMhvOFOj4N0mCg8eoNDudvv3FPxhKMLIp1E08QxIETYm3JGuap+tXqBsF0ng
0wPSq8XmE0nArrAs09DT8alApD6EZk7Ar9AE348ddISEckRjG6ATddr06TC1ozzWWnLEYzA/AGS1
IprC3Q8eDb9FwbkY/PbwBfUsqdl+AE7r3K+Bobe4818QVgWz1SQR7Lj87qq/601DXJWd7LPCdhk3
Sq1jizGJ38cgq9YVRVhsmFf8u2Hsg7fKPuhkdfr7WEwx8k1TP1mw1ooLs5YIkywulZGwSxyY9DnQ
zXwEb/S07EbkRIUeNK/xJbX2q1NWqH56JdyJmAWyd7MomWoJroT5UHBS5hWsqVz1N6GQC/kdBSGk
X38GPFuRF302qGSMBe9RvL0BjWCBwghse/gsl9+8CAX0Hpem2FMblCAQw7+VFFWSwF+MeWQ6b9kg
n7eykjNLS+a24qby1gRKn1VO6on+y0QXSKiuItJ6mJSf2LMfn6jBK2YdOD87owldaRnzSQS7iz9r
Wp/QVTPSz/C0b6vpeuLjHT4OgCNuXfn0kt2mQw5eFQXGMpAoUMx/eBZnk+9LiOpZb6Zye8uhribf
94dP8+2WeZy/AdeYpzYB14kcrfTMZmFVjHmbjoBZsVwwfC23FLems14G/yYHJP/48D5U0Bhx1Eyh
xOwLFO4bPgUYavdGlNBZFz90EGZ/LqJtt5mQ6hZlhhGiM1GXxXdzw8pyJWxKbtERonceTEdtbRFO
Mr9PBp/7TyVGYmUyV9TSzZfHoWCrknTe4FvnNLNgksLtky4gXTEWtJ4OSLU2DukZeApfXEY3NMkD
m7GOdlk5+ByLAM+WlYYiXI0Zu7J9khYwUZdvGJuz1N7kWL4OU4iOxUrJsij03Gsg8MiI8YAlAqg9
zhUz/ItKuh1Zzq4+rqRM1/1B8fGt6dq6cRo6fhpcrVP+/bGRI+HUAyM5G+C0XXk+cfWJAMFqQn8V
/K+WVegYwOWraMFJGe8tmRXhzwzzu3s2YU6/uezCVZswGUSVL4UGG0uun/msm3HJSqdFWu7qbWB5
9aXgxnqSK4DRWymkF/+8VXwnWNMP09j7Uz5td2zWaHKbhE8UNBvhAnme6OXa2IEsB5eX5qD/8cOH
YhGwxWiB7PmXQOd2s1Y/64+DMXY78qWBAvkRAMwKcBkBuHJnOCHRTHG7ncCL+aULeZfNXwLYUE9M
gUmfFjQkP+kWd1tUy4QxVJb3Q+d2Qo+fEj42y0suQ5dF+y4Bb+wmG5w/x5KitEMZ6z0xC/j19PT6
NrMkYX177A2IahpVRzwfZ/1MbfQBzDJ1gUCyBQmgK/TH6WMWv++k2EB9FLplBPcSX5sv/febd9/y
X5muy2toLem+D06V6T8MmUr8ewunnEKdlaqp08pzF9R4ogJQNaZUqQD4wFd9VfobcUB6LSUdRLgb
1A6hZxYkh7Qi7r7IoEYw7L4OeHmVFkehFiPoDIwcerkUnfnH5El970c8siqkh9UtKdUnXWjnz1Mb
JPHHLQ6FcHoAKyXGOZrta75Sx3vH/uGXOygIBTORPmq67HMvo5FpdSf/74tuLV9+avN2veCdLI58
xhOILe214T3mrtHLFM8EOlv/Jy03xNVQkRvs78Cm4mWrguzFiXQxKZmkjYKbA9zXFuei2LTh4Ne7
3nmf9JWi12eq6qIOKRSRe4HYZfYN0od6e7Zj0kW7AxrV88GufeqlxgWhg900GXRyKyRP+Qs8lO44
RMixinWE25tFB/NuC9Y7LUMye+wRL4C42alTzXADlpTL+oO6DT3o4ge1HP9FV5JPKLUedMVaG5L9
jsSkoCsbCZucc0Pn6iZIKCiYZWcyJ1QQwBJ+sZOeH+8Ch/5EQVx4pjkz3oXiIQG+uW2CCb6EzTzZ
Wu6Q0R1sB7k1c4qItlaPlxiTiO0Jb6rLDSb2yeUxNcL+kZXCwXvE+tKZiIY8KLuX916r5CJ4cqca
RAdfmWfmE2uxVmeouCN733xgQRoVvcQybIhMmfrri/5FoqYr5m6W5xdPDrqv+5xv0nPcneCS/TbN
507nZ41jb7iTRl2gFw/Mleq0eK+eI1IfrzEgjOXFNC9E0DfrcQBswGeH3EhkQCw5BqJBNfMpxYrA
4Gb9KiaaRfJDZaKAsGjMx4BIoHiRNEfOoRpZLY+6kuK8GGv9OOwTsb6b59j0Op19loDhIZn/2juM
05ngpGFrJt2wz6ZMvOSYpEILWEGVYMKEX83wir62INDTYCQhZ9RzeB54chHOSYkyD/YOSFFRWDF3
4mb7IM1MQvJaZbfpxuPu4fa9cEtPHY5VwAxB/0mVSSiPbMTWBLxkhGkvyBKiA8Vb9dNu9akj++Ii
g5/g4+LlsMd36qQ01M9TzGZzm2sLdlTiOHyrFs/IKgSPW2s1w2Fp9NIsZdwb4whsDzTARyShfZqu
0YUxcHcMxPZ8aPpWMZhylPOz+N2V/AA+iMbbFDXseobIcy/pnhaleX4Z4G0Usibe1JZWkxqrHUgn
gJW5vZWqSNBM/2SYkBOLNFAtybRkN4PKmE37f2Cjvi1DIEZvAM8oCGEJwZxQZJRr+8slc+8MRuR8
pWyNyNv1ApKv3xbsL4N/uFcZ8f2R/ykQAjDoz4YwXPQyfTBozwzagPYKuIAp1QqaHQ2O1f1AbqbA
R5ciMFSSlXOvJlNDvGV9XT9q3Wtb4Y/i1+1QsnHvl0EBAACPxQMfHqThs68tmhvlN4hNmElBheDW
RoNHyiF5p4WBL+aPpDGZApHzAvxOm8sjD20wE30KFyOkdTNGdvi3MELNaQdzcPFRUx76x2ZZ5XLp
rrc53RZKRJjjVoSABjCsGzi+zDHl5hwOc2HaWS7N+5hjr7Hwj13TnRhn7Faax3jNOvElG7wt3wbg
ok2q8IQq4/qhYx73DF48Alb4fk3qoBxwce59mG/y4euONF44328rqdZXolrqRR3q1FVOEkoTucl7
BxxrwJu8UqCkEjDy0Qy/nVlLXj7gTIeLK49h348pooSzEnDLhgt53Bogcmweb+DRboYL4KH1EUAt
mwy5U9NUtt7psvQ65+7R0yJgwDjIjjfDKxgZjICMynxf+dnmbf8w8VC8tXhTe8ArYpLTXcVc/EQN
48n9n5tz2X4OxzpsBAmRlVSVbNsKhopiVYKCDD5YHScDRUZGBBWiyMnIZIX9ys40XDUJ0Mcuq7kR
GHpHMBPYgPmJqobUJ/yI9FdN44P16yphn1/9PVHY7G82sZHVEZS++Oxmj68u3jnwgopuvwiy/l23
nHWA/OJ3btWcJT3IAQoCnEm4QLQjGYcoZZnzuorOHWQJiNAJug/cZmda2MmsZ+9RTYOIuVYA1+Yb
Zb95xgCuEjtiVP2hVv3T24U3qGVH5+BQjJlUzxxWepsNLOhUoqxIntc1b8ifiIUy+58B28KGiXTJ
J+vxjTVlGCf7RzgDOnl3DuJFRjHvV8w2zYYdIwEsPEXS6dS1uOj39GR6pfb9OzlO+LEudwsx8WF/
LaI9yAulEZNE3O1RqpbZHTPavX4ezTHjj/QdwTHrjooWOKJkC0efScq9E2o0puPK8vvr1d4HoEjl
6nhEKc4qFbUHJrXOi7gKWLwxy+iitUUpLpzfr5pImZwkllyc2VVRvY6L4MTS0f9SiqEgA/2rzJQJ
wnB5gy3O/Y1gWxgcEMjhMCqD1X6iJCImWI8qdEoTxql+EUFrM0ftheLzqKJ39ubrrregJptAIZEZ
qtb3iyP0QBO0apRT5s2Sa89jv5zAMyXaSK/TKHmt/S07rRmVfDeVPLS5+4+bf71i37xW6Q9XAOPL
1OdPqVyjWGMC7h27MgSkMBq8mO83i2k1hSfaCJ49qtUXDwkHBM6Exn3sMYWc+EKtx4u0n65SXu/9
BVe7Os8gQ5ZsTVuOcz1k3BHiic6wP48g2a6phQxbOEXMKInKGkBjJcpuGkXicjXJ0tlJXOPZnujN
s7d4UHJTwYecjBSJkbGyG1qCGgbvXqxSgtIiRUL3oXwX4jt8m9/UjpzQmisxR6iQmbyl+dI0pshZ
amSeBJ+R/sgOTepfqzmbloNzdof9n+RL4ZxCEomzpQJono415/3g62pwGa1x71TophvP3MUnbVNZ
OKyq7ImMj9MvBhgt1ReCf+FrXUXY81PWfrzhe8iYYpd2WJd7CvphfkH/Yo8OgOHRY4sGfItcZjru
cVmV60Ufq0Nhcb5Itxvfg6NNceQC8UA9yKfpv49m6iiyLbqa17dzOfAPkSvIp2hhLPRzxnBdAlI3
hzrroX0K+K7ZUmqbWVINmUAjb/3SKvp9vUyeMv8zAfVpUeY8ms4RhbGedp7H9lhyyudvwihBa9zl
wWSD5JrJL8YGXimkTdNzJkpvl9fwr7F+rNMoRNfKp5i88ygwNvOXfcCTg0/2BwtRLMnFlEATpr2d
QyeGFoiZ5S0AznF7tn/o/HeQlSrJNVE5Xtw+bNIId9Z4vxR8YtrVg4xxlwMPyVYKeMAAR++Ti5tZ
31XrTAMox64tDA496EHk6tewwFWvRtZ66IHInGoMYsAxbZxPGdp90xYai0RVyHzOfCe86dxEspd4
Ev+XuDqedCA+Jty9dBdMjLaWzcXZ7Lc9DgOv5yp/8FCl4JgdwbZWorQiA1wu9LsxZQkurHgTN/nW
t//AMrOQvNwWcenByDouDuVck3EaYzAVEapen6FRATDimo+QCfNPbNZFNLu/DfsNNpu7tu2dL6He
mHOgCSl+TT3XjBpGUcNq6nDqLOKM9J7YyjtsPOg6w/hh/AESNKWAAXSwtInrcLnkA3QwmuzO0TDh
MIgH1+j/ok05XApXJaONzaQC1ZqM/MJp6al5YX/eyYxjYrdfD6FhzhU8Eq9IG1ez/CRrdihTJe4q
/A7+IGYhiUoZIsUIqLS/jWAF1IvmrfXdepgPCA5DKqucqRUdq596+8B2iUmI7cP2xwIORIVkbaRW
vmHZGI469842h1b0N5P1yC+fnzP3sMJgajmE7Z19+3XPy5mSMedNx+7EygXP7C/NmMZOOrzxYL4E
aqETyuVRtziAw415K3TAELOZatu/AIqejeWb1+tAKGsWtEbZdyRRmFXF8S+V1vQVYGfmeDUl8pq7
Sz5j17rjhtWnL5zEsWas7NGkcqelfVicpQBlhhgC3lJgSR0MqNd+d3zw8Twt7jg5PoKOfMhmeTK2
26JnFX5TWk8wQv3Faq54TDbhfSmmt8Y2krpC3ElJGe98prqVk+22DNlbH+VE/P2w3EMvnolBw1Df
mXHHh8ij9zZFxBBb74LmusCVgu2fOqaXuoiejo9D7/maZqDDbwBnb0aDKtNhWSVaV+bFJty1Smj+
bVfKxvVLNZ1lBft1kHWN5Ez89umfGgRr9olXLOMgMLvceTHaqo6Su86pV0T3i/D131weGGxAj68Y
OA9eVsRSQ1Qxw3636CJzkERzVVSySpYy4m8p0Pvwmb3qThR3wUDXzGG0k7rHIK/WVzodtaFfSTFs
uks2CEqhom1PzkAFDpQg5VzfrpsrDDn/s/nKqLZ66476kKYSwbe14P+YIG0EqJ1G/lx6FNopuNvx
DaXIOkx34irmHqHzHMJLom3+poADBRqlVIfhXADZZMj7pd3d8kH+2Zky0K0kGqUu0rxKClse83bP
8i9MtYFxNRrockWtXpn/PDlwkx3vZQK9hL4ApJipzSkJ8W0VGKH3N0AbPs+UarYqoOq9g5DdDfM2
sue/JD7inWLn7r1c7votWcqxiF4QMzg0tiX6I1yapVCFiBWTm9Oog6q2w6Dw8wfWr3a5EcMdG0az
/ZZMNL42dTl5tVLNxxB3egks7aMa/hEBmqz1lJfpsGe5FUA/ZtxG0LfYGrMHZTq2alPNGdmAQKxI
sfnGbFN3ksOFjrcFn1J9mxiOSo525j4ufhzz8Cs6jZ0yQ0rlNApqjtyhD6auK2U0+18kklLBmLUa
B/Rk31CIUprhH9eq6VLYCEPA+D2OwIMBlsTIte5Qr9d02SQj2g4ZgOwA0wA5RaJRNEEfJCnJxHRp
KotjBiCjJ/4Pztu4URMSfKW4kkPL3rkXbl5BsmXGoF1+IUTbaTuJDL+fjwNtTzqDAkYPHstYgp6l
H6k2hYABq4KmFrIoLFl+vkTN2QDOif+dZLUPSUT77aZniVtHX8MU3N5sl90ZM9yyTQYvEsuNWV71
IPwfjaxyj4IsLKB0DYz7XPImKqT52igDrPFVk39f4vJz78y0H0uSfbh9gOTerDnJpwio+DmoIEcV
ruWs3r7RSx91YgoJqoxW/9vvqXEtgkI1PCr+Oz5gtmcT0puekW8eB7MpUr8gC/x/hOqD/ya8pjio
4Y5EE767Chv/Gw4+ptU38+da0f9+OiuaCMfoH+kjR5rrwa8D0PfeXNksOT1om/D5Q/1ealg1rjp0
wt5j3QbEK8tcJBeLtuH0TeD9zkRCYPVI3ioqrtlXI9K4/JJaMNKMHi/OELUKRl5hsjxTClS3TsXZ
eJNLLin6ehEXhbnqcGIWw2+FU6WjclapFICV7REhevtsGHcoYZoyvz6bsKZYDyR9sF8UTmBQt5iO
2lcxdyEz3TkSYv17LxKzs6xlUMP49c5mGPA6eRIZyiGD28bruQQzs++XHrnzhsogxeSYHlfF7H3D
HibGeJi+w/gB7RmUyZMGfubnLUTPJUvgvYeDsgkqKteING2mIRQA4WqSiCvzmxNdobmfGL61Q/JA
tg1L4DKA+WQpa1RU/VFzr7NEqgRgsSNyvwqcyf0HFZGBKDKQGm4LHg136x77S/iB6JO2nC3jEch/
kPB4Vw84vJ+pkqn2v/JrKSr0r+QXD9Y0jZP9/3NTsrT+MPCSal4zu3boa3vFKK0QX9/LTEKk9k3J
9e+zf0rSTd9jxHzWs8RGGhAaBEp11oGoOWBxpdU82jaerzA8lS1daOcaSJHkd9QLWdGYuMAh2rlp
jhUsHLK00ak2sSYYWF4vNloO2evLv6eJeMH4c/QwDsWM+aW+fVrD2X1PR1eHIBnalg0+2KeewF2m
b/pfQSchan9ypqv/BXTPtBoB9m7EltUcMc8navz+dehkZ/uIR1OnkFOr1o5MzT0+ZEZqL7JrbrTc
k6Lte+Fl4RJnYFprS9CRWc69y954J2eTDi73Lt/0DF4EtYivD748JcIxz758yGY5L1xpm+JtdzS5
7Rf6hxcJHZ+FhL//o1iUr0RDzlb0st9eBvo3yduBJyHHQfKlpyV4UkF+ybhxmTFo4+ggifrLWoBO
+S+mw+w0qnVtXwO85hR75MOwceEFzKAE+4M/tbmV9ofjWGOQRBPXFJ1yoK8tfWDQj+o5pL73Andu
NIpRzDkvdxz4MRaxskHu2JHqknM15vHq+/B90VMhU5tiusrPO45TMJfMdd4Vk4H3vSxleQlnBYi/
kLa4p2rDa2dSFpx32xeh9B+BqlEYqXvU/BbHBzd712sRsTCFqa+4CZxsNv2A9cUpIVQ4wF8e3pWs
hn0zPu3UpJpSBcPnoYrMFasIK0gpOxuTSRHeftJEkLOhWUs5a6q++YAWn+R80YsET91aWB83gMLT
dy4MV6v3Yul3fkMVUifC6LxzlNfgFFu0VNWx/qcdSr3YpHgbin1vn4C9pMrngBVpQWl16VbicqRP
cMy4skJjkYLbe/fcSNEh+zO7Iy8BfI+HT2Td/PBNyxuHuL9q8p0o5yUdEkjVY+0R14TrxtWxjiv7
OZJm4TlZRhOWoVLFmxx0a0lBnIT1hrUOQNJcH3QxvHzCgzF8Sum8DoOIqkup0XSZH946qyCHhdx0
Nwz7KUACSPJkxZHECtKYhQ8yECvnZD3lm1iNfATagG4z/I2Tlc2NyR8hGg+JmMvpv7c7xATU4qOV
jGKwQe04giEE2wLFC5ijbnlMnq/rQ9ivMyT6VSYAecIbUiqhWJ0I32kiiL/Ul6Iwb4xT2doAaDgk
ykcKxm+4Sa+hC0hv3wIFNWCRpjmD/ZDdv3sFpZEsP4B03ldEEAdSZX736NyU9rBPFNlYBWWmllOe
XgC+wGlEOOzm5IyYjb8jQArBlLqwQq3Z+NoecbdFvlnrUMPJLokWdQrzAVogiXXGAuVykgyt6NnU
qbFrqpK46hDG5BrMcM9o2DrrlgT5Td73sW/noMAm/z3FKz3IsyDVbqDLYUp1I+HyCZFrz609n7VY
VnUthiPRV9/V5PSmsiVW3D+mdbnXoIT3PXkHpDWo/NtV75wjGSiRfbjc0q+t6v8EeYEZEba1LQad
RzQC7lKtZx+i2CI5J9i+DTbxhg0W62Jdj49KB44YuW7yQ8w6VMuBMo7/xaLZSe3pvdtYOJdErhMW
czGE0hsJw8B64DI0b/RfMb42s39HCiZyx1xhR1+7nqljE/6vUxI5bcvlXLlq6u0ZGcFrNCn/Dowo
cgm99gcLxxtWoLlNe0dYomyJ8hsRFopkFjsBMXIGJItRjwatJ8Ui4DQuf276SYS3i6RwgrqIHzMl
T5XHBtdm3nm02k4q9ziW/ASmqymbMbRnplQtandai+svk688YpfGx78yi+csMwHTzGmrJU4hQmGj
aR4udCDbpI1onuEN16uKui+lW7GlMICKZSF9OcfLsQNojUEhjJ/nuLsZDZm3uD+g8A5XDFeown2y
BZL0B2/y1r0faOAMZmJ4AtNFUcNqH5TWa6rnEhk+N+OgdoY+4YIDfo/GXNtz5jJz6ATiWdrGYS2H
qkKYU7W4PK0Cm3Q4jtHTlzBOc1KabppT5pOghoRYJFuZlrFfQAkjMYS/fEKb7xTAYfOg8hbAKsSd
ec/69vgAlbRvQEpVVk93Alxo/2lK55HC699pxxpITCVIoN6JhreQsc5WzAOlwp9vFRMBHVy9L5Xb
lD9o/S58UW0tpRs4tt47GctFIi/mLV7A1QxMIWK/yWh22ovYEfx/uT0FplBzd27OEi8p9kF5reZY
039iBGkqBfW4DsJohZ2QL+fIG6vHFtUwyEEAnmcOBHT00CIGTjPSjfNkCBYYcJOAUUMEOVzVMjLG
tHX5Ti+E2xghABMYFRQWQstJJWO6fqKw0G06kI0k37HYIGEvrR0KDzP7lgjAMTGzFz6m4VWvEOno
574D90nZlijTvQ504MLOZMsnaTxYhXk1m3NinXsNKp1cOdWfbJRKRFIW7jPRVMubbWiXEOWzVd3C
zLe6oAlhAaxKPPMbVxi8VDBN+gL6CtB6xQHcashFsVT6kbnSyBCp909VNE/OKXPq6lvW6BhJ0rLq
vAIaGE4pDzNhxuH7s3j/ymaPaaD8OXl806NtAxeyFHlmxP7MfAgUYoypWO5giG34X88dvauR7lRx
lE4T/6ZQRC1bXMT0kR25jCjxclsjZSHanHfWL+PSEhiRkP6vWVYWw+CK5zKtEXNNP0a5qwQMSth2
YRz3Y7BH2iX5/BTsKiTY46H9xC8BdugbC+x2jwN8dv98AejTKZPuMydE1yOR+mmooVXb5Ivgc7Eh
+I7vemL4tlmP6fkId80hDwvv2+krNX26gGFZcTC8+I3EWeHD6ccwTcnEo99YmCSW8BX7Ikb3lkr2
t7zUEHcRt36mcbLWbYZ/iZHX0F0b4taDyCXb8YSrWzLrg1EQzWubFIxGDV0ToVHQr0oZXMqIdP6R
wh+0v+dnFnCQT5xr7BHeGDCrDp+bAQ1odsYhZTi/th5HdUzZUKgbp/5weVGih7z/cZzY4cc9NB6f
QYQMNNhQz9s0vxvcia00NBL48KuMlxWi0i2gFG1QQew9uBoMxE7jSVyuTiaEgFottEy17r1Hy90R
JSOxPSEtEOpXCRt1JTVmCuTKbfXFmXB9fbDbBDD0Ax1rjtAqZsSQyLC+eEi6TP5ko2ZQdH8m7wz/
OD6esQ2RZDVNhwBiB4uKBdZBczcQHu3lfhmSdlrrj+uj1S8j+t8go6l/n1OZTQkkJIeJkP4VGLr2
7LYtA4rWwt0PJcSSrCEbrFKwgYgDRFwKf4O3AXzz/PBeT/bNhSqIWLrBqEW92iyIFv+9kKJLikwK
2IgjOVuRX/+DyhL8By2uouKdjA2XAsYzl/6qDIdnLmmvHkvBq/120VpleJ6m6OlKc6vMM2M6ByOE
gK1hrM6Uya+iWETuLKuxhUY8b3Hky7m0jkIrKE37lFQ7H8i1TBHZ39Sw39vJFYiskad7i4vgDXX2
e7rURa83b/Q0AnjFG/EI43Rk9425ON/DpPBZzd3yOthh1BSYJJxc9l0ISjlRKGKtNQ9KDMmHxDfk
dzfmlnLTT7OmV3hBH0RBEWqcFEHpfrYtLg27jQg0m65vz+roFQYVLlQtJ1uTpEos5n4tA9b1UsDF
tr8C1deX747AJk+vJP4XzKtZ4F9bD2u9QgCZqBdCITS0TenDKGiZdry/Q3hlbrU1LOjSQ2HoGLWX
a/PKs7XIL6EzkL+22zvAFE/+rKDryxN9OI+itmjTI1LkStqJRlxmjpG/PXr8JBlhE/e2e6XLx7HD
I9WSM4uEf4B8CUb2YfvrWz7kWwHEpmwa8X20gRjIKdil2piLAzM6KOnkOWhGZrsM+O+LtMHAT/vM
0UJx2CBmcH1NTNyRK/O0aJNGkYcTMtb13bP4idyiI2aejfMR/5sfxmQ16DZuQNhS4/dI0MkYKdcx
A6xq6m5mrGf7x6yIcqch/qX2jDKi5WhGzsvSW66ftbzB135GWPy872uiPPCXqedvpIU6ep+lX33G
ZKQyuh6Yq5nSDUDveFT+e1SC7C+qKr4GGer7UK308sKwKc2/3m1xM6QfPnmvsez5CBtmpnHLnwCH
sVLIRo3h6et/8t7LLQZvPOq+LhTELLEwhNwqx0cNDULhFPd3T8xu96caiyejYgnRAFoM+HMh3fl1
5lFsRjH5NuFG0TZDsmfyDCjmczp1NBKQ39VHOe2aHjyTGhROUWdex12UhPKyAo24fdWLtHgZoQ7I
ssmGu7JJYuMryBPuhUpxfKMMBFAIsNylZmkB3XNcFckVIavQVbyAdiMvCn7mtrMaXNe0OvjEfGmA
oMMsygXX99VyF/4qfCU3Hrrrno/CSbHVttRfiQNm8FTDaePbQcWKdzWe5K/m0XUsY55KXr0fu0gc
Le2+JVjT8BLTeyzm36cDJBGuhpRPRQc5IGdifxKp1SgqQwciyPl8K7T5D+CgzSUFqTPmH2zeJBKK
oSoavm95Fqavx0oTD4rquiBiukbe72w/ktcsI33kR11niTz0/9IA1IY/zybs3bOY0+sdq+Bt3zUR
txKZmDop6Lch6bqE7oVYIqsstIXFtaGet093w6qW8x2t7TSRU/hwRCyXbuezSdv+DGKZjJ08Lxdi
rs60pg/stFJjRaS4/XLNaMXbPJQdYif1GbLU4hABsUo+ONAQik5G9LI6UTGUDm9pNhmeH2CEbjd8
pF9BtCSOpULPbBYK/lrNL8MymJVfviYDeHVHU9SMuTS0e9IHwFfCRvW3VonNnv5vNcNiF9OKxcWv
PdZvMeb9WI4TuDJgwN5EzelUfKCjhkPADeDbxb2xHtPW6BFws3YGSR5IH7lAPJ/es/gwmydDtPPX
SwzmB5WCH7pElzquEu6o1QhytAnxGB2HiFTd8kC94Eu8t2IprXW3eyP05i7XPzHN6GRyTN/BGPf0
79q91kFrNwA4+nj/q0VWJkx9cllf96pi3cR8qxLgdRICQYaFNEN+O8yfED/GX1/8TbEk6eimEN5d
IroRxf/2ze0YeJ9f6/cUV67wW6I3QYFHxgQQIeZyxm1u5LyoFqJpRMZb5af8lTbrgiZf6g66R/dq
9fh5Z7fxksG6k+wEOaaiTTUNlM4MeLg+o6Ajx4OQjc0R2yPl+ykXHup6cl11gAj69DhEX5Ipp+s3
2+vSCxGxA6wjvrCwcw2vA2NdTWjcBSDPd6zK+Q+BT4DZeczYrrlrGwsY3ZaKwM72uxXNM7RLksVj
zxH/VLSykp62QBYmMGikQAJhFSxBNNSkd9bm+Je7mqTZTTcu3pjNyyl1RMnUjB/RliSz41/icqBt
Iyo2O59NMHxPcaQW0BavtE5esESRpS8YMg7m30uazDfEgGJt5CgR87shr60nuGm2uYSvzNrSmjcb
hiBEopuVd1jCKPZISJ25mlalwRxXSKpGjnRArgBLJkXcg5va+Yzz8cSpeqonIDIJSdKwPgEhwP/H
WkKJs93o3CY5P4I6UmrfdETYsYw2akEvhIK2Wo/cBEPFFPA95SlQzndVRfsZFwyKbk76+rMyETia
2vwfn/dxPzn49og1llC5E1jblobkZjK4WccYhkyECIf20NKPk0lyOsUAujyIIgXQ86XkgfQ/biub
zHYcKyO1oNTI5xUYaO6UTE1mKRIUte+8Pf9pBbUSq6Xs9V2PqNhF3+j2r4OZZzSm1Xw7VzohGnpt
1y11j5WMWtvFIw88z1l7GhMWT/V3QpXiR1ZvFs3lRu+qEiLY1qZ+8712bo6MG0HThNugMrxj7gH6
orA2seg6hKJ2pM6ytHjjoiZEfuyNuFL3u+7AfCf/0WPKzGn6m+f+7TX6O393d/+APiQfnBO99Eno
sSDEE0P7AKWAGf51AM+znxiX4nuRT/Tr6DA6vJWCZ26mEqnwnRxD+BZkqIGScZk9D3qhySWTk4T0
KVKRnZ52StUf+vD70uyFzNUftGdug9oKaquK9Uc7Wmj0F+CvzmS4N7j/u4VEYFOAXYpwlNfVD36O
9wKdk52Su5QTgjtvcuS4ZZAbQOtdaeu/8dpqJEfEQf511eXboQfUWV1+Nd5DETfbrLtQpR+5uKhL
14oS3BpzGbjQS9N+FFsTJx3E7ajnkF/nGcerxGlyoOKpmX+drdC+feTl7fXLfhgVZGBjRmFXfj7j
tM8IgTL7qj3qti/kvOzg4dhx10ZeXeguUvMX8w/HtAYyhy3dp7iGcNR6jRGM1+SthFHQTEaESrsI
lPgukIawYJHHmF5SPTjHYUdpBP24VsfxhleN4Ectyz+6mAZDX8q4uA0HpPXUIKpC6Siw+L0HWFQB
IQZjZytKNRJnlyCXNDidsTTW0eNQE4uyzx8DKi9DV+XE81yaODB7wFkhVWmtJF2tGXRJjccZjwAG
+7LtM4VrLsViRNgDpTgcJI+FotvTYFmcl7+jOFZWsyJwemiJ0CrGEABJ0TjNc2INBlSJDtdQ30zl
Iu63w+NxIYF2y94fUKzv9Oylxj0zKJOuwZr6Y+scoud027vCujMds9B37y/EzB3V3SURkM4MwPJv
34StVBcOzdo/ugbz8+sIs8DINuqKhOUcIrYDvexehYzqR2p8Ti5JHgvKXKBPt+B5lEVj+eGSrOZa
ZZVr7TMDhtFcC8vjP8Vp/C+ar3tbav9Wbd7gp956uTqrlrEqsv3cBen2tF81Q8RbXzr/581GZbS1
Mx/D9iuttpQbB2o1Y3ECHDIMnL1/kN9isSvxxg8N4pWX3rFd49+hJ4zLIAiY57xabtVTaxDhlXOm
3Z8L4SKxFtrFgMUzcW5XHNGRV4cLjXfFuyblLn95Eq8QC/7KoGdwIHVuXje0znFVRel96gR2vgAl
fYUpxRwJ9ypELgg9Z/s+TuaoWP5JLWDKz/WoCu9aSEpxWRzUCZsdj+D9kST/oed31Yooq8tyYvar
W7cnq/UdioSyraAEkLqL9eeXYpAkILJVNXtssQRyOFwQIx2jSHEcSHGMu0bLdj1iQPpxJCddS+5E
gzPLRdcTrAUj6RtxJdtgqLiUJvkZSK4Y5Vw+TVt4/P7QiEd8JrTNm4I/BYGGOX3AVeZAoPSq67aM
eMBZ4UCMvuK7bL/ci22gRC/JADnHHZxtlyVTLWLolVCWrmyixNmbJvdE055B1hctBF0RoYaeBPT/
3Xeagxp24b/njtkmOdr7ReqtJfd3FxWs47kwiGllajhky8RZONSw+Vbo0AFh18x2uTzVu6N04TUN
2J9nLYB3n5+nl2h4wiYGaHp/a3WZ6zgmbFBQFHvLSTbXrL7BpQGThhR2Qe0tZAjW67c2BojXiXdc
cRxTel6FgZqzCtxR8RAZGMRwgLReFntLILyrs8KW4UUuccUuFqjKaCuj+cpS7+TB3+Al/zpL8Q6+
fGFs+9EqGecgGVV5JuaEwID6mJqvO0ZwNU3vMoDcXnjsT/BYWED5H5KWYWyWoHInHKZLgYwDIVVF
3XNua3eydCPt88Xiz6VgIdd+03IHvqorX0qkZTKRgclxVEHJaPOBX90zl1g8VOmJhYGtjYFqAt1p
92qIyu+FOQDrwt5Bd0ECJ1c3/Sxk+vcF/q0KKhv9Oe1GW+QkZTrJpOdJU5WBsjQ6F4g4tgtxZ7O9
HVatyz6cDDYqwrv1LVSrpXQNj3AzBMNqli6XlUC2Pzqd/JW5haXaTgN+mitBibUj/rzP8yJebMgG
IdmgOwm/ISkrKAWWj+IdS9FHuFCdUBpX6uy1WHJhkc9laMcrIKhv93+fF1hVMLfFiTwgy6Gu5bUV
hNL/KIbYffo5Dh3pPj6l7UjvsgTXiTC+TLqZ+PRJf8Fuw7cU5tOTLOye+jAzOPsKPn5A5g7Yyo+1
mSluyUeKgaf1AJaREACweQ1RCzX1alFONIY8odVXUsm9wTrFPtogLy9jz8J9eqJDI45ATuwJAUXN
XxQLgQcZqzPFmsTO16GdObgPP15V+z9uOxG1DUkrlgVmfQ2TyUmGgG+mj3L8w0QQ3qzp0J8WwDjw
SGnxDGBGOoV8Bjg6FUElQezvJJFB81p7vCHUGBTFWpbAzOKtCEBv4txyb1H4IFNXu7zyIpI3QGnH
JO68vsmy60sFUZajkfLOr4rdCE2EvLRqKcdM76dWiD+C0sqz0NcqOpvwUIp56ialSa/eVDrQW8wB
AUjSro6GeRjqY7WyRW2SuTCwGs4lDWNCrTnbmyzccOPEVqDFFeVTVPosrgGyLav7wmwLRuG0LabO
NwsXaA4S11ibra8B6abTDDPcfahllGJCHO2YpMGG5BRpjuV1OdiUsBcmc0wmebHfCh8pUH8n8Zxw
b3STWkFnhs332JLct+yopPD7mnh8I7W3FhOWtxb6Nt+PPW6YgCmk+wEvfQBaRf5/gJCC9PsVvkXS
EfymYF9hBCFw4KqHvps2GrnP06OJg/6kpcRdaV11V32j3XFW3IGIbcA8g0slLdbElH+j+50lz7Tt
CxoAhrbtHfjL97Sz5GLlS95WoQmHcp7FGYht6ySJF3QYesT5Kr4b4BigkCX7enfqEqz20inrVQlw
dVku5ygWhdcOr/qEvdciMK5LmLzOgB8oOGSI0gH/QRBsy0ruFvf83rWou5Lc2518seXOnLWeYZwB
BGTsF6+9s64LTLVeYmKq/2cuc3Jeh5LJqoVSm1uHPYnn1XxOug9utWO/0Dw6AoBkx2S9psYYB80m
roeqp0bUfTMKI+2GiN6cONrJHICy3EErNaspMUH69UOB07pfqf1qE4Q56Ue7CM2prBJBuAcverW8
1O3iFBd6pnO+JFs0br+9y2Ha4OYv6DK90X78/B2RSqX0LkTUHMYHHw+G8oZgYtgXlw9rsGwNiDEh
QbM/fAQRVdHfj4EcSesTYi40bI3PDJZDcRcp+VBb+Ar8G4mbJoc9578f+wp4C2jPnf4UYJVw0tVc
st8RnRgwXpKfET4aDB2Oft+mkVjLNMzN4xAtA/voM35jWK4QQ8hFw16g+DigzUSfl1Ba7vA8tx8F
NDu6/ozL47De7ENL/HLpMIhisiEAyNrIQE54zeUkDVCOUlfjjtqVcyPwxYhO4Wpbx78zspfr4MZZ
sEM29NW4+6Y8ZmlMwsLJbWJF+1QWr4yGYTyaSvmnPVtt4to+rRNgdquIPsH6bkfs3D8U27X5tSsC
cM1EGX1xStC3BGJgtbY2NiY3wNR35f+VfvZDgwzRbjfU1HXB+/MR4twx8b8THs34U1aPedl/tMcs
66oxZkSXKy1rsaz8l86UPLIVuE/asU3Iwmga+QD3rghAwvVvUU8PeCFRRFyLeQBtMc53uxZSFIVr
oxfUZLdOSEiT1O+YkdQ4QpAAQ5km/c2LgeAbKvU6/AmA3uxaT6UbJ3yL8m12WtavsyADOTS0HSLc
HumLkNe0Rsn4wNGiU7/SRKQxYoVRe7kCBOIweXiRshkezcnwDi+VEVY1GRWcnJ+zNSXfJpDANw+m
lXIEhREUC9uEH8GefAVa0w41mx54kxz65IAA+a4fDgZSX0sZ8uWfDs5Itu+fdQ1u8MLzQqHvK7Qq
/i9XLCfRBNhAgKnAZw2ljwPh+P81gDJJJPgZizg1uQkln0GEB437LROlGiDOtHnw10mh3GMiizfZ
ySnN1upm7NMIc3eFcZLxauP2XCbgyMqyStsc+BP43DCtsfcsyfMstNlsVkYDaemTCjLOxkaZ9Pr9
UBnGMw4u7CU8XSQqgSCcyrYjRIjE8BYkAwiUAAnOPR5yrLhzjlj9HrIC+6nG7PPA4LbEcjNshZon
NVkCmMX8E65FH5mOeOU8WiZQJCihPoJ2rV9ZsmRbXa5uTxOS75z8gZYpBiiUAEvp3xeF6P+NGqKy
cvCxvw+6gxM1bv5XTP70dXSSro2c8S3oxOQTVvOjwmX3WtJpSIjW6L0E7f5cwnyoz7PA31W86Shg
7D/1ghwL0H5PNEq05cEyAlHvh3IbYj2mTXEuVfrZAjz8BgtycH05++2jxULu68oCZ1ujICHRQMjW
vmDeZ5lCJmrNJAu34qbsxG6WMHTaOIYaSSpKzOn7wnm1x8aGx+HhNvxcXb6yo+X+dEi6uFwxMA3z
dXLu1/6qcWQ8jv1yXG+l64/dK1YjEavkLt6kHtqRcUAtZAqCS1DwVwy+41gwvoglTijNfVTQeg/K
GcVqxqdL2OP4aytYgSuJvokPTAqFSrofLOMYwp7+5kSxsIVP+dvYj/tBNXKMUGzl3tTFO05JUhg3
aScGIO7+FURVyXSZCEuHRE0Pv2565gdK0flpUieM41d5NEGdxzKsPMQO8FGZThylIaZ3/+v92eQg
FO5cDHckDYDUT3xBEpA3ya2V0jyvoeo+lAIme+4YaYQG8SpS2v8wkmS9G07IkImRVgtVJi/PzsyU
iIwYlNkvfcY3oRfsDJPO7uBi7a5Ho8P8shAJ+uoCyKEYXpoOUl39RlOaFQG13RMjo2fRBjfqbhvT
m2mt0hpwU7Yw1BPwcREdRswqCLN9RjMMX/IKAS9Bwy07F1xB0YBBGWHUhd7Wnxklv1cj9BJya6gW
T3EiewLUh7L3J7dSEFfMCp0dNkRU5rhdvGY557dQayYc/m/I4xjWCjS6fgDIJqGMEShZCxS7E6n2
ZzcFcK5SLgR4j9FS20y1QKELTGJe87rMfpB05csdg3VYjBsrh8u/ndtxDTCEVqBfU6GLNsws+ndP
FgXsXkfmFOQOk1OXWILvGAqBiLPXyhJW/6J6AH+6FaewSsQhcwv202J2NNvTUrk7+G7xL7n/2/I4
PypaM1dN1Ymq2AmYCImgEjRUYZl1H4Wtq9cfHxcxCjjoMhMXcxOPbHscPXg9eZX9JFv9khdRVhhC
KNFfZNfOtTqsh+ygCKfZfDZfgSqi1Cj1TXvfblHPiuZDjBfHAUAqloWjTrfFwqUSpt4tN1n81KpC
aJSddqA7fCtKvo9mMkPedNOdxjmhM5620fOd3Xsh/sTYi3IQPjCZTYP3/cICZzUcb4wBMIgu9HLz
7wgRGFNt0uiVT1VqKVbwvYp/WDAb53IfwIpqlWGfprBjPb4cLMGjjVNAZYEcLU8ElyygQCf8jIUl
VShirwsmSXMLF50DNJOZgbKkAvSPi/V/MDzZ6FuKvcVxOCAB36r9uyI0hl+Ms6aotdbbqxJF9twO
lU/Ws33K5OsMfLd1DDL2go7g4fy+kvNZewfhwl0BQ8DiMC/2ubx3YZsevUIpAKw5BwTrVr2azCGy
vWQq3CYDQNMEe5QPbwE4G0dgEn6velQzwIc2AbFK+nHE0mKAulmcR4I3g2+A6i1tnXZVx/3inOhj
TdJgBYyVzcfZWQpXNS5f8svOuX6z9OK73aqZhA6rOkFh0Xb8xrtylhW0SKh9PRnC1j86ZK7+L/6y
drVka484hpoy6EOHjJZzriR8n7mcWZK97WpVjpsGX2/x9Ge27Ans9A/ieBfH2YmumvpT4vv+Ri0q
5XStYpK0gU3kiqhetyF0LlJwNIFtnf6d/PpP62irYEFPjbcamR6Mav1nmBIIEtGs26R5/kJ14AAU
F+SfmBtTS3CHjxIDSE96OSZYowIYamlWlu0OUM/ZBZIgLYwA4+4P1EAc9W76DGNIxEr3/j63XkmJ
yr41tEdedN/5Fi4XoYT4BG6bg3m85MUA0upftJqAPG6UB5D36HmcA8dafXjGrA8+06wAxDTTsPop
fAmuo741Qs10fvwwnXrdEDUHFR4pUn/R0J9FRyVssmH80fBdKjkwgc4bKEoOQG9nGz99/3GM8hBf
xEIhzCw4cNQ6nnvcxCCms+aaN6cFe5QedBUMCCSz/FNbo2Pw+e0+a4rJBz3VMCrLJP72J4rQAkSX
mtN1Tz1+whexyn5lZdMd91qsIwttKAT8HXEfPiC08Bp4Nzkyj8IAlAg+b1LUocisukGqe6UJmdMO
M5VMJrwVKkv0iRwqI9M0GJnyqZQNBXw6GcagiUnF3zLUtSmjAfulUTSzBE4Uorn6t0IGfoPEPMkq
6/ZG1W3a2HjUbKUdZ6GRNIOUkTxgDVRfa/rIqrc89yrVoccJpIOrkSuzhItWfU8phUQaQFPk2wng
AvO08fVXGtClldf9ePQr7F6mLMO8i7XH2PwHZCYtVzn5flxhHFm2Vg0gVo5wLQhs9b75HW4b32cy
rjmtwRG8/jcW0s8pn/ExVhc0cFSuOyaqjrHTY9vW/LpvjKIX0FeP6DrRq1oDkp2ll/oGsC8Tq0wm
BzglYqHfnN1QqMxo0Z5Sks5I0YU1hhWmMtosH6b3ouy/QKIvF5IMT83AX+9vIg3exe2hFM49SFgR
c34NdhHyi/55pb58zigq2l8s/TGv1Q8PEdxSftNEwrW292s5klck/+xoLRbFIpx+KKTKjdWZUuDS
gyZ2WYeploBLlDCYZy6gcI6oAcUTUGlabm7sUN/MnP7FPlU63nA6MBECr4gtNZAxk38IiGGVvriP
t+QS0OGY1tB+5IlWl/JZnH9B9bF57PZ48AJkfcgxCod7ZYIpRNLbWREOgwEHFaTCslp/heSaTl+S
YmsOxWYsg79cfFc8qcRDiv9u0BUZ3Yfml+An5RzkS9oRXcgmF8ebGT7AxXTSVU6NNOQl6v9d2KBn
udY6Jw3C7TfS2NfpvT3gchii4jLTDyVxY6roIwUf96hA/oRsffRO6vRJfMUh6rcC0+SWXxTGs49c
7QM5WBslRXJh4aLWXZFmu+iWWh1sFtCIxrkzP6m0tMxuT2iFjiEiH1gscSbKF6kQD75cM50XkxDH
sNhZ4hTPw5+W1KUCv3/H0XwWOeiWkgJkvFEt8stdDafr4yksdZYjnghfqUedJ8E2uwnzsx3mcGFH
V2eJqldUTEJyxubg9J4mDwS7kqSJ5Brn086gHtJ3EyOcRT3f3FggQ7oGktHQZiw3SKGmgmdtFVNr
lfED8Wwm8+0tQvFCE7W1+X9zpGZFdwZ7S+PH/x9IvTMsCaFkwcxz/+VdfeO3hxsbPURG3cMVdJ+W
HV8glilMAYKEe+1HTXisy7bdlEFCg6tgiBqOW0hZzR0oVKc+1wy6lGcdFh/n4WDuJslMjWAbziR6
0VbhfDoKTCIqcr6XJeqZEqrK7Mum/bke5Ggq2RrwymSRgkx2i2U9B1toN2CqIFhMw+enGhXDk+jd
2wJ8rzkBQcJkg6uZVePXHneUun7SYGqL+vmTSOJ/R5qsdA/lrbgd0y5Au2XSZffgTODFpLHjiV69
vkmkxn3M9o/5tuPP+TmwQu24mUk5EooWgkgieNKU6DS70gqCuB7jZ2dawLHONHPnlTcD20L1inPw
4rST7cAMhhg0hbk01RzZ92NDJKf6KkbHQyF32M7qlDlU7rrkHm+h1fIB/6FzjKa9+3nFlnCN+MJ+
wVDeeDuuAwR5JVx7XozR2fejU3xm6Kvu2sgZ8pcrIZjhdfO3wDPvpEML8lllkc5fytYoAoVCF4Qg
mOpXw3QyKKkiKVev4KFvqSawQxePZiSrcwHzNrxSeEznvV4OLU/S4Xo0IByRgRAVd1fgwg4VAG8t
/NJDA5kNuZJCFx+iDIWXJ7hVPQ4U2u53QrsiuZIpLfcpNG7vcLevDf0Gj3BlFHzVUJX28ykUPVkD
fcfEFj6pI7fKdrWRIlZKm8I6SUVT6zQK7dso1zqw1fwRMeqek2MvWYOj6AtfDEflSnIZRRVMycFK
4ExEYhvYalNnIQ8wOztcuVvIDFLg/2aHUM0imE8Ki6abPcuSinC/5M0gy6amJJcpkdegG7Dgk0tN
0wxuXaLB3AfT6d1bdcRB0cZo/qmtE9XqJySM3oNahuo8QbE8Jvb65UBYX9IsocLShzvFAYSyVjds
B6WwdzZGFWztcFRzeHqcHBU5MlDRfrCU2ZCety2V/fpK0vPYuV4SeqoLnUs1egWEpySE9VUdToGj
KKMpIxaMEcn6G9p6zCUcfDfA5LKCuAFvPE/EHdWqLkqs99vHDf7gpZ6NkvHYX9hM7xCwoO/U/b/X
DdnZC80BI2+DDfvNxsB8/TqD+c5xMzI4z72RmP3TYzEET95oaB8VDdGiX7PAS4vhblMZQ1tGnBwy
Ob4jRw0GYHzjpMkh36MyO40lJUAG8n+hP96UQ6EXITPKhTYDkyUj7Jibj01JMpd80mO7QUV7HIdE
pVl8i+6un0cQ3DdSyXW2jkYSKr14MluF+CBZaOU4ikAYJzR9AujP6YzsC53k9Dwmhs7BdRtjLyVG
7XyKNOQECFm0LNEjfbkU1pLdiVnCVDpvKzw/UL0vi26P8MRoTloM2+kR0bWY8Ticiy75bVsE0fBX
mPdjIEPTkXiaPRmC3FE4TsD9cw2R1SfHhepzmXb03EtxvriOrdYQF1vTJOtqzkpvMWo2zt0WRWlh
lsthGpH4pEmoK4mwS3rpmHKI3Mw4nVTN+l4oxP+YJrERrPXnoemupouNxMFjeUwcD17sRIguuk4v
tFdYsdawtn0YF8XfBrjHrddqW1/SDlG5KJ+Pziqjp3GNp7KP+tsE3dhpMEgJAVt4ORAoXmvg+LbM
rHPW4HIr6yJJhjmVLJsXH1Vm1bPG5Xab9lAd4xJDuggtKzJt0YYBhUtnwaDPgWT1ZMqEBWmg76cU
2HQiE2NtBBvT0nwzsyY4C8GiZ6jH1UmbN01ru8F2Qa/eRF08Rmk1ADldK5zlxVQkS75wgUqLgFxj
fQXjig0gO97S7chq3X/rQmEkFVbntzB78IHfI0D1rgsLy46XCv2hjth9kFpuXXiUmCmF7FZFCA38
Nevq5EkYPcMIxhDL/MYd5GGTXmwNW1Wp1r9FXhDHVoAKxck/AdS/bBqZKa+53VDyTHkZocNRpxrI
M7ETqZvi6Jg4raLWHobEujk85w9d3+AeHRpRbBEpo18fwToHMmMI5Qheb2sbTFnWwGpweNFyTq3F
RiG6hocmOYbSkOLBvq2uaAuTMJEUGvml9LzLpr6G2xagGpeE+FoTmGiC4RZEB74f0wCWVqurhBOL
BX8kHL3MfK4jTIBo/FTRHzsz+KRt01fjWsrgXwYYVRmGLfzqL/YAuCL/K5dwnRYPi6cgo2Pnb+y+
+MIL6Tu4aQ57Y36IkPyUd94rG6ofCeFTB9WD5nfXDYBpP67qIDNqs41pISFpjix040mwfE0njEV6
F46cJlnwPLLolTh/9vcpuSrHaSYRKWXb+LxcQ3mSMPeH8je2K3hBSqZ6Xr7213jhELlVwZ4/ERAD
g991qqqlZ8YCgH3auJsXKUrRmc9qwdruQuOcgLnt4VSKV6Ec0IusPXOb+OKAQZ8AvBTKRlLvM15t
XMB69TuZ5oyYbUhOx2KPjta+th5Slh2mPlSJ/EZvMSLi1eot24R/R54vfSXm7Pq1fowWeHkt7s1C
UoHsS+nWD0oiXBTWg7PCqUqRgqpZHTvH/GcOPGDVfROK6YWMr4le6KjCyjQQNjgAnTe2kX51NwFK
fvB1aXIZN8c9XgqD50N7rriIDMPQco26FHRTAWecBB61ef8Dg0zaPu4SAmEWTxxBev+tPP7GqfNi
cAS7uPOaKs7OXjB5dKnP2U6R7TUVQ/bh7arHGqH2KPKCddbCnkItloPATpXs0pX+TZxGtR00tJP4
b7l/26Xga0nqZZTCgKl5vrfAHOazgAMgeBkRTwZ4zZMm1UZgdwh/LxvN8q0GMLBBnXkxV0Wyukgi
mpBXVv0sMktGV3m/DAz3weZdAXTeL+vyt3H6avTmUjh0K8RZB+7GrS852tsDVxESTyhhJi3C203c
F9epDS2/ln1XovNAh4jWRcZix1JhMJgOUEBpu0oZBObVhYtZ/nWiiqQJyhEJFLKYelv/U0AmTqXy
Rw8YcaMMlsOfI/LA042KlOqGv/SbTKQFYG3p8WtcvEzoGY6TSf7iF1XLLaxj9BzXoCBZ3BkAIb1j
ZxqsAF0zwkW8Babi0HzIUXPqvIiC77Q+GSYvG+a///RzBLBOnRAgpkGixAcCpGc/r4X+RNOR/8lv
1Bpa8Rhh2eGu/U5XRURv25AR8HO2nA+VLgeXM2sHXvhUquoKfRued1oG6/2oueh9JscuwgW+sks+
jOqLOuon8edGlET4Fk23K24cAkR/N6eiaeBbsPpzz8rNHBQlt8ipFns59k4Qyr0Qiwzgddj9anye
4zgS+9mNCMj4XICFz0BHSi2tIUbj0uaQqH9ygbh1zxWZOf8/pQ8tGIiT8PPFrQBn8hk0C4+J7z3i
Wy9IeKvD9NN7Vd4+Bi7neHslQMo4poXhNFN6CAxEIA3oaoTzyczuRfx+NlGOUlIWsYxb5NI/t6dS
FGuFQUC4Ivi2+2qiFzqS5RXA7J7lJydaaDWt6KWYOos15wUoKixidjhUan4WWM2WNBEr9Q0ZV+yH
mhc7/H5jD8fzLz8MTVaDXunfL+30BbTf0YKTSnYKmXZYltonP9o7qjyqqARpVnuZUNvKlIKKdYE0
/nH1GyKbm6bosUH8FHTXz4aKwmc4U47+YmhMQVWOwztgCq5sEC3PCngGH+kwHhBItU1au+IKXVuz
nWiMeDUubfjqSLhqJlSeqRDOf/UREQIcoJ/9BocDzmYqdfvgatjvHL81y7rNwxbuAqwCLphuplTm
veIx1P+zJb3seTQItmvMWdH0XmPfyIJ7NYS0KvqbjMY2A+VGyCRqduwo/f6LoXEh2Li0saRF7vet
Foq9LXEqNEXf6qiI/Zgjpn5bVnLa492SkaaMk1doUarY2eb+eeJ4nExqnjXz4VNH0CGVWzXrESla
3gleXdo5KFDz2q/SxxxgYkhlICsXaQBiqXjGbwWDzuOlgj2e00kZKDQw9tbST11eIBe2P+5VTNIy
6DTu+YgyHiDTK4l1FA95m0fP59t1RbfyrL3wg3jLhOum6/cGYfR1f5mjGPhRQdkVPcKKuj6/gY8h
ltkKBU/eo4uZM+/75v9nh2b5FqyWrT0XzWOPXAjP6qJzs+KKCDnLsPgm+qJuE4CQnMpSoE5oC4bJ
CfibCTpjS8riuSXO+9LDV8yHL4VQLJj6NTAQVq3+gQSN0YeA4xd9MRBiF9tVlLy/8nIRsS2sCXfh
kgFftfJCrBzEvPxi2Cj4NJJDJAN7J5IjYoNqViVCmwG1aixYi9Ygk+oTj5qrrkVHzN+RAAQ5d/Oc
cILW4pytezvILdiD+AwOJllXPoqrkV1DoDocVXBq56mt5Z5cizQ1kchWRjx+w/S8Tk1m+60WFh+F
lXHBFMI4NsQh6aSq4KjnxZi/mmrsLzj3Ilz08d5m2NA1ztbV+5GXqI8s1aCBjonrVaasU/6anzbB
I2P5cZ/Cel+Hs9CNgEJhgh3f8ldDKR+U4glHQa2D2KN1v/Qal9HQiPLW1fN321OfNK+5AipUjtkZ
ZzGP99DTqu43RLPsFT25qu0jZOlnMEdsLmeejwBEZJ4JS7CpBwx0+IlEvEbIsHrdFJBHzmOAwJgK
y3my/CQ+HUqSPkSGpjy0lj9NaqVPP4zdWMGEgf+emfBB71DyHlyxemmBY6M327QMPCVDshHxlXhI
FmCmyOhdNuKCiUPE8eYikTCTX+wgynjZVhrJw22c5nkpGNH03xm0xqTYk71BNqP1zXSItNTQbgV2
Xvl8mS9s9NRZ7vp1d2Mu6TS7InlgcWraMelvmiCtyKx/SVl1jMSF7gDZ6e7tnxEjP2Nz6RF4hNuw
/xa46a9ZESJmT/WIuuYynDwQ4GHkAlHyR2bnKxNYalKzGW2poFHMDPk1HsgDPXIdP+QIpIlhHQZY
Sa0cnrg0MdF3vOslEpuI4opD6xoBmKxHk8Inc0/fIEMW3lEVWc/1e1GHcX6w40Fo02ndoQ3FlvEQ
QQuqH2D2f250wSBsvkVG+N+gAysHaho5tgge5z8mprP923OfBf4Opd8mMVQttNdSLY0Im9x4pK4y
0yovB3ATHLLOYDqL/482/Fwkas7+Q0NccBT6rieCq1l9C3xfSCH9kSGj/5AgTEUFfa6R8X56hVzs
9eLbBWgBrfvQ2LIdVXgGf1QrUMG9knrj+0mOe8lTVuOjeIiUAs1iSVac1qUxahaSS0+oe9ZHD1UW
js5GRHvm6BR6AJhwIJHqkOT03BGb7mkDZ7ROOE1YtNqqr+VCM15BoI1silR4yR/3OD7nHeOs7OXe
eyah4otYYdsDO85Qvdp5rVRS6XL2Xre/iOXc0XI0XIrA1cehefOHQVglXljG0Fpd4UzUQ6GV6agZ
18AgPlntJSRHt9ElFqp8u+3hz5Bmw/IKDh1oOME4s39cY9yBKjjjl9JqtlmgjFXmffAl1Aby9/f/
Mn8NGvn+q3kZVRKSMNYpZF942uZes9jgXBB6KfyEgSY1NHsTLc0hxxJXKabs1sZZTSCzyyAwzAvT
x/lJ2ir7/L99TqDf972zj5EEVZszeCIbpuO3d7bzbnlsjzmH6Z+1XLlRREnq9f1nlncvv4Eqb/GU
Iz0qpi20yUBVbbmrAiz++BxtyULFHVDrIfUlzJr8uJNcQ+HoXblHZMHzxOJwbCTLE/Ig5tVVIYAP
A8Zswk1iwQrH3bCzTZXJFXyCnDwl6bcEjqiDkxyEWgzHOfUrkXvgY7MTWQREtqikz0IitIBpgN72
1Eic2kSqfEqVZHhbHfOW1OMs/BS7473CAxXwQ37rjtTIM4V1RZMWfjHq2A/juBYYu24HLxXWYkOs
TM+QEzYKrmp5YDfEBeRP4oVNK/7lo3lkscUFdCxWPCwldo1UC4UDzqOlnCJ4esdDNn0g3V6bzRPI
ddz1AqBUHbA5Ex7hqcg1Qf1jXkqSIxyoEK5xO1Idm3QjiMn2V4VgKKw5DRbQvr/2VCgCUU+bd4lH
8/PnpxmaKU7CRIDcn+5313q57vXKHNgL5IHxA7ZQavp/uFTIkbOPOHmkfGBta2tCiHFDrsP0wVjX
YeM1WrVJZmv4QOztsy/5lnXhl0lgscwJQ0XO88XcTQVkeqRC4aX9/5u1vLGkV3WSn1VuEkvyQhQj
jwDY061SpH9kG0lc/S2sl3Xuca4AXUcgfcAiT5w96LvzEJjBZBxXowFFUO1DVhJm7jtaYL46ZcdH
cLLjXbSBY9tP0wBY3kRGT2t/xJp5SUWWemlkPK/FHaDBc94gtJheBbNOAMnQNjOfeQD5ENdYSPsm
ie/RskKXUq7NA6LgIosDQX60EZA5nbZ81ADyYMg2bDO6MGtTArKuzwmayiSwjYgp27rQTA8BsMFB
90rfTyIUQ+f79/9BHzKRqnkpGwP3ma9IG/tQGmvwXYLVe2Oi9i9TnH62KgBWgMM2QT2ioIynLoRN
ZWtJ6BhjKK4nsPFHWpMuurZm60ci1dt1/WMPD/8PShD0aP7al5EvBK3V/4YIPxUkJocK67RXTDXv
B3wb4j1ZdCab8z2kqq35UQ9lA3TRkX/zrSLjbXCEzP4oczeiv2Pdxh8+Ao7hzoHveLNOkUaWZZe/
NyQz+AV4KNv5v4sUzHk0OEHrjzTer962cn5EC3tdLUiJRSoyod6ZO2T+RxTb0JI3fA5VWK2UYBT4
M5bpJzGSv+l8xsYBW6pl2tJ+0/XSnMJrBQQA4OvEg2Ack/8Gt1r3C5SJm/AM4mjHps+biaBaszte
bTOoy+MuEMfFNE1m8e290zE7iZSe8HxLAnnXyqV8lvTjt6EC1x0FKT82b/D2Zqbj38ZEg7kkJOGt
OGt1MclJG9/yf6TkCHgr5CJE06KtnXy+Xv7pgWDOaGAtqSjSn9N6OttPK1bfokGvSgaBvCGJFveJ
ce6RVBw6vosHI1wPbXHRnFPr1FjrA53LVRgR0O9PJRe4o/11VyhgbAXKHuplTBslap0YjU/ISkEM
UA68mQZYnIcUwDwh7SQ55mFoVVc2N027ujY1/4RSxCUmK6bHreArL2LVzIap0Oqt2KX0peuCpAaA
33PL3rqZXJKpu1+pwkydhGkGqe4J6U18vOO6eEx+HPtnXyTeecR1PQyFrXgiQchoEC4t6YPuKMD0
GPGX0jp0JjrNDzUKZBk6yaizghedBZgeEvVhUW55SFig4T04/j8F1PZ3U165ujwcHQrkFsQaf5bY
if4HYyWG1yxSZtYEhuJnuFMLjv54sIFZbD7oxolQ1IE3AhmSc7eVNV9HNxFDfTzAhx1GAaZOddSb
CppW7WuSieT1SfPI9934bFIdT0V+gCuCzkH6MJ0uv0gkqjfEPSr0hxoJh64YYTm+lor5HqR1bQXw
wpKMOpfnZan8gZsfTpocAluMspV6QtOfCtweLZghZXHu5+442RsngVbiIrs0GMA0gNYPWdYb8v1N
5thuyarMzxKjqOi2qX410KKDiTBFw+fKFjiuDGx6YeJoNOo3RJP5iZ5K1Ldlnp4AsBOsnFdNPRIf
TWeD4Aih3z4oWcn4W/HzR+myBFLL+Eg+5+GjGNtErWJyIbcftSFRZKHVDuD6xKkpJmdM7JiJ20VH
W2/HKFM7/5YfrlqwOoxptUumZidFH2mqkS6hhET/8cIMOup2cGAPq/i2BDAcItz3eikkz93NjEYE
BGvTuRs8jNEk45acVTVwnHgY94Y+7HgAdFgvBUQ/VYLiApprmvwZv4lbSWXDUPMvU9AyZPPhrYsK
+ACey/RcoijwUXQX0F0bxr75WkjXQHnFA2RUAcmzDxpoNS63mp+jeU04mD/3a3JYxq6hUyE3d32f
DF++f99WzSromZEJeaaQD0/7Bju/RQ1Gw4yzDbNOcv/nMQTAEJOX/KmGW3JbItBtVwYxYHijqLD8
YuBOIPYSQGMRDKTDFOUDxTdvnH8oHYfVclcP+RMlK1gE3f+RPnov6aleQaHuLI0fzi3azzLk8e8j
FYBwY763yV7ldX/mB/U453ycYJGYlOIaGchGVFCXbXBLv4CyLfO0IVVVYR/EPHPPKqPr4u4iu6cQ
JdB2Wbr3VBuD4DF20SQN6bWtJI8uk3CXHU+/yXCEPPXkfpYrqGDksiHXDaIb0pUa2MIeB1WGAajx
LUJwrafsRKy64mZji9ldcbnsmOjo5WzweeeKAKdqQHtVK+8ZwubEcmhtCw74SzfjWxUGt89svq7D
XE6QsgYRUYQZsNh5sH3O8px4BZHUv7naYRQ2q745K+YBOTgBU0GvngtuX6XY79Vzrmofzuhd92fB
rNzdf7AifVwOF67JdNgcAoP2Lp9bKegTarSwMdYiNZkGCwhhx+IUran1hacxtFVocoiuyEVoF+PR
/9b4WZqn2qRaOGv3+ZJrL+Gy5zr60BqxloweGLsVkSpB5rxqlpTJn0G6B1qulA1Unx1n7x+rxilt
yJRnsMNMR5gQYCHETCdCF+qtB5IF1gvWp1C9bTJ8R/y7+gPhzEXsTTM7RAjdKI6DQo20Q8RXGThC
nJwkcn7YSOyAZrZfe8htt6ACXKrbC//Bxqsje2rlqI1hjMA2DMlvqbaKJ7wWcmbF+lBCUTmVcelm
vEqN5k+g1UD4BZkl/QD5ciFatPTDen16NS4iavIWIu2P1PixfyoLZVG9jgVGHlJxagjiddzgTpYp
WeTSU361sBn8ia7U5AW/4eP0/IW1w/NVYd8HzU5w0h7zwbgn78d0rKWii2fteDvdAxBSOkyYyrRx
wDvdVO82uRW57cI3k8z8ohyK+L5K3S0Vxbc7Bk/aeP4jSjvkU28axKcregbgdJrdy5Mp27Kbvc3X
1or6APA5+1Dugr8CSsnfwucMGG/OfU+jGYI83UbrdiKiufbCZ6znz8QvmRYiwiJIiRknmJ7bY0ed
HNRwjp2VeElDAqFRwSXVVGPb8zQ/52la4Oa2lad7H49Gip20CKUSI6+7u8I/lIsRPq2w4pUh0TjB
hqhPo5aCg3AqCf95oLp/KxKC+csiRV85pmKzCpUCleLLP6iwBqoApqKzKoBEPXfePhwwU5er61j5
22/AeWUgu1iXl36MG0jsRYW3JrzCoh+XlwQIMqrQlREHmDWhRn6dDqINzjcAqs/GAfwrWdcuR2A3
m3S9QYMsn9poa7+pESWTWkSgqGxH0QbZ00ZED3fBLrHl0cjLMQPhkz2wQRTjyd9K1KAGel5bQpv3
91jmsamX0CTtlmIHMnmXBBUuM2XUT534unAZmbGrzI+SF5exY0LKQIpWUHP5U31fwwn6tNUptaoh
qrCi5RtjyZpvMY2yh+WSQQFvPO0CL/VWjPXRBtpA364om7xdcoC3tdIXdku384GIB4CToQJLUKPV
BJTPX0Z/9qdfxPxu0AjrMxRw0e92lMaicEPZm/00D2XSWPz26nNdvTGCRsV6Nn0IqM0MmdQycP1o
FgmSqS33aYmCTuFY1RpMDbMZddNQre1G6rDmQTGGj8fglUzKjBBLXveeFgHMMDsY8/tVHXXKigo1
n8aAtx/gqmzTE70IowoKL27IOqkwIAcjZW467mtKdfkL2dq/WGP7aS0xwfyYJyZL0Joztdredel4
8lHYIqLAgmzy3GzX16M9xLGCoTnx1fa8YtNkvZkprv4slFzRy9Mp+fmXQ+5Tfv8hLrqURU8Es/oW
MYmXYsSaN4Ho8WMeUBULNVWWZGoG+tR5uTXrr67Q7uXUWS3rXFmZdZZxnzTxhO7pmP+7lCHhWmhe
ggR8yXu2q/M5iHS4STN70dafZaydPe3eVXeQiluQYCLilc0cVGyuCEMIRICg5YPGMiNQW8YDJAeq
gSrNkPb/xRzJ6tRgqiqxChqWVZ14gCA4A2Xy8qhfyoAcMviTAFg1/vMpgddyrw5hJT0zr3bJonDL
Acy84y7J1NRJoopP0I35wRK4FVmU0Rq1xtsA57wyQaywpK/ntDkSyar8vzOzD6Ok7ed2MsSTYuc6
utdMgF2Y9RbTtsDbxq57fy4KYhYdGCGg5TB0fRYxXqmBmpQXRDMkpwIpkpsIeEe3re8H4FFXAcky
ot7jvv4KAK0WBO2AAtwiOEiCorz0nIKy/KW6SiRQF8GYDkIJc7vexpYE30UJUTSmIOKhGwAGCqcO
3mbMZBKXD+MzvDaHI7hdGmRng5SKXkfuHmpTkpMjW89xEOUbdFtdEJdiUulpRHJzE5srJJnm8m2e
HmbsK+5fOc2o+flkEOyhClvcp7E+4Q3tJF9JJKPf2ITSR0qd6d1OWsDBX4h5TAjMbYjmmHvax9YH
LAUzYbKtMGLnleIMy+UJyxia+Bv9Hrux3NOfNod4roijMTNv2gwpSZNtfLEkoeK3B0IBWEmOF9zY
KduCrOjtB6BOM/FQPQxbxTpPoyhnwvpDdjQ6cjigom5kq4sBAad5MRBu6y9pE7johxL2d1zlWZl9
TIFa7E4R0nm2XsaxCREf9xzM4bI2DO4oGGmd7x6XcCWOKq4mzR+Phi6SV/LpDFgSOmY8wX3W/TJw
03omFv01x/J/L/VyXOhzE4OCcTcusfmfJ3YIlJH67zLfZ21FIuBNd4xvH83rCRp5HNyf1NWQQi+X
s80PI7tr1CQJH71jBw5vofM0MXXCZxy3h/rW1+Y+WMv80ni6W/25yEjaL0fjU/e4VYMqTLMAwxz3
J2dG3V2GEpjswyrokq8+EoZIAAFqCsfbvG9ZIrqPGREyGbjsl0ea6cgYU41hghqFX78R+kSU9dZB
FRDn4VC72FskRWQBaChOh1+n/zal0fT0abS7DPLiXjPjfzTVKkmoipJ+r1vEvg/vCY+GIsAH6v0Z
8EVeiS1bRQszXCq1Bp3obXjPtESyOKiaZZnvtkP+e5hU6dl6mgzNCUHmNLkS85DEsAf134L8rhud
pRdjoG0BdDHn7cpqPqj75HGKfx5vpZLbpXgik38uuA47N/Ojbd5wJ6d5vg+nQh+Lp8EvpsYEYnW0
5wTbqRqSQbw8ouQ946FFx4DK/rMc8mSkoNE++jl0wBYR79g08htiDGBKmGdZ+ZXWEb+JEU/qDG4Q
tTKoPGBznLCkCIXbBsMcfsWP6h8jxB7LoGZZWmrQc8I6FaqGRSsGkMAQz+eBFAeBU6/b9+hvmLnO
aJ6j3cd/EsroTpVdOemzOFihnR+SS/xeBO+4mX5JmCInc96gWGp3MDaC5CNFDXAx3cuAUzStAc2D
eCYJyTFDYu8R1GrhtFFtpfoIxGsbYhobsjSICaV1oBvZrwLeLamWIGhjmR4tQnrI9s+HIdsaA8BT
lXQDPbXgWvfhr1mo008fyDuZvGlbS9igUvNTEk939UzsKwAEIpFr2j+UT1SNVLOtPLa3+pKntgeI
US4zHYwG0AG1F4U6s94owJLumiuexsPdtyJE8Jtwc+/492jXqXH44R/g/7t4YYC/ZW+dVEr68QIc
zCA/Q17OtUnNRfo1NOZIRU1wUz13spPnrff2HeylCSSWEuG2jfa+f/f35WYKUsndGN8PnfKL0dit
tJR5hpagf9sjHt7WnHJWwEfXdmm57oCdH+Ynjw98+1BRsgl9DxK7hDd2pKDXXEZDMhFsgk6jT38d
ESa6DVbUnOis5SlwGgifnVNsHr1XuadxGVHNeGn19lxpOpREytqMDGIJgHjWD3iZTe1QdtrzobNQ
AXYyIMCj8l9un1JcgOJTGaV66SejFZ5A55ALdsbtrPeAD5+oyxH/PZIBg1+6qjkPwH48861ustiM
JMYLkeITwwuEWNdRacpMak30KS7ujrVCJAotb8AtsMkEttY4DxOyVvS8AubGIC3FR60zakDWwN9g
LV594DtPl/RjY03w8q9KpL2F1RbV+oz1jlfPnL7mSbGsxoGQDRA1W0ZnYp25uskKWKpsXFYHThJt
dF0ux/mTowriXNyiXsJKYN7hfSxc5OroAOML12IDM0ib0C66dW8bDGJVwMJPBXbN3tOj4cKvGPn9
vSm+lX/IoK8QLiOIe9/MPR0jy3t59iswfcADNiltdulpvcKCfpFHbCHS8IWhkqC1G4doky8oIgzp
XrOmfHUA4MsjCvJWkt8TiAXUkPp0hwxnotbDIwfHvH6S58+ni6auIae5ETfXWCzzW/ZZh6CgkfHN
/I5DFSGRiLjnnEqoor3502LFuEPvM6WyjacH4CgAdAuR9wbsaOvSJVUBIyFeie4fiXAge96FNYy0
3psx8mQd3zqWA7f0pAa39sGhifdHcM+4N90KWySvuAy5AhGk3tEpbHersjCOPcD9e1H+KG3q+aDx
+GG+X5WMdpUuPuzVXZ3064uLvULnkh+3l216vlCCAJtN47J8VfLE5SL8J2+4F1mKz7bUu/XrLUaZ
fQ8Hkl024oIyIthJ4G+3u5oWug33B+9j7b1OF0Dw35wFqxCY7joggnwZB42UxzpydygW9eSrkA6z
LWZLZ2wimx8hn8FKY+UA5CRzxKEX8kkF1UfxSiqQmU/iDytR7fJe/LWag5O7GmAGwQ2iyUZ81N6y
i7PYXe1HbC2A4zf8JjpnyKHTVIB1aEbT7Ctwz+n77+VsbBR86WWA9PPljKJtRDcpbbz7LyHRHSXJ
C9C/OSybBL/6ND6f4K98P/MrOYuopYFs1gPX8ATkzmGbLk8E6K0oNpM8UjWEk98SfepAuMNlU7BG
lfeJQUj5EsP+zC7vOO2FasrFHuMwHxHDPM3VTR9Zt0CXtbVDugCgljJTjo0aXQHtKMSmNMo7+/X/
8sbYhjx0wLXO6ezN+C/+Kt+pMzzjOHc84B34d/bVKckM8h+eMjldCuivGxZWB9VqsDNCmrfNUZCT
HzxmpgCNQmx+xv85FO12q4zrzV3lGTAjCyo3RQCFvFoTJLaIyTHSkiskV1MPhOMjMyz+wSkrHyuK
sPkQLWC+yiuKy6Kmlb1oLcQoWQvsNX1D41FAddI0UjXe6sTAtAXXlZZ6TlpcqN8YwPB2uYm9Dfjs
/fpBsL7zWmrWA94hhLecBGBN3Fh18qUkGvnuOmeHm1vR1qAURFD4RP8Ul1vqyQIAwXLFYBAeGPQ2
1IloxohZX9O30K7Pitc4fV9bDlmNai/kWTVfuUrZbfjItYQgRsK0XWYSV+h9/Rv6T4flN3issac2
8sY5LXieISYyQfFspSqxE66N72ZQx8VXsMvlTdOf5DZdHtthE5icFa2loKU/EHjyByuL28fC1DGm
fwvkoAkPs5f4LwDGssOe4VJ7tfHCn/kwA75jZnAJ4i0hxz1wNQfSUydtT6SDo1M6jaoNMULIAv4Q
VN6TiqMV/xAXEkGFQtCvOM04D/D1jtuX7m74dt7PONsLFso+gT6MmwTDP4i3lJW2VmcVE75RhXgc
iZ4vLAZCtvbwa/r/LPLEc7JNul3WCQQ0vifJ6NmUDfBC/jd1SivUcHkZ0Vl2WbFkUV4huD4fHm51
iFcpvPrCVYnTh04FTEa76WHxZjgkQR2NuEh/Vhmg7dmxdYKMzBPL0sdzZnMLlzdEHqR9Xj3R8Rjb
qympK989+ydK8Sb6Xvz9j2CKSB/xkqU0UOiU9xjVRa9Wo08SEoBP5WjUKmF7no+FJWlstgSRjn+h
LdTUBCfQmbBLiR4gMaqabHxEBsSfGAcwCmklM03Q2kW0cZNFK7G+m+DPogPW76splOSkOdtVj764
vQgi3qKgLCUOAb1fMQmHXkKNSHhOeAsI+rOMmUd2G4mgbsX2AI1PZmjXrOzjuJwz7OJj/A86iJse
VsGHSumNpsif+G53rM4UGrvHsEXjRLHwuKlb4ReAwTlraGnOFvL9KBRo1jOJ+iKYD16Ic10A1Lxi
z/zgwzyDuufAxquK5VDD6aRXRMSvR3TtGEUbVw6vKLBgpEFaHBzR+TFLn8ASP5P34df7o9xrEqiF
fjyzR5UaS11SBGLyCvKEAtTiqOKjqIarUCoTZ3XMDY9nG3CrMLZXT/brbq63otzTdrZQLpW2CEE1
MPO0dZduoAZ3omSI0ZWxOwTcs7vmu1/w8B2DPGF+9TK/uqXwhgSJkFRizRNExDpK3jsXLfV2xFdd
oMRc3MvjMMA8jtgZD2EBNEyeGCtKzn4T2eZHzwmkcti2ee/vYVRL2v+KdpAZeU/KgEn86RjIdyWX
8L9H8WNXMQqq2kIr7gi+/bY+hFIKJgSEeR9cWKcUh7IDbHLtxtFRVlH6CzIo4YZmhIrMVAcp0qtL
zL/JBTybRId2Bx3FA0G5TJ7pJog+xbuk+1dmUw8X7s0HelycP8fJwoBohPHNA0Bvb29gSVdJvmZc
iY3FFRd+sjN7JONe+PmRu2TErGXIpokPsSmDogghbFsvK1qq9YPjD5vmdOUVxpHiDrO9ze+xU5VD
aASq2AgXZUDiN/kmOoDbog+zqnwusHP4ldDoWZobWfGlk8mwhyFIv2XccQ/GZWms44MyVl3n9QAG
QBzF+0sycw3xO+hIof+WhPgiv5nrMBM3jfbt87Hrs1TS7avZrEeKvpjXhIqLxqV5frFw9P4MCLzG
2zQYoSKL8qTdxzr8e3B9IAd3t5br6g/4H/NmMANW+UyN2Zwv19yvgTwcKu1HTb6Jz/ulzdMLHsr3
3Wq7seSC1x0lxP4emAnp4U0lPZylSmJTxZM3B4BOWEqmbS0JboJMSK8KG7Rmm3nU8un5xZTHKWOq
6PADyMnVUc8p/HQLH4yAmpyr1CVwezT9sm6Y6wskjI6jRyQA4SH1aFQf7WNRsE6jPZgLIxc0ljnO
ZCU4Q6uY3lwaQWJyy/bPCgl5jYuw4MUwCkHKDwo1w4qAlnRv3DICTE9PXthcfY4yyjflssXqyF9X
6v/HiIbl8EoJ98NXyxJK5orhWHaUbY9qwNN8Wkgu+d4gTbLYGoY2AUKODvdiPdZXeRU2tVM/evE5
DR/DUoZBF5D7KE9byaYLA8rU0CxPsNgTRh7Oxn3YcvBDT7Te7TghzL3IUtBLpMRn5tiAU59n9mYn
7WU9AiM14OGDk6xQjQIoK1YSPW0FZMCWY3mkfQQAMEdgeW9eCgZ7kcVrcS4y+CyJCAHXenRH+s2N
uPXmYHSQ5nlbEfd5VB1uDfnB9EzG5YDJTeKG7KodJ8+zINX/kSYib5a/AWae4FILh8UPnXQOmiVd
NafluH2kqh8C/wpG0IPKlit4psRBYxrzPkizkLdewVF1025vWvklMhB7VPfj5R4nSA3byeZfDXH7
R94EsB/VONLR+uI2ycw8R96VM6bjIMgW23IKGn+LGc/Nsq4LFctrDbklYP6qzs9HTpsycMNaxbri
Y1InR44X6To3ORva9b5G6FbZV7KeTWim574vWYD3/GV60gCNRylcSd0woBUnT3Ic+Oy8s3d4Rhql
CdA5p6AnOR8OQYRh6S3iWboCeHYk7q4PEQ5oXMBhijGHp0wjYbX37WZ0R3DYWr+XrHpyVheoYTQi
No9vTueW6K3orNB2RFL/MwEQekYdPA4udmbt/+JEiPpTFAlxXFZNTX41162o8skxTuqz1K6RW2l5
/ixqPt/FVJYPYiBR/58Oeeo6Y/GPXTG0MIwVzdajTgpI5Ue4ZW6fdTVBMbZ1ODYP49Ehmq/iiJCq
stiSgJwXFPC3yoveSUBnV9BafCFLzuC2cqH00WQfGsd9D1QL8sOu30hfbZAtBYtMSVjckbeMrAD/
fAfsqWek5+6pw4dgY+VfvwVNfRvnY5CvU/EngXCX9z2+Yo9be5UsYSvOpc/MyWOCNSjYRB9BbMo9
rWfaGcrR6651CVN81IR86B/moN7T47tqRwbev4bDcmxr5+UGq+rdow8/yRLAYu2Mr+Q/7tAk1bmh
+V7RvJ78DxbN82UtItGgSByUrwERsOb7a5H6MMkhjFzQC6xlmLoEJOosUqXDvXINBgXcSwPk251I
V+fE97zV/IAlJuOlB3hkfge40McKEqiUXZGjp1J0TwKxK6w1816Hs8NbEN3ZvVDYIEo3BxzQIPTM
7nYyS1Uvym7PRZU8ehiypXXRByj9RIqVUtU9s1W0zzeNzfTm5ZaeNVPdrq6FzkA1YoD5n6LAQw0F
HZHXfzo0PyllhzWj71yOS9bbwWPraYxrwAPp/O3ayJRb66Eogoann+pU3Rbo9HlmsBlYBlyqiSXh
c7j15YbxBTc5endcnz15jf9R4kxNtXR3gEjSJe2oILSR9UZMqLdgPEE0SVWJ2LSjzXskIq0trQfs
fKZhUoairZXt9tBSYNDH9hv1a8z3xJttUbIo4PwZYuLMPh/FeqjQOhFx9TDEoetcWgMJd5P0uS01
/tgT9GDPlRsSABtnUhFKl7wE83ooNpARP/xw2hW37kkjyuIfGk7klAkzMsUuD53fQ6ogopjl1yyS
jhFK3uE65nUX2TsSSYX8C5jaZuol4Chp8x1HTIcAMk0lilCFJfjxgpfQ9GOoHp5ANo5G4KLaPOv2
zs21ruBFPzO2TCZBlPy5GB96Sq4MtlMKYbKNk8KoQwTylB6SAeb0RHHmc8aey+0p0bVpdTwO+T1W
y85EMJGdHT/AH85wuFPOLOp7A6a80MTSKMGtk9HBJ5QIarLw3D964zNI0hrV89EQf0i2FGJAfofB
GexkYDGtn58WWYAtY1rpxkluYbr3lf7ZA7KiV7Qw/p/VhoJ6PTMYUiuXC1uT/x0oNyEBgxyBmnyp
za3GUEHg4zODzsLqzraG7dozqIDnOrEEkDjhH8m8ZBPDeprNWUyvcjiGSuN0t2ACNtgYou5GBApN
ofSt1Vb5Y376ZuecdkQLKDWgplQwNT3naU9uJGet5bZc53eYvhEEZkd1UFKlMqcDHw2QreHE7s48
5JMeKjiDIG4sz6xC16xl9L0qi8avoSAYNeXXVlAs44cfDX07HjDWvbEJZ/X4Y51gX7EzSy5uF8fy
eGrNPtCbvG2k0zimD15kvU9HiI+ifEwL4+hfFHdrpEBXnRIgwKsb330+yZIVCaix/DNrnx1awTj6
MnDw6ZFcXp+HU24b2jIfzWRUeywQoVzNlMn9GrwhJM1xlxg1Ilello8pN1MBTN12qSpz78HhSFCh
698xxVp7OoOLl3GF/err3hti6psu0gST4HuL5y0yePEQZFk9Zk16Ttxa8YNuSvXipVDWY0GLaat3
EQHWnFIqI4C0ORE3fRWxZp+pFwmTcVKkAB1YEACInXt5Ie1LEBUvB3UHdF5OeGHMbRxV4LFZzvAO
lc+ZrtwgNBbgqpggH32AWwf5nAgUjXKK7jTJ/hIyz6GizvQ9F+sloV7ScyjLy42eMivI4/JppBEX
JXmkk0TJho0X50D6mnNA6NHZKOcaXg6LgkRewTMTz+A1KMQcmVrp3KNX/pN3sfOI81OE3WDsd588
Qj1g97fwYkvC0EFzE1JqkKRR+962ZQnz9QUMIsg2FnN19KpJ4rOhc4BCP6tUYitnZ4zoenADYRPo
wn4HnpniGPiRK22Bx6jTxsCgBMp2/IC4h6qqwMxNXWG/36me21PtXojQnvNBWLgAt2CW4TlEqpHi
QQpkrjVOzx3RLeN0PyN2S6ooL5MwEQnun8C6VYbCTvImAuyZbksPYkzlL6pyU1QU9fXvVTpuu/XG
2dSKno5h2Tz+EX/lI6lvYK84Wnl9OA+E5rPnqTwb8KGyXYGzeyJ5zAod8wue8bLF3jCdjas5cFua
w6gV4g+re9dfvfdrtnmzY7ZcMT2B0uWgaJErUbggZphOs19ETbU/3u11UzOfziwrBpJxsUqAeTuh
OjfY2Mb86KbANU31+fZ6RTi+Br/7PwKaD3QOjXEXEjyaXgLMHgfIIIkolMc1gMPLg0wmczL5Rr7q
wLIduMyBTcmudWZcYLiXsLYWIwWtQc7YiTvTL+DYX88Op19xXroqupD72QwQk7odmE6pCEtr8TYc
6MAQaJj6PQ14xgVBZCkgpeUg/VedRVYYLJENIGWRqFvOAMLk9YLSpG20yILUszrlQJw5IBQrv24T
TWUPuC01c+eT5g7pk8DoTV1btHi8xP2uEuAz7QJmVauolCP9loArDXl8tzfY8AJYLvle+3rcNFQn
JbB1cG+L6oGP0ZvL6v/hNMQh16AKIy0ELK3pCYJJCIok2GXCEevpS52Xv0ip276upyBLpX+c181J
zBkETktaZVuurWCwuyh7+XQOL+Y0t/ZfsLL97WsPyEa8kHQrrxT77aWg7H/hcnBRh7p2sZRQjiEy
SU4GrB3fFr1ASfKDttI3A+GkGm+tYHyr22Au/KX8ukKdqRWwJ1NwfWaCq0zTm70wlzWtgYBTYDH6
gTrC9HLuyIMW7yBgfJ7qMz7bksemSjkD5mteyD1ueuuIanZWGcRzWdv33GhL+Mc+ZSyoNJS8xdj1
9xV8aNVnbgcT5u0U/NYG/47dOXMtDxU9X5qmF5iosrWkXG+J19pt7oWOc2fM8zSMmPwf+Tp3BOc2
RGe5QBlNGs4cZdn7qRfUUDJBth7LpTCJaY+mIgryAvGMPgXkMFbDLVAgB2w8efXTIJA9ntrZFfvC
laNBD6SSLVMt7tvh5ayPLrTuXMCXNUdg1PRtO98V4WDi6p4nBh8Q9mccrdetIYuK2r1MPMvcxsP+
ZFWuzR+28aZx4Aalw+PwNIwzIbFB9i0Uqg3N9EdZg8SeFd5cbBXURG87erYN3UHvZ4DZ02m0SkVO
J2olO52X8SeASJqcxrT0SO8SlRAj1v6cU36fKVZsFvutLwk+6+kZnprWE6x9w2XS9ZaedzW+CDw5
+fsrVn58/8dzCV65Ngl/hqFoe2gLDyFezylmrtbO+wVcU/3ZNOu9MxNXmXfgXkpqBj1RY7IGm7hc
HAT4PrYrcAtrcv6N0xq2Z+6ZCmDVfKN4Nv0QzlP9PSp9aiauw5MNB4lfVPfrtkiuFOphKM20iGMO
kyJGL5ycuvLZG2f6EwpzrVQPpgjiSJ6ep4fRp7TzcxKZ6aTzOZTzk5JGzduqSmM+fHPtF2JA7B3+
0ngcbA64BFhJ5WBVLH0NofKZyS8y1ryRGUE9CoekeENyluZNnjb+5TuJd6ouJr9k2+wb+CMn39Tl
WNnLTXaT0VnXKzvXgTudIE8ygMPMi3ecrgyoFLI/19C9tgN3XOIN1abrUFnhlBYRnfINY9uXry9B
PA3wT6//aliMyVJHrvlcQMLezsusW8JOlHX4s/0RW/0wAo1TYJB6xByuDzEJLhY9zwnOzrCnNpBm
V5rjSVBv4l7DgQU7B8e4AboJNiaIf+F6VQCI88oIspVP2+ffMeG2kOnd6tsi9HrrlVNK/jC5Uy9Q
NHpZ4H2HZXUNilU9hfZ/sXxWCR4q8nixy1G7ijXp9ujlzVZpLyK4y4nEGk19kwzHqdN6hoTj3Rb7
tpkSYnhC5mrR7GN6sjGvL8p+gxf4qE+almAYCkz59fsGFkQaVwtxFZDsU3cxKcRaetcrXLnECh1E
+R9rLXzGV5NJwEl9Wp1E65PV6IIXqpEzEzhdlt/cetAQz71bKK0/Cm4QsYT3/LgbBRy4DxC/0+FL
QKoKyQ5KRunrdirS2SZW9mEkoKxXDWTfpytiWld0jTpYXi7CZNP4LQJsvD/t3cvFlqwMb+q40XM5
ySNjN072TNBlgC5GdDoc+2bXsocluzMgPHLoeKNUguqjEpH5ujEPytMx8tqMBb8YGQQyPQzd5QFv
Jufyfsq2yyXIuLPyoL4W+FNq2mVoed2AX3WP9voiE1E0VCM1ghsP0MxqvbaiS/HE3CFR1PVF2hSn
9LhJZfOqCFTmAsDdBMYZKoUuciwetQJEbDRG+1xQCq03RjFCWa1/gNHMJJt2gCmyvM/pilFxRPem
KzmCrEwJAfOuEO9YRioUD0hwKhd3Twi20jzDWrd7X1uDdZ7Aa9dAOzjK35I5HH0golyZMoRkpjNM
hXlKfjhLZ3zPkCE8Hal0TMKqXVMhsOfbvQEnFbjRrX0xf1XaTP0nTjv45fUWleRl6en1gDubTNsG
FZewkSj+EWaKhFll8TtZj4HEQUfT15s4uyP61PAVMlyem0l/wN3NW7dT4Egz2EzYC8OhrOd4sp+C
fixkUpqx4sUEQ6vVBl6WHZOlQPCMdDjKA1Ofp9M2PYmkBLUaLd4LxJLm8kaWTEFBe1t4h67jEO1G
sh/4kL6WFnY5Td4qIv7Kj2t5lszPmM8D0G7TqNtyLMZleKrlSODXqAaEa3PypfiQGLQJpo0+CtTO
3B1O9nc5yVCLe6TSmdnUSWSIhSbSzc/xnBf8bjM30qWBg9g9yXebKS8h1oCt7wU34pssZ7lnHAMB
+rn3WUWqSwpgAcFShcGxskqL/DZUmH+uzoq5hEYIg/pK/3FNFPyvczYGPX0SnNdmjphy/QV98MUR
wId801ygrNvEgLzdJIDqLsElmVAVd1VzN0n38Zi/IrPCxfq9FGX1HHdeWHhspRZhOd5lzbO56gWM
gTtMNdffC+YxA7ibIr58AhKOMSHqnbCXPqr3R0XsFCA8PQ7DEiSFpf8hdYpSohoHoTZob4JcRiJu
mIWarUdkHxxVn4EgkiGdRjIwAjdluR/IsoWHEK3DO31GG3by14uv7PDbai2LlIPl507ST0/2yQYz
woswBUkqU53uj+bTf9/tXmfSXLhnQm+x5KRvmSEw3zGq3c1ICG8wfjaho8pKqexPFrllNc6NcfMd
Am6q61CeZ4mk7hWOooiu4T2LoYRm0PHOyT7VjmyqFnWXwDsxN0CW7y7EgcBzZE/UPd8YjJ/tIIJO
fUnH0/fOnQxXMBZ+7ZQCcdv9i5KPcbikqLLZxfxKo73fVuthCN1K66GUk3t5c2yayWMRmS8woR8X
UQrpp8QiGd3HZ2F8eyAWDxjYkTFOBJff+IiSYcrTIlQ23itBx5vdnC16gcYRrVyhTlH4fxr1Ab4n
2+IgC7pa3Jtr5BUV0gHxVROiJ99RWiqlSp+qSsMB7tbUAdp6mYGQLMIOZYRk/na7Cj4ER1zNElo5
v9p9E/GJy1B71lFtWLFjrPa5Ti8Xil640YcCBl3YihLv9M3l8kpAxEr1PXZwJY11tXl+d0LOMOqo
tq2hCclV+CpCWm0wZlB642mE/uVG2+dMWGvxJuWqpsU/LRNdmnjYpOAdmiOmBIF4Dxb20zbqa+lf
yYT2z25hZebGRP5wT/w56odIgZbFtp14ezXkBVwu3J+seqBzO9R71CY+IQyRep2Qq6oxifQzNKDt
MVHiVOmg/Wb22KNv7XrWn0YeoXWc3zKJ1uOMznqJmcZgFKlcQTNGQLOnYhbV8xGBy6x1szi6kSVG
oHeKBxhvcOPTi28rK86LH/0UzniaVxEP/oiLJX2E7u9u0v0lelUE9Ltvwz3415dAKId5iQS4w0n6
plLLzA42w8GqTd/zVzACJooyu/y1mWOb4D0TdLxZRRwe8GGBji0a6ojCVOwE1Pn+T0NibEBpQSv1
khN6LYvetRVlhsiBHWWqJcPkh/6rQMyeIepSEi6ZqCFCcP6XMa04EDcu+A5Jndal/3a/yRt5JFBP
ajWhanrVyW4yHDsSRjyayHUgbZTRPU7rwopwHQlN1aX/utKa2NyiiNVvJTmXIySO0Lhj6SpSIrxv
nAWClcyM6iZ0ZjGldnnlCU7zKTRd/b3qGmYjroqmpNFaEvy/zVzsfsNxzXOKACALS+vqUrnatSKy
ae1dyvRoPBQHA5cVyixbQoNy+43WuTRWqD9BMZjofViXGADWwmc0XS7bnfh3Fl1eHxUIzmlr5kaJ
4QGK+3/Q49Qm+DfPy1YGekJzXEnHewdN4ONHztJlQE8fTsQf0rVWZBXS/fAizFk7vr9jd8s7f8dE
4f7NhEetVNY2xBKneUt0aPo5OKU2Whcno0uCxQ8wyUiFCOvrPD0O1z30NKhxnJcspUq7mKmtR0So
/FaqY2sOjvjcxT5aI9G1OccUUPKvbEP2pY5WjW+KTkNIAsZNbjb+izRi/ivgtRCwvuDQ+meAka2b
Y6ijtj7gbC8r8Rq/9uMcogRK3rdte+TP+XgKuxVNA2POoDEzbUJyznd+/jfWaZT3VOY2uF4uZmCG
2vmuRsuLEfA2Myjflpeem5N6VYyfhsWYYPiDA648fXK7lojKqZ10pkFm45+4ByDvAFo0hugOsjO8
4PKf2QkWyRqVPyOZI093PN8GSbcPlUq8CNC1Vr5yTOSOCZSEdZw9b7CCDDrQO5bmQQnCeKkIQ5di
vQRwE/sRWuHK+PDb571z5aOLCeRFxJDnDo2k2B15A0At0CZHyD6nnliT6qgT4wB1jQZzi9D5T91y
ovDLEl9D5HDWKfO3Ye8XhfIel1CSB0ILCLEvNwnQC62X130lG30OAitQRSzfpGA422V3ajk7veOu
kk5cWMP8Tn3Md1qVuEnD4Ikqit6MnXg6LcLTg8s19h/5LSGFClVYhpiKnxa2PbBe/cfAd0DiONIf
y20b8AYaHAxBB4b7UB6+P6NMFrGZ8xqp1I1xHm5S+4iW46RP9+PSxpszfa3cXsQ3ohrxHsxX0w8M
VXX5vp2CP86gqbfgmW3f9sHGJKi5yvWXXtCPrONR+vD0oPc1RkPSD2ng0L1oCU8ursDQeml9+l+9
3zFADRioKeB1v03IvykkJxlj0fvZ2PlGFca8LRypnS2QLkAkwi6kdI5FovINEizsGqA6HO05CK8R
qm0ObffCb7MFrgQtvmNRJfLVNM5pra4a1/0V9zQX4/8DVG35Svmu0LzY4XUcayGsfQ2QW2tpkGdo
2IAXTeqmlHFoeSA5dxQsVfG/IYJVMHTTSKjP4qfj6YhnWYHBC7zIbHZr4SHnobcnAMvLo/6JR2Ir
pccna3Ee2+nFLeGSvb5DsDqR10y2DaIteqwaEgY98jdIDRVsH7ydnR8IT16jUyubaQwyOtkdYBUZ
MDoTmqFBysPEsKSjErNGNOGxPM8mc8pB2SOQTohFe/3CNEHrRhdkjoV7oP9UcK+RzzeMBi7f0mjC
p91VlT+70My3+RKH4mt7og1hArrWRyDO5uvekZg5WqvI9e/nWWyyOWe0RBeMSyhAA72obbevVM80
XPmELky5mQ2syK6hgErzDQSPSyaSdxk01nlcSB6IQj+bFFsbt71Ox+4iXHrdc1JQeBYSEaFt4Q6Y
fIsBMlMgjrukZvfJ5yUE1ZhZsFYBs4JQv26+dCemqSVBjJGRKqyl+IT6Mc+58cS+2XUBNmkqrLsQ
l8jkgJkwd374TwMzAXDMPm7QM/KXoXFLv9a3WxsrNtMPvtXr5R9lwaFrloRnBQeGGbTUrlzyprgo
AIDMoYjyw0MbCKCe10/AqjJFlx0CgRAH1x+zSHA0nZPwfpcWd4haJNbrTqpwS5b3AlnZiujeiAuW
jatmOyFkm3S+hqpYDuQl7r+T+1uWqTvzt9Rx9FpgACS5ITk1PcwONeFGBjJX7OaSJLyi+mlYckoE
btNEKmtMJq3kMwjxlJAvY7d1M7Dz9RLQTRsTPJeKgWBIx6e4/k3eOemSP3tu3zOiqeOXd5BZiFKD
4CZE2P4BqwdDA3x0xkZTwK6b770UWz0yS8JntxD8QBw8E6KTcouwoct19vrisbaEKZWb5aan0Z9d
Mt3A6nznHEO2q3l15B91FDa1YAbTihQq7PC/b/ZYbLyoZgz4a0tLGgKjbbrkHIr3M5Xs8SmSHVJS
MS/Iy5S7Tps7pHwaqfTO3NdfVCqtdECXZGahz7/+TyP+TmTIzUFXRdS/zBmuja5OZ6tg5jOKNZXO
X4bN6NQGDAAx7wy0d+JfLyd8jQgL7wtm/9nVh7EfKDl3OR6OMTnE14eLpHgNGanvRV+vj+fPPSe0
HQA655neL0aLoB49yQfUCn0hsSrn10sSBla3cDC2uA+k+J8FnuVGMZpNDojY4dhiT8BSK/DRpvzd
nLO+L8IizAoLQHwgDcnA+GxuFtyjcSlQTZHwMLTJ/cbxZNobuSwyj4H+cWS3w4jq7PyZEvmJl0TM
PqoH8NJliCjqkKa5t3YpRNiXpSBUz4bYQBHkWOO6hBzmwKjQ8M3npwWZEgk2EVheczgSM+7Xgvlp
NK0854nkuCIpWBloFX2DFBo4s3M3Sw+mJUfMIjqckvuv8DxhGUMVEVSCDc4u2sS1jU/GClMo7Mff
5l7mengClCYRTlUEFVUq7yCzkgxhWXLADu1PN9h6fIecWjULJoju7BA08FXaoVB559iM+oWn5cCT
0JWwDHz3GFuPxoZ97DgLSiLntXP0MeIfcimEFXKwkWJuufOWQi6SL9wX2lkuI9/3Y7b9WJNp1x4L
xHl8hPn14ICCoY4JbdeBpHWPFmqL5jGbU0dxVb2vT8UGzHeO4E5E54cjg9zBNWBVOb24tDyvcV4r
M7WG0lfBpGk9qFjrk6QEbY5pfPnu/xH0GE9eneUHheOuBo90iMMOExXp4FtNfS1vAMSj3VTrp0/p
MP8VA7vCCwUBek+M+YZHhgbnptUzsQF0VScalgb4wFXyfCb3fCM9fx+Ebx+fgJb8ECHiEv1XyfXY
Vxu4WyVT/nu/jw62MMln6oFB0zSI4GNW7R4aHIWRYrQC+ooyX7Vo9uwcxcIcQm7s8eA9GrVz2a+g
sjQpauztLSeGmIs8EitXg3cYX3EQ/KSSRypFvUYE9uXvZbH+XAhd1dMqSTdPX92u+FFjUpzlVBYR
DtWXqA9IbSuPLDyfiQKpVUAglTa3DdyOjykOpfLrnW6kptlQSc18k44imC5NhXmEZMEQvquEjo3j
hrsg+Lv8F29sjNWweicNkEe0kDs/wGSQSd7ERnqzDe1rpSfyuYRyp52d87reiOYa4riTF9xgIDvP
Nz40iFqWdnisIl3ODRczvM7qbjrpXUZigFd5F+KzUG3tJKyc8Til3SWbgMy/c2WXk4fQGVhOPN07
yFru5HqFfRiIiHAbYsz9A7C3v5GZ6dtLomUfMelkv+xOO82V0uFBuuA4DtD+bk3KbV2H6HPGJG08
fgOtPG95fEsqk7OxU4RqcASJA+nn+jq9NTuMWzJWvujm9G0flN7OdIiHJqQ8cHvDXtDFeKSB0kAL
xSSh8Nwoe3GWRb42Jj55ZLWUhe7W+pg3wtuop1If5Cudr3NLXXLnmKL2I8crNeLHMg1K/Od4AhcX
iEy8659kR+mTif2G6Kd9xz+1wNjjSHVXa+iXys6eoDnszCY7CPU6lo3VXtwb3WYufmCcEwNfJD0C
k4vD1HBWZ1b7vLv3rPJYDeTUJB4fbLBGL/kr877qoDl2/zbgYORMjSV63CDJgsayJ+8UvfzXYPOR
D8e82KS6N7oyIhVZ7lqjNrWILH2wWIb1jDkwpIZKg04lk842ahUpVuzHErGRoVSpH78SYtnZGVbu
yioCp7L7XmxI/y3kh9cHg9ki3w5jKtl+ck+FmVTYxVX7NG8F1p/xoonAZWy/bcpPC4JahWNui8jn
HvIvu19rE4D71VHVyHZfddLsmcGknnG9EWA16D9XrDjKxqsa2EGVSsj3mlazSycNqiNatiNhrIrt
+2sovoXYqryruposbxOgNonv26lBs38mKeR7z+7L8V9Cya3GThBipDa5Qif9jo0s4vSvH7K6nIR6
JVsNaO1sFiH6rLJrLVZ2TKVmsqtxrGtks5PL1LqYsYj7cyRqR9lblTE3JXrRuLyG7WlXiRMe6naQ
H50Zh472p33OS8iWXw3j+kRWb+hB6ibEJbbn+AEgwTZ21V3eMRw4xZpkqEtEp1ZdykgNUpJObzc1
ds0nk9U3XcAhCxtRuf40h4Eztmpohivs2Q1idGiXksCES8B0L2jVAoO38INqkpXubweMT/2bEYBo
jT8bUejFvwxlURpkHaQ0eLKl8tPSPyNTa6flgLZUtuau080ZvQDha7T1w9sYR7RB6RaGvfaJ4DrY
qyCHn/5EhD/wW4g4XyQCeg9wy6wQTmRvzUeGxIq8wk0vK/P2jUIohOhITCgXLXiyUe4Ivz7Qgzth
cL6tYNUCo0Je0jJ0JGTb2l9iNLZA6lf3UFexJxEX/wJG2h3euwdlBJxRt3fNVJ9ug/nH86k8jkZP
UThcQcQzzIZMy4Do5vBogepwK6usfuQYUhJYxLM6NIyk820rzkTkRJRe06NCV4nOtvep31pJcNSM
+adKHwHZFuDSqTdVPOAjLTwoJOJBR0NIQK+IVk/UI2bfbH16qLoOmIBwUDItZ76BGwwY4xLMppUV
TDj0Cqha4SsjDWtymMwtNrOVMxdW0NgYvD2lIpniDAiKXJK3ECg1BD1vBkuV9jXwV+lpSkFJ98/x
LTk6S+0b8YQ0Mgt70XZToOA70WkPOcVfVeUrL1Oogn5Q22RAWOsZ2+4sPf8ioXE/wp94j3ooKHCl
53M3M/ugSnyLt7OzjWL3lR0TQI3yqMnvLwJuHs+59KWJ4mXk8EpoykakgyxUqr5uIl/PUkLUuqpe
GmbCZED0baLMGV0u0tQDjcB4LtYRkRxasCQwRab8x0hVdJddpjNzNkDFN909m2tAB/iidR3gXJW9
OowxLmDFDn8Vw1vXjzfGmCYTjTD6jEFU+CXLrQe+0u2FusS/eoybbQEn4q9RNs2RWHpZNEDATEOR
kmcRq9yJPHlRScV4mbnw3W06IJldEq4yZfe6WZZGGfwMXSY32AzDf1TKo1SKBB6SHUXRmfo/k1uc
OeWR9B/9p8tHGNKzze+M+bRbi+CmZD6qDQpCR5jb/CDJ4Xfy/+x22FXgrftMHHIJyzg8zoYbpUV2
M20DadtWi0FfKVgiZXrFF0OrB0d3y1g7+Hvv9Da5+bt7omYvk29ms4v5zzUllfoBW48x1h7PdJJG
HokMepziqoElmrrMVBTS2zdvx5rrqo/RcHMfpoJ4xRHCCStc65amx9aGF/RZ13Eq+5rYVp9Hs3X8
JwBXxHSFcHIac6mFYmRGm5GuBuk0mv1LtYA/kz2FDvLNX/Kks9rHrSa4d2TyqdHHUe2X487G22nU
ee+2g9V3mx1k51TkMvY8qrxjykzF6XYdGYnrHRQuZ80obYg/Ga4MgtVnu/Vx4PnxPgqHW/nGAffN
iOrlKn3wLDdMWFv6GXD6GXylrYLpBrVa9HScXghn67/1DXsHFA7ri8sjyXUKsOPxhu7KRKPWG9Eb
dDoGFScLTujwkwGc+n6ewasRL2QlvOgokkwPoKoBamcLWKPh+L0lrZ0kcZ0nHZHvFh4PzioelkVQ
ZCRKADrq/N1Is46HEF/vang26ooYmCyuZcRZRk+ff/2jFfcx7epz8RcIR3bhvx7t73QtM1elfmP6
2q3nx7Z4fZ/aVYA3D0GAwqy2c+hJK6+EGaub94TszKYKAm1y44ZNgZ/tzzy6Mrg5noJ2NFoyLZNh
lgMI8IBYzSwMtHDpzdygLPTFHYXTFNtcY0Yst+A6+jQ2p9BIzwW6pdAGbF28R+GZXA4ueNV0Amm9
m7HOaS42WMvzLFr82HJAtHI56DHIH9Y2klg+Z+wpVdSnSBx7zRHM2Ynk2sqDZ3dK6YB2tCjI7WT9
MEXI/1e2iuOvVzkv8rxgv/LiDjk8+0ZG43IeKZgo64Qtwh25WYzHjsUb+Gcr9BsK1o0ZKO2hErcK
49IDu4m/wN00Duc+NttX9sOQH64mk/OX7ymxJNHkOKPV8Suy9c8qquB1Eh5IzZnZbgXatq+FpSDr
br80riQc76LwpMrKMI/JTHpMeWcsLSQTL6aQ5dKRVFRtcTvRDxEvdEiBXbZdws21KkExD+ibuWM5
j4ao1agE8YH1bgeVuE64n46Zqs3787bCu3Z2lEA8OID6hzsatPiA/83IqmbxVHZ2Y79uwQsDdSmN
JL6SQ4PQ8g+2NIq/ugpJYxclHr+cTRHD8zwqeokMaw6Jb7KnauAtKB2sVBiiKZAmW6xy6EfMttms
CNo26bGn2UiTLHX+ot5pguaHqGC34DSIDM0IJQo9wyBDCV3CJMYUCkE5fZzu5fiQiOEvg2OdPaEo
JcdiKrj92vN9heD8/KTnNQnewS/Ws4pAeYhfyZw9+w7kMSliXkr2Fot4TzMGPEXu+0dGYTACK9IB
SYhCSRSrc+zaaHozjxAStbItWyBzZwXoRzFYP9CqBEhAHgTMar7vE1XETM/BcEDxWzY82xtowPUI
3Nvyc/gUHyJkOWPgkp2EB1xpPjJwb09gNTLdyP5Bpg6fYcJIQ7NRFsuComvT4gXh4n2c9TLVc2qw
li2g1twp7uf65Wof3bKFcT3Xd3LmDETiozrluC7vXVsSsgKiRO+9DzdoiwS1r3gjN/cWGmnlj6bd
YUEWR+w6Ph/ZGrA28GYbYVoSikzTbhsKsScTafurvJ6G+68zWuf/nCCT2NX2Vkt4PvLn+p9fSPyA
V0CQvCYBt3vb1Fj/jCCNidkkA9i3Q8qKZZdWOBjJ6Cl8SgcWDlXjget+H1RqRVuTCQflABx4+nig
pGr9ZkpZQq0ktB296d4bYCwgOUdQgx3+Zt60V1uJqdEUOyt+rWIofnfNYddeHPKuWq2kzML/gFX1
h0+NhjPpk5Zh8XHhkIT5+CTWZbvcOv/ecR4TAsZFXVZ52AukypejDm6ZZY/odPT7EhPLj4BvV62M
/33SVMOPU+a/EQAgqzpdcOUEUvpF/wEiDMsrgbIi0bf1eo7tZRCP9Ct8UDdjASvuyT+h093WLZwA
ciiRWB6Q1ZPr5+wHOKHjpSihUuc7fSFnyZXGHsAohOcB0xHZPDoc0xDmBRWQvopBTe7l6Y2Vmdtj
XgbTVEZlMDZwYI7KNWzkutRLFqtY+yozzYx/kVEUa8uAEVc7zTWZYI6S+4uJ0ttbvsmkpV20A2/6
aEpGGq+dDQURrKdQVosVikbrJ9HrM6E2i1aJUYLcd2Fz2SOqs9rfrnhTRr4wtCoPgiGywwfId7/k
gClMAzC+4AIWFkbgnS+sSeRvVuXMIi/701IYJVuR8fhm71C6iEFyA4ABf+Q1ftHaZdttMTuwrVip
UtS9RUhmJRxQV+h1hKmpTa4klEnjWrwpkFGG+4cyNSYD0ba2L8J30STP0A+gK4/qMyfU/PHKX8be
u3SvdFibRkgjVNIuAtjkCvlRWdZC8wyjHGzQEIU0G5gVexOlHRjtK7Ao4QMALRsaw64GkRxRbjCg
1HWcVhPLSszHIJ7uD/rG3XGpPqPyGjbSHQCaqjSOZUSXHoGBe93zEvL+TDbnFW3otOnVfc+t5Uj3
ogFcenV53RXwGXV202f3Bi3A9wvzYQtLnP6lP6Zz8j2PPnh2eVMlxJYfwfTE+RNZd0A7zlDFpR0x
q70Kf8RjtijA+l8UyGqi4aahGorX7u6KjTDGIgO0QOr88Y7KJ/slIwHTkAZn6dYOee32oVItbQP8
5x6PAafpLDDCuiiFgyTtk+JWau9D1MeW0ZLsUMxjyEzbfPxA9ikC+zDRRH0qPKT9WLFigXH5uA2q
Pz7TntKyrhHXr0MygKevd5gCGSS/lr62+VzpnaJj/2rNACvB4QoynJi4kB20w1xwYcxdR95FDH4H
Ho2OR1nSyzCESXReM1g4EE6Mpr4XES57z7XbOohdZQIJQD+FMN1IfJ/Ka/jQx/XRpuiQGScBJS8s
6lv9n6h0KfFbTWyTAzXNn1SHOFG9092O8ckLHmGUkITO8QoHwQGMQ3AgP4eYwi8YuywDx5cvUczT
P6sXmd/EScaQ+HD65ZlquCI8RSRQ0mAAE7MRNC7wz7yW8ofFYXDJQiz437xh8X4gNPdzGp3VIi+a
+TaB3HK1dQSWL7IKrlQNycqTBHkMKkHV3hxmXsO4CetkyK3yAtBVhZVZA/W6N+VecWZ1QAAxPsTF
7g8412fRuQ9k35/G9iawqM3D4YYmFjF5vf8lKYXsfvxsA7hLrhD3nbkm6aBb7R1LARZLCNIc8ZYL
ybUiAbox4AAgUwDFQqO1T3e0PLWHtulynhxAHYdt3b8IgyKv9aPEz2z/JBWsQvNLGgMdV//T3YXF
CI2z9KvNXOoyEDmGRKI8RnTreyF5LVG86Z8nwT2KXJetotyGMdM3X7T7AkrUXWy3LGty+XTLU1gu
MrcKVEu0sfVo3O67UO0+0Y5IaNxTBkbX5sxx4zaLWHXNAhbYWWUAFLp+8KEtRrXH4C9+CBMF1U+1
Q1jl3kbqTU9bGkzA9+OMedp897Ry3DsxL1UY51knbn4dHwdzuFWw5Yi2xtJKvh6gba2uafoH797O
reEGQ14NiUNqoj5ooX7+9q8B+c7vlXsWBWeC7Ql3KlccFchtfLUTeSXs8KZ2nR25tl49t+RT9OH9
9eOrMw08XYMLSXixasbouXZxCE7rSr8+sKneKcZoWXoo5rd3Xih0uB1ro1dHBXbMC36p4otWfIWk
ChH17RtkaWFy+CvaCvGYixukYzs8/ZZJissa9Ui8dfL7gl0GjktlLfOU92egWJrR+LCiyonxQBb7
DempOp+shFlDYTrTpCno+toAVumwoMQDKQoFv0JoEP8c6TZvQ8EI6mC6HoVoYevTSkdIORQFFHKR
wB907iyJ1GJpZ0Vvc59FYwQ3M+4VV7gC7YixHE+2d3EPzNPUpHHqa4xC+2Z5twKSpofB/cZ1qQi2
6MGmBTIDDT/huImx/i2V3dVRZdO+29zOX04IxcxMf0r+BUFIsrY5vI0WFg8rhdIClKAc1e1Ux1fg
peWDrvYXz7ze3l0A7AO1TAg85s+sNT2MI86tsVnhjSVsds3obc+NOaTypZyfTGmBh/3U27UFj+2B
x5B1vfj+XontpL437gDdnnt5mLWCRR/M4YDLCsbFG+U8ylFbGqn0Bj2aGShOX7ye/IsbhCSUCeF1
83HSc83wdlS8H0I9n4QhPjykibrVOCdLBaOrK1ZWMh1AL3erg+2677rKaaOEJ0V8kXUPG306X8JS
pUNH5oKuvNOSkBO5YVjqfQV/4RpkfWXuNoLauytT/VdEOL35KUCfjvF8C9sUGdPXOQNJ6RuQtrtW
dmcJ+3o/KkQ5ltEkGcb6Q9v9O0/wq0mqJ8OUvAQ2Z1o8rDsRPebR1EHEFYxdi9WRUAukGAOB5j+g
Mr35UM62HtQWPsoZfJH5cshHI83SdEgPZRHwiyfiCrWFkeCw3Z1kWXLUEPpnAgmF6ZhnlSzmhVLx
JirKxYdwzw4s8M+1M9yO7KUruSmlxfCbGzvSI5SjGA/d2awMrzE7Bk+Nn8Z3FMqt9TIoDXnkvC0F
vIN899UFu1iihvv3BNwp+KHhUpioHrHXGGmxHHB+NdxZa3uI/0euRcjQkyw5BIzBpDkCfMwn1MgW
Eve473XIV21KQJ3APTGoZR5e0vg7X+R8pyUyENPBYH+CRAjMKQ9P+ZBKMhFM+VciQKgGhfRt99z2
vXUQVJ2yrPbgnBibP4lhfoH8jYLZ26jqIN8Zw+bHdjE1Kn8MGqg+XBp83dzmTFGJcc0rPsmoL3hr
97dX1NcBqHdHKpsNnad9WEJLLlEtUs1Jw8H4NfH89tmW8oYM/7ON9i4rcwASlhQSu128fEPYF1gJ
YFcfYIv5bLp2GBVhVQHkCVqO06oXx8Vh0tn4CM05tnj+x6JiY5ZHi/0ZUAkZ79J5nu3cVJY9g+nq
pHh3Pml+th7eJt+0lVTQRhjd5M9pBfsFOfXW5vBGiN1l39CVTjWUJ/+xhTpTZDMyt1FAirWin+M9
gIuKxvTsdyIzslTYO7MS+qv1cWY+Fv2LNY67mu3mtsl31z0MRLUPNJBQC8H96vgLvN+1rcuiSA1t
4D1TLWkjxAwUfnKY4wFTaw0EsNhrivQ2u30EjnAa8aNRcC6U2t3T8nrrLXA+jZxzzWyAOMiqDGQ/
3+6/mHgkcnZe9VMgiZRzlnGQ3cOnn4n0PnuBVRVd8OE1cA5Wv0BulrqjfxhpJBXYwMv+hieYhV5D
i44uWdYYvrGD/VAj7pgOouUfBnFsDRmgogdTZit+ydny+izRTQBBHJyvGCTsdXvM9+MU8ZzKicCN
dyLx3rzK0iV5UdNjcIKJiiIaoG/41vmwIVrrTcfpUTKFTyuL1m6CzetqOunWH8YHfg5VZr1WTh3Q
fwTZF5I32Gohzkb/FgBNjrCgktd3kYp0OqM14mdOCgtSZx8XjKkZlaZLClKniUkkWxNUiIMKlSgF
F8tntKiP0xgy4FUsWr+0sDBVpAg1DuIHDTm7I/LbR9eXHu6UsSGVme7liv9p7x3zMrAYQLRKpVef
vn4s/L4tU46k3VqQu0Kz0SWom8kzXeEiJ4WlZEGWg2ybVEvFjFk9IMhytSmzXKpS+9SMDaboPSp7
EpDD91rD3eh1VsoyKVpwl9N8NDKitc3WkTIx7QmKoCtx1IcUCZuQVkRXb2zYk5+s3Dpe3ATkQjTZ
2VItsgUX54kDV7NWTJuoXCT7fbI+e+HVQaM8eDYEQxF6mQSTunmdmdh9WP4zOn/96KftdeEIxGyh
v5yWEMK/nbFKUtrRJeTvb+YEARH43/XMybwTdZ9qDXFbiF43fgYKOZ6MoUS7BInMk8pqVtqIkris
VxH2bJAKOJaQDw0nNHAcnv+JqDRvZRA+DTxaI5rxQXhXWe2qEGnbWggSbVuy8i/yKIovmdSlzHDM
HJdJ5l0O91ef+aAXObTTYo4C/WBPB46g9G0S0lrq8MULIt8jFs0ZHxi4dpA3iAKOj2jHQsbYsUdq
FYuDc4IWgttVZRScVlQZDTVOmIuNob2zLavqrDE7cCHDtzgPpB9AgitCHrKpq3RGEzUqufAkRXP+
i5SZCmhvu0CiOFBcTUm8jkuq0DpTtSGfERjApfdqtkp2BcrK0kM4FJtXUvXys1upiN/olJhdXmmJ
fqxSlff5XF66K9pH6LYvWGBSJBITd5CsZCi8gnoJj5X6Nl64/DbgFqHpxGZdjiVjyHk6+K83XhHg
DCroVhVt2q7Kzk9ImBJyGlMWA49d1HhgjETwdOn5ivbiM2fOXUFgy9k3EKgM2XGlpdDA4dMqB8Kf
RqxmQKQTO+6Xt8NNDNN2RGOKc06t4E71bJU1INuRmvbszTrL/esqlzoK/LZU/asV7ZYVN+qK/WPy
FLyClUs+l7k7M12GKxOBXXbfjZpm7c83EuKcCYnlXZiduQk73AvNYx/uGWoByGh+20qlj8M67wgc
jvCwB11iNTZ6/lVVEnADJI6IDHmR4yHr2pUVRaa3BgZDhw0Y2JpIhS7IJuzx1FcvBv7XsUSee7dZ
4+i4gPxuSJ25PTnE5CRA7h7yvoD0Qh0NubX7Me1cYWTn7XQagJY5Af4XD7NBX8lF8HhDTwrzZDSv
bbQc6QA06CoodEOjCZqeF4Q2C/JWXUnIKF4cScENxIDUkgi40jLDo3s95JGIjo+q4Luj/JfaPsQw
FZrRVWXK6s10TpHX2rt9UTAMdesVxXqgElZtZJw5ra81fnsiClsSRcT2nZWDot8JES/4nDPT7EqQ
cKz6WXxtDwKPkex1phtud5mEzVMdvuRs7Rkl8KNyud18nCxBdixnNEFQ1uVjRtOojyWO3fEyWXi9
OtEpaws1IG2lDVwFLBqYKe76I65ZD+33GNp2e6IhRfKy9VQHOFAat4JVfLh8ztis1xRWvHtRg7ey
CFo8/bJD+ezeo/2qL4ezX9OOsBqspAOCoF8uIiUCMdfV9Egj1+peZyI2VfYOqXshyvfmldeAVPNl
o1naTpgTlSUMiqAncOpQfKN9hMURmAAyifyOG/6iv9xZhc3ENvV0ihTVtAP1THq32gz/8W9GX+yf
1arpOj2ME0EMe+TEK0sT3lf5nLXv2G62DklmtjqZ69U3efcYl//sTJf8nMG5sz45WQW9T+SNShVA
AAPbCd+XQMqdu8cVZ8BYmJWfkISujKXAB5y+tSfoWKT3fweTaDtcXu4xdj4XRpUrqlnb5/o1pj99
n/iwQFV60uJ9w4rzQZ7j3vPxKe/H+rh6bnhtnsQxyFPvjmlqKeqRAABFjlVNBJNiwezds9WdiLjm
peIMddTwW7Y8KUDVkQH0J2BDHVxuGjJk7HCSpagEn/veyhtjC29Y85WA7xvYHQqxdeYoe7N7j+Sn
/KvA/yfaoUk9NKXf76u7WlLd+u+vnHw00g/y3/lc5YYuHGIJJspWUt8p/Kr2iessrEJWwn5f8fol
kJpR3b3z04NoeikvUJzMtvBAkPgt6Hcjz8UVDORIL+XDxr1KafRny6h2lBq6FdK2IQjvebExSKaR
yaFSfz9YZ25edN+oxd9KDA6VwK03YFoUqTXpaHzrWjqTYJI4u4T5a+jA8wv1K1hm+FQ2BU8lM1IQ
MbHvAdvV/9VeWeioipRBaQD8KnR3qGOUM33wo+I8nMAmhQioNYYnCDbAB1O+tA1kSbaN2yDfgSoU
yEszNNQGPW+boCRkYViYGHy+5CqBL2k8vxqo61gdM9/O6bzWy4My6Y8zl/475S3YpC77Z8x5kL4x
nyOS5jD2rwXVFFY75mikmz0f4HwK0Kfgz9E4EXlhcALM23TXZs+T+6GpowO2CQq3tDldB1qbDZW7
DQKLfrhyihfN1dZYgwriEOGMPS8VaUJVe0SFWTeQCPoEYIbSSIGjAiPds9xeWr1jjUf1xCwo0QMB
12N3mB8ZuIuVy0l9r60rRi2OMb8ke9Fd6vAYtt85vLEdl7ZaZopBsX3/EBPsF1gjOVqMDtxiYoQR
zA+Ca0NMOwDA4CfJZGsGNK3lgv1lFdTL2kGquSZenIsHmUhOdEpMEXM1kJocl43Hf5qOehnx+HFN
SVnTHVDSLKu0OIp2PifMHPkpPQnmM6D1nHBDKoASlAb2JtDMl8PLuP8PhgQD9HCtXE8YM1NEOOVE
Rdqlh34HaIkjNO6iv9mHs6T7GCUNn24LDSsVAbAd1OXY8Hv6jqaiyKL3V6RkS3Owdv9gKOpwCzOc
dR5lLiP9C8CG1UfRrhNkTWqY6dRxRsEc6lako5lnKQ9zVEoSe6mKvijXFPgaaw85tNDHa9nZqvZE
NTFDprhSj2MSGUJO3Shz7595e7WDS0aKUQ+1NntIvukbAWfDnU2UfrbqUgR2am2G7eqqgQ0orS88
OfuUlhi8w8qhxgIZwID8VwCIPePjPnLvxpXmmmmxaxBz+Kj6o5PWBSnye/7lnmzRMakoIcHZR2gZ
AFRqgIBeOjs9qYtBT1t9+2Zjd87q3ymRnwmS3zprg96cmClmLvOxPhScyD5I2EfMjGE9tIHEgwyK
fWiDXTeAZdzyi+oCRvLojuSubBKhl5ebnj6lBfWr72IO9ls6ZYnpQ/KA7vpRMNbMLhbCNcygaYug
gsvMpZ1pv9GVsw9L4oqA0ZMrEYD2+eYdcEFZ6wNeCqR/IilHPAV/gRprGU4JxLhjpbd+UQoH2T48
aY/ZlP78UwEN+4mVAORm6UDa2Fd5Aw6p4j9apgFpQ6xsKLb5NH4ciZyLBhqyLqaW3SqnU2jYFk3d
6orTST2r7H2B3kMx8MZ0LS1KBSFet/kYHoaWkH6Ds6jTycEcM9VfBP/a6BkJ6+IyKBzopjDQpCun
1dx0DS9TLcPQuvnXlz0k/XsAKUKGydwoJskwBzTjD+LdvWjIrrI7NS0jtVL64eA8j3HjFb3g51dw
3JuHhxXKlCFJe9GfZxKsFoxcGpXRr3ckXfY0GfH4txuwJ59xRKr/9Xw58i4dRaqJIiYo3gZiq2bN
dX6B7tdQv+l1qiccWeTJaKNT+lvJxHlK5l+lILmxxpUak8bywVWFbUu9H647YdqiQIBQyoiA5oaD
LSpNg1cOWWU2qWF0lk9JoOQWHB8AaHPzaOr5+DEK6vTXDtPorA6qltcrf6KMo3a9wrflTB8OyNN0
BuaCvBo3yGeixaDD/MMqi7d8qX9Zi5bdRxB8nOj6OcOm+VUCpAexmy0bdCuMtr4puzcQLor1E1uk
CNHxi27y71hIwD7K5i6CJW9jbb0ZI2suzpzuVaL/lW6un53ni+DG0LLs3nFWXgvyM2tLd7PkuWSy
UGndCQi/PR7LXK+iGtROGiGuJqJ3OgAgJmktVZdv8h4mmScExNOuiqef83T1PsiD8vytj6F1y4VB
OdpVIbW4E+H3ZND4iaD+Ok4ecnjc/SDxEgp7LbpP4yyL4NSHeraqopanGoEfGFjM7UE++vu0lMPs
1IIOqYaHQCE5n3LvLTFk7FSfNucelCc+JFQINuf9AOvDE0/iRFa2CgdEzcQUjAIzApWnVm+LdAg3
swZDuWl0Am7wuKaZ4htBbMu034ZFoZ5Lfz3QCEoaps3FqkA+BML0UWeuzBOWimypmloyEhalYFsS
T1rsNYimBFDMZ1XIBx/TenbjNiLemoq2+j6YVttdrnbfp4KuqJkAx0bQmAUSHxMe6T3Oro+8KaMG
bwN/fFCEuVdCk0C7eoHRjxH1pAU3XNA/zFUklg4RWpNLRWmOLRYIZAX37oVgELLGBzBr5XyuGB/0
2xsW/X1tiHYi8/t+kLEDupCLMBL5I9TMKi9rauUjwvIiDsRuCNz1iJWarVOPzbi4EZU8NCk4iVUc
M55FL8NnjXsTHSqW+7VHLfYGAjCzOX0dluQ6YZ74S+JK5yHdRecFQ7mmemyD72KoVKZr/6+Jjhud
IBZdfoa1JMiYiqgYzE1fRynZb79/1DwseupPesCmSeG+4CJO6Un25V75OMz1AWXDtbeSAtmsA46q
AsajnZZC9WhNAVgvuYSqQ2uLGwoVlbZwY+sCo+Wg8UFhQaWNWxuKkOSFyN/Y6A8rjK1uiTidCnYO
SEVud4i4uReYjltuGHOnl4t6Tw5kwUzcnVWxjZm5J5/LNeayuLFsdYEso03WhO9bBzfl2k6o1kMm
1354n66tbe0aGyJ+nYz1YuiJ5lmo+rgMWgqMnlUovD06OacFal00ltDHofDPlux4TrOsCwbgujc5
T9/tAk1i7HE/Zq9A7mLQdqj4YBKhQRhEG4lzCh2KEJKxiruteSuhzBJ0/vhkWXDp75+qoApNP0an
k4TuGaTPwpgn+jFWGU8uRZLKrb/AMfdaEn5fxEe9lS88ONJWb1R+LGtDRMafq6Nnt+PiX8z9DdMn
a8CRSpwAp1B1/NCbpjWHwG0+P2VBvtKqOwDCIAuvGR4tqrR4RTn7B6Xz5QIeNJ66vC7TOZXvfu9i
cSopgaavz0XDOx4UAM+2CSkJLTAlhkJTxyxOGl/e8NSlRPqqZyZzwjsWl9+QVbf6W8ZD5iWKQIEt
KX8NLTz3TDjxr8sjjNg/MQcUPzjU2t30Kdrihqvjne91bcmQARqgR+DzhuvsOP4e21sg9sYFpPw+
ZqUMMVPrdbvG+oyrb12/NLus8yJyCkn/RQSVNgLoCSvKyhWySXlu+zCa7AFkzofYnYzP1Fce6y1V
SBaPx93J7Tm3omcC4HIDhWTgmWskAvsfl3qdQokqEWZMJk4k2aMt0J+t8DzL/GNhBRkcow7sYstF
Vf/bWgc7xtYadbK7Phzd/psWp4iFsZ3Od+YgQIOskuLG5WGyVtSkJrIwajpMVe9Fku1nD52Wlb9B
sN7YsTh/FsdJkyCcqNI6jYjeNBO+eKNZ8Y2jCS/i9fnrgfoo8/XlfT0cwECi2wTVE/vz8d8uTnvq
9xS7zSZNAHI05AtC5TIx5HC0Sq+lzfqy2cj1QOs6RX8kRqYIzOpQh4xl7qhMYkt9+k645S8nRvnk
t85HTITIT55zx8MOWn8tNSqb0yUo8frUtXRKPAKAeyl++arBMV91Wux257sDU82hbSXadeV9isXs
zU0ocG3wc2JZlx5pCWeKIHLMqEUXcgjeMreDxjkYE/b8uagpAbgne6ut9cUrqNyjBsZfl0cBZMCr
4zufNBYvhJz1nPFdds6qorX7kwXPmqZU0DFTrdVIESZFkH4TKyt2iVoK40d4gfBis6SjPPV1lcbA
UKMRpbLmlSaQgFeBp5rD/6/j1oiUnuqRsVY0nrvnEvWsUlyw44+mvkMFPXOPRtG0SaeDMeoWbeCG
ahZNRE3xfQXEDC0YFAJ8PvxWZ+Ms9/4rXqjo3/OwGhAjiXKp7tuxBXIx+PuvnYoQNA6B9lmgkiyF
lMPomO+aPutLdBaMJ64ZFig7kBj+Zua21VR73Zgq6r1jC3mvCKFaVujl4rGnF42q1CIsfHkDJZpV
NJ2uDG0Eu0jVxpf9s7D9nilIo9UnIednuT/UASW/yYuoQtd1mASiHELN9xpttPkOcXGhxoqZVZpM
+WwQ65wW6bM9VlY2vvwmFzfHCKuG09oAzbbCRp59WAgF/UeHbtdobo/2J+j/9btw9Tp6G9iZpMvr
q/cn3RNsMDtjUHh+W5CwVQiHRPiA1blX2aCdmkfiuAPp0cAzZj4Nd77Y+SyA5ueZP4VyvsVZ1O/Q
S+engnC/L6ophGCzaEBGnkDFcleqLrR0Zx9srbNvO4q60i/gIpGzAlBhch8ODEK+owA+IRa0c3kE
tK0OpqNtQSbFs79gEcFLA5uWvYmSUu9ER/1bsltCWh10tvocT5mNB46ct64bWd4OlBQa1so+S+aZ
rBlVgcF3MNOucMrAja0YTf6gidabTKGmYYHveodXWoafxwZaLR3SQHGFoii+OvG9mnpKmaswnZDe
bXF+DaBL4HYo7mP9kcPJJAgvA6/iIIGM00OrvUS7UTaTwKUAEx3KcWydfMrLq2/ZRI642VJdJOBO
Qy4ZVsXTYsTLHH/XeogEBI3bIUI1KpTXAPeWJbVEuDOhnlPAIZM+qX8vcd9GFTD9IFcXupM5h1Co
XdPTtMimYHqw9fzSqNi307a6WvsYK0HMJeyu606TiatvEfFzb/1LvnhzSxpJpIVzUPXnheVImuc3
DOAekY9uJ1X1dtsQZe/WscZR7ZXpppsSTsLjlFr4RJmudrBZOammSL21e6AbiXMb2j9htVnlFaEG
13g/3QH8M/2UX1Yx+55G5JJo7zPczqFrp4QYETn/HI0odaMviaoxiYuf63qJO7QzEQPZsdFMBB3H
ZCFsp72m0IWZibrsvxYgIQOwEX+zje+ns+ZNYAcbIxhUbo7uheMmRkm9LZU3zBkW/ioGjcsvMmEe
mkfsMfl9KrVoBwLClwnQCCuI3XeFymLWpbDFxV92vcW0kGoJJgiXSQRklfLzdbfEMfdRKfJzxuBY
OYzItoYBdxAyScioxKcVyzc5A6CSPFhapBRDQzhSy4pBGuf8rxNI6ZblvcFyX7bDP81q3HuuCLU1
i5iE6lt9o8pp6X9JvoraH1d+0Dvch1bhNdKZcH9Azhc+CTYOX/jcNgfLEHttzQ1UfeppFDl1inXZ
4MedqS3MX1c953UmryucM1AXhBq94fawsmYJh+Z62wqqsHjGjTFuSjm5wbST7kcFv9neX6RIv+nZ
tSSNuqhZmNqEtAEIpzIlmnlvzWzub1Cz+fYnMFnyAFDg46BQXaFeNFE/uVZEQd4Pf2fkvD2Y41oN
A6b0GaDlpbP03xRbwdD6a5Lao2ZUxfrjRBsHdDSYUoW7/0rbg9+nFBeOg7ylB1iMj2uOtmYbbN5V
crZGI9/OvgribNJszJ3NN583YeJoXl55KLHWDKvAc35OACfKebRT+TblNf6hCy+GngXco6iVgcWG
HMPmkMDkIY1uW3QklFxkT303HOamKW+9Bxpask7TaKi1NBQab/DIJw2IOPnVmRxWAHdLAbMDO8oA
yJJ3rWzzKfMioxuReNeENuOjN+PFEV8b4LSGAnG6CyPx9lPtDQdr2HJnmY9Hm4Lb3aYRIRXo1DyW
VkT62K6USxykDnmUec//sITpsCUhWFmdj/yZXhAjKOReLc17Mx+YmyVfdXgmsTuLnWefgSkBLyKb
grFskQ0oq1ARC+F+25B2kOnOHfkX4b4QZvq9XiF5Oo6s/h2baL27zjMPC3/BpkCdoXTp4tBdYetz
0FxDs0hvb8yY5xOFhZ1TQ/Aokbw7D3jYhQbW467z2Io1zwsWRfUtKCSXPNpTB85dTGR5V50YOfql
ELLOTlblTKxIEpHAS8/RSZ2JuMDxNueO6pFUWr/DuT5IIzKfkccL7SZ5/lmxYfufjflNmlSumwjX
7Ndcg9C0JwZnG13HtGHfbG8aNLPRLyxmVS9e2XytM4Vg2UW5mzZy2H0kpZEhAG3SZW+Q2N5Z1a0e
uoniI+UaiAlSHXGFGeQnW2Hi67QawdF1xWGVpGNuO4rZ2kjXW/PF8U1Rl9Rws45fIWvmULu+yxtm
ddzxpMO0SyfuRefiOe/3ydQCwz+rPdXBP7an03GqyvRgRY9m4ehigIVL3LGlKksWCdhOPaOIDJbb
qQzbTB+hIuZy2scJBxl6ay74SUcRb0CGqjYWOVaghmDHib+wnwBM6wrv0dA+NsF3pLH4ZNICFV5S
niDxb9rdkGC7V497O12S2YP/hmxmP7rlPNy2HWbwL9VAQYtJOrFc2WrPmvi0iZWbPbhChljVrIyt
N6aS6j8fudT9fOlDTkTaFQ4UhJS2HszjiKgZ71z7mJya+PF1QHINjpaBap7oFy4DkfGmGFi4Yem3
b9WRAAuRfDoeJ7jxFWp5ACGWdT4qRDnHR/dzAF1IXN8p1uoYYmBUjwL7+0vzRWqgP67lWRlBOzyc
8t1JILI5WvOY53JRHyHES1qCB84NgMW2ot99ugdcnS9Nu9u1waoWA5WwlTRvhwxUeqX3OQ3/zePt
irXZt0xAAyrZbuQkED/8qL47RT8/MGon1+o2H6oJu4AtJMc1QMQBfAGlxU2vJJvkqzKwqZ8KbjTz
enyWWDLZltKJBBKomXrh3yXS8DSiJfHPQnhnyK1qEkSKvD22CvdRplEDlkZ94jPLVxN5tHrf//mS
REVKoyy1Asd4o2Ifgf7I/mE14iIpu+/OHNg1/CQrQFEn3Vpguf/WpK1M4VcnTD/C1dEVx08/Xdim
W7AD+s9epPmuX5cQ1wSeBOAl5Cud3HDnLKlTNvJ7kvoDmlK976SHqYIHc915dzQBDOKHimGcBRbT
GnRshLq2gxqw6WaVgG4SyYT72af0TIZ957PZ6d4szwTeIKkNRZ7kAj6hcZOPFBbfT3ZwHmX3gDJS
mZgkf51civV9uYpZnwuq/AEekYzXYs3ge8FIlOvKXPgHUHVbbNBgBTBGPWeHWANDPbERdoKvtofO
Hk3/psZ5CqBXLtI2mpbBRU0KqtG0zYAg7qYYqwVQTrd/m1Qxw4VXKxluvefK0x6By2gXuIOPHii3
2Az6W4i2VwCWqinPPUghOSKmkfZoR+dL1zy/rEzhviDaBLW6qAyElO+XDfM9dG7CNyOl9+anP2x+
WDtKGIj8aC1dU65g9kVh38hACYshNTxPeE3bNw82sA9tESozdGxspMmA5wTqzjqu/E+52jf3toKN
aWfaPtbD7LjvXIqBTxa59IIvTIjMNiX9qXqGvCYZWQmrmhrvlXlxtT7G98/1XuXoMD1emoGCnv1/
vGo0QX4Wzs9TbPGF/X25T4RS4p2i88nlk1e7y4ncYpkkjyOG9/V1af+ecCX9CRm0/Fbj3waoZ5rm
2BtUEQ4m/Xt+2UZq19weNOCFsq0Ze1MOIKzeMRKj5HS+2JjBXniL5oa3SNjvJpvDo0caFJEpjBKF
V/c6QZ3kZHE60T7hD+QnUW5C2XMF+mpaZ/61N82EJA/LWcBkBCvYLbk4yRceqp/VoocTFf1SNZ2U
ziyjpQrA80gvbH0y1fTO4qvb8pvSz3wVeR+DSnI3HynbhZeCElVlWIjNvqeUQyEk0s1ovbZOBcY5
SLnSSuWVcD5bBDSCWF5Kc+Wu1JT1ecTyPaz6GvsWQZV9A4z61vivxOt28yAycQiu+Nad+dNwE9Yc
8GLPA5HeiKw6a9nml7ObJwOX/6FqkniQcv0Oo/uZsqL6JJglMXZEz/C11gCXBiCm8t58z1n79ipG
3iHyGg622XHHVYPa9gHYyU5+OHgubN7TDo1OWl0QInEFsfffciF5mXmzOLr5yHEM7TlewRFv8grS
qm85LPYWQtgh/pN9+wK0Z9csHSDFOq1Au7ad1p0j/h4ztotf5Uk+BLuXGAYKbgbRnUWbmJtQnOYv
cjUsgzyEzgfaLN5Y+0+fd1uKns7SeYFvG7ald6O4PbMIatAkOSpfErIeCybvkSVtrzs9NscYYMsi
Kt2JDHaIYuF82hfSNQf9X9pvofmnqzD3rnvcMD/FBrdl1hX0W0wRVIAhltuxqX3xExDFMXHhBvhm
LPu2TP5V9F2e9k8P8z2ISGnCzT0QnFDkLvhaIkkMSDOTAIvF+PhGKpCwk+uu79AYvAgGscJzV7wN
xO+3KfcqCG3Eqkk63htmdYkxJk2H/O6BbOTAT6pXldDecVC0q4ODu3hOMjk45oTzIEs8Qb91ee4D
e0+yAojKMfxUY1WGtoDfz2C+ZizupDskTr6h3dFrLH/cE8Aov8j9mmAMAKxbhHTU63Z1HjwpCtz8
/h0Mkhtk41jfmBd3OpBiYH1WHvun9b7v14jNCuPs2jjAlF/OolnhCL/to/mT4Hz3bqlS24Xct1Lb
rw/dePsOgORfZkzLayszqc3kYQZp8wh3l5F9fKAwNdaY9guoozxHYTGy0c/BafVSrf2HoC+pvhzf
djk4qp96kRng6LbrvwfPyTsRSo/pE0Edf6p+8kSTCnAbClZMAW21HZastQjK66H54cYRK+PXRfhM
KeWu5WgdYNv/IAGG6D/BiAl7ja0mxgSvTXVX9WBOWnC7TBLG/a/q50ZJLN9S2sAKe0Na5jmhKn4e
E5Olo5spGQaMZ3TJOFZA/SqcgGCmb74oft6lmFTui+NzWDgqphmElR2YRt+SCsYSmndOTsKokR0X
JVMIRjWxeVhzp23LeHcxKfK1qiKZRS5Lxw1P8YYEYLVV7ctbKch4DP+624lwpuk8AxFOzCEX7itD
aYFz4ajA5Z8dpDt4TyxMnPwBntMoGPvObU1JQd8pgDUOFvbej8rMlijerd1Ie6jmJTNMv3mQt6PD
AXh0qqUYmabnPJFPHcInYuk0aUVAvdSIL4f/CP13jIXj8f+eNUU7CS6lhZgWOsY+ZwpyKIr+3YWf
6WswgNJTF1Wo0QZ6BI5Tr02/du2tqmhkUSNT3cHfMBT4TS/bXGIcQXGLgjzlvo/nkJZ0TFjp1OqZ
OIXJlFec0doDHEkeIMrm6oPx/CJa36sxSE1RiZCg7YF901+4c1BLueudh6sF4lzh3zTjXKRcz/Av
OeTN7KQUDUCCGTElf0SnyO/cH83m33WGZhJSF6vQ3O/DGJnGUAkUl0D8UhUkm3S0HfeKtEBGSikD
DmCoQfu3mYnkZYnjYMU92/bW/dOO5Z+sOuFoSRvgR9yvHg5p6g/MT8uH+jDIOmKN9luKlVkpFQkj
GaDtqy5B8aefqYfamLLrsLIXEKzzi9PWD27hWZCMwTOepeAfTVxeCsMQq1hHpKBg1I35FalNvDZp
RCb+tZMgN3cxtqNv2prFJpiRKyRST+Ur5VhDf8fzYkF6BeOLBW14TLfydHPn1//2j7YjtEMHqcqC
6lA7AXwzU85+jVXMm38hsmE9sSBidY2V/0nHND8s9iK3IdPcr6R5CvSYVuXeVDEGjHsaUUTS02QE
B30zzMdE+JJ1ZxrzSKguxb4PrkGoVtE+PkixAjN8Sf57VQqPnN2Nx2O8k5YGqTvhWLYCAUOmwdXy
p274y4OYvnDQJRRS316IKx+mIvxIRiWXKLJHPSa/LU+A+5DVlk8LRwK/zjpHxEdjQk9R3avMHHzx
ueYiCJmVVFHAkv4z+CMF2r80N1ubPGg1CqqZXQr0kkoZCnQIRPTV54flifrlmxGGBJm9HTlz7LBw
PT98zB3W6L8yk8DtCkl+1jfLI7cUtwjxIqbDeanC7WMZYx9/sEFcn7pt59fUkNjE9yOWBcna47do
kz749HD9KiQ5vaL9E5k+DHFSPWpSyJsh/a3OVuqKx6LpsP9VRZeVr4qO6J2qVCA4ADDdRXZn/3a5
Lyno6YU1S20tyXCtgjHLkeMMmhdaKMoOQU1uE6hMIj12Z3S8axcAVccFh/0s+h1w9pVsvRMZZDg3
apvaVZr28vbkgw9o7tk+CvfX66sSbY7PIjLJjIt88Eg+SbbWXBFeLfEYuXBM6jboZQ4aWKQ+TiZQ
gCI17XSzoiHR6k6J82PKjUOkMRuKqFyHpwwM4jTylOhuWw8WbN/urcHTT1MjNr3tTIczUYhMai4D
+rzv93GHEhAhof1hhCI6dMhC3EEAOG+uvhDY1k+yuQ/mNjv9Y/gMcIS+FcPk0b9KRk3JrMM3tx+y
WzNnXWrxudYbjMB14Vpr7gksGH6c8ytRU2BXd4d+SFeQwSIW/N6PKTFBUQ7t3J5k1AQkv/4WigsW
06yX1q7bUIdtR4BMZg9P0a7B88xjzg8TjbLMmsxK9/Iz9EGSBl1GCpni7MbdpiOWqOQql8TYJARC
PWI+QyMF6A4Zwv2w8Dtb+jFUD0cBViIUuvUCh8NCePoTDkKp8yk9zFggYYM/HU7Cf8dNMC5bYGrc
toj65EGjzwpJ/91IiZuYsKhjIEQ6rVDQStU5WL9KKIJEs3SDlxGcqkLpgz2DYXrc0lkZL5fXFSGv
jIh5rqXNd9iS1n/g2OK2vHYeg7AtlS9sW5vLvPblbIr5Q0tCXAXrE8ZAJDzaTh85TCJfSuC/BbtA
dvggSvNtLeWqg+m1hGxwo+lxPbjPcVrFs6MkrJH0pgyOSFfx0Z8TIag25HSyoN1lcCjiREMkZRI2
E+pbP5vdVUEjanjeSeYn6PP3CqWGpBnW1vaGUbbxyP0yS3tLZDAkzilTqhMJXCwK3e6k1uzsnofX
URCRGvERt1iIdltxc4WO++AB647TtfuCZcGEXc3prM0YDtMt0Y9LtxBgZ+ZK2AxmmHB62Ep3EW9U
V5NMa1wSbc3DqdZa0lHWLYSiDUDOvWU1H+PtqwaIdSMMhrHVFLG9Sag8IbRLsXZK5O5aYhH/lxPg
Xwd9edF23o0k7mWnns40h6AhMNtUjsWzjLrofT2Z8BkUz4PbwBC1FJ471pfHIkf9hXjwv3xF5lLe
bf2auz1QdXOjtf0zeUrysISA3Vsknf3sX24lTBGzHdnGRGZYQo0dCh0adJLOZfAfmUn8tLVaJUFe
Qb9v1wws1CFlgGXTVph3XGioK6UmGUOKnnp9m6LTElSA0B6nqfiBYbezg7+M9aj5oVL9AydZl/ir
0a4l6KDKaTB1QD3cfxnpzveSEY7iC3hRBze+9GF/V+VT8qcrvNK28lQB9Nw/wgsnJ+Z6M7R90rzJ
GCnT5/So08cWPMxhuxyR0D7vUBSqsE+pH7/XZeykJl6n6RVxAXfTFWBAtUl3D97hmQa/InXvFVOV
M5rzHCPqC8H8IgFAMZh4ANsQvbZ9XeHZY1uTxmJ/R6FAdplSa4FiIkL7sny6mi0WOn0xA9mMLt5S
5GfNceRnNdPWtUKgM2DfmnEsqJ4xrUbhUq6Mq/BspRL95E10JteX/HDqBHO8HeD8sOlzPY4Jf70r
PYde4AAMY4tEdpy7BKcX9niHBtspPLBaok5lz+nvLbDtd662CM0xlOFpNU7Ziy60hNhnsfmYmFYv
Auas2Q4ExydahAmI5VxYKGG71QfNasK1Y/d0FUsmAhA857MrViEk2MNjuXgl/lMOd/hQ88QKAvVK
kasn+H+gxSFP6O88JTzuga2GZ25bJfHa9R1CZMX40N3XRHnBytNSHxkk3b04gDngz2iIebOq2uKZ
jjKFSG6vWhpkZfLVJ0HO4eGQEO1snf5UxlY0s3G9WvCf7GpVuXBx9zIglY9kSh+tIz8fYUVENvNZ
RtTiSouCj0vZBNxfOnD6pbdUxOnHDwQdXzpkfmok0gLkO/x/QZ+2Ll6wu2GggAIy6n6Z5zh/Unwo
U16YGdRLCsnuAiu8DRnsA4pue3gNt5T8QOXAi3Xikju2qnI0PbZqMGbcfDOMpjC3/pmWkYVBYFg2
3ave9ysPZL1oBvJrTerMfc6pz46NX41Qela5S57bRwepjCaJSlpvUx11KH1BGwlCG5CXc99UnT+7
Dopq52IurkEe9X3/GmpQCVktb+B2W06S0MJD1vHG3MPNyp9/Z6o9J/7oV/99q33Pr4AN5nn9zF9+
0OfQ0oRuNMM3SiWbmFs+CEiCk8jQsCHWeqb/n3ba1w92SD9wy3UNyL/kM2EbapfvwqfjsrSjyRzT
DETIjemWgJsTOUL/svhc1vW1zTlShrQUTFrJazUswDL9Etd8Tc3EJEAU8JCpDeeyXd0XYU05AtAp
urLVTmkl4ceFps+UtZfFa6KHxFPXiM8jB6GZ50lh1XeIHhJToCEXy436QeOJlYVDjxlTSKw87jM5
xBEZ+Q77vG6LDsH8IaCV51Y35+2h3MMdTmJDLleseGH6mTTYKCtZHxTiq+ttjczqKLvOCsrlbkU1
QKw7ViBwRLj3UkGtRoFzQdzOzCLqOPSKpu0ivdz53U4n7CqoSnJOmxBJ+CzKfSDssh6SJNGqX0uY
nAGCZTj6X8+Zx6z9Rqz9i0uC5vqRTNBGaiyOHl4sQ37IVfh75nku9N2oFS2z8Jvl4Eg9HHONgyWy
tizeLWhDc+Y/8C/QnAxhIEZ5ylyhCEHmb0HJp3kS9yqJgqIKI1rr5jAe4QnRWhx/AWPCocPqZnKp
Be5VH6mLFECfDWv5Z10Rsb0TZ7NvnJLLAqlAKsLUm40ohzZblLyfYxwxoPsvg8f885ojq+BSR3t8
6RTsOpgeDXI9qcmr/wsd+5Kc4Xx9k9nkLI6JCezRIX1dCE8Llzd+deCitgRVIK3IPa0sZoVz7jjd
91ZbCqqgy4f03afnFgj5VGu22Iy8QWrvuJd9id17Y7AtDQsnsd/BFW70WAVUo+exNa6vkTrrivGV
n9hXqXe5S3x8ymzyfE26a4NOwnW8itxmHgMLRUAsezZUSI114K9OcwxXxkF7bX9RcaQRAnEESYvL
yVlXxtLtm8ioDChhO7ssTRkeQH+4P3jX6AF9u+JX/sZl79GdT+/SWF30VHACG0OtUgLssm6kZSyB
lHQw3v825wYnhsVjng8+unQU3kCQ/dE0q+1tOM1Vk6yFKvtGz9s1KebMZbw32jUmpAASxAor2Rok
i2UEf5ZSxKQ71fM7khWfPKZHb+6IRsxgJ3DJzcKODabABFjRD4H6wO7xb+YMhaddp06oVFen8MlL
cjXfGNPq48M0FxO9WRFjBQ/w8WpZ/BwkCc9ipUblkPEWav9czyZohfcAb0KOFjAkyDwxbGssXH4l
ZmKu+2y3ILq30ZNHD8e83e7Aap4E5eOIjgfPBfkQ0N+847yCyomvV5ZhSuR97IA8kbIEksArlldO
yQEXOHIc8J7WdwiCF4vhW3sv6RxBsJUQA+17yjdKccY9lKgsYfhP+rzEBXRBJUiq3WPcY9ibdeWe
BuYtW4PlmPNAj676rBCWnRj2nNKSIIGxWPzUU9ZSLTG23RQFewIuzc3GmxFoXT/Qr/Cx8JRB3eWk
wYaxktKPalrz3jfwKMtvquIyjIAsnovJQwGJP7vH3Azcta/Gc8HXt6H32ErLTkc8st/lrhL7gNuy
gg9YDTYa0sKwFTuiPyj6TMK/jthIOxOVDC9CwRy8BfMy7AbXvyu90BA8UtBIm47BLqSLlYK2mB+k
qxqWnZ/MWnV/Nr0fxksxQQP1y9+RL80/6v8UqrVRLMndh5uRl9+ZYkmR35+i9BrjZ9Zar2RJoDkb
L2+B8e9wLa6VcHzAXbPCwMtP+uLhE9DGYD3jxf2BmSLRugHCwi3/XGDNUO/utWfGI8yWxeFoz79K
85WTSyZBboqFCKVVI2ajIP5R32rn7DyzmdqIVTn/vpQOT/GEa936wgyuoTWVClYRyW/An744OkX1
IMTock/ec3o/1VQiSicmciM3mJ9BEzVHeTnRbHh1Xjq1rDlR9Imce5IuXXCCtTdm6vAkxOnvlSWY
TsKhZOVHiMnLtIiCM8gtSBAI0lmkDJvfZX1mrYilKzBk4p/VNOdRlJE+fiFKiq46cIX/QBx5tWgh
kSF0nYjG9PGGKf/1VpBfMabE1w7wTlH2Mjf3bsWXRtR3T/0E5QVOKo8Z3ji5jPshidxZydLpADw0
Gkfnh2ldlWpPUWXEKH+JmTFm8hmqZsIyvAc0jAmvO9rkmwemJYSpsfIvBFQ5tvp2Gr9QEEAsS1QT
FPqyfctQktFAxJJJcRCrIRbLCntKLXEQXgzdI395wIy6lbhdXumrisxnsGwsD7sLsH+XbONTtDNU
gbzhVMxeuDxwcYAETKTn/st5orfas5FX98w5C8Job08+yf0hp9XiDr62uFrkUyNXk5pIHg0NdRHP
T4lL8plNuXhZ0vo1YJ9ct+XTzZH9D/goAYuUSWB1LC5HOPU72hvx6HrxJdcTfhS5akip+WF7DM90
6q/hqMttax6IRvEzY/nHCQeQbh/bk7HpLERwX0blqDbg3xiROPiZumAAvsNGk1MhUgBUgHwEiKG8
VpEigRKl4hBsD2XWyB7x0Q9w33zwq8gxB6efC7yxJf0nNWbC+DJfi0AYSSQmgjcpt7xaUseTJ37y
KBaoXqvutx7BAIUrqc1QyhpqZawJpjezmNwaj+maUhEMuKFMltTFoet/ztr6kGB+mCyLkwdEHh/p
V4CwhoNkuUuQoZkFIL5bWDXFsDXLoMBx3MiCHN7VB+k1nkR2gwI9jBLhgDTPzQMDNPeL1MQE2MsD
fkGeJ82e01gyRKGQdvweMyHU0y/e/Effc4xXHj2lJF5Yv4hDlDDpNzpEYZOMq4w9l8OXV6ZBv3QZ
p63RF5Lk064FPi8uArWInUGcBT3zg8DnP1zObWoHuUWVemB7/MCCLJTSe2MZmNPlsg69I+icwJsa
irq/sJTC6tI9SfMUFNe1oFHuMWf+nl9606yvxXrCiu+UWbSKNKVy3MQY4YRNcvq0ebcdsMtr7Ydb
rhC/58wNucZP4ODQMVjFYcG8VoMod67LwsnKFXcf0PNrD/3GSB8TwqEsgwGOz7baitn7HHQrKOBS
Xn3wFnpWCydbgRU6AW500E1WnWUgqVeD8PTxbzRp0ov4UFArnFcSFqwLOOxtQzhEbDbkzvyPUglp
dwlhqIuzNJChbixUOODr/duaFAIuD3cz/byz2bRpwfkaQ30B6mDmU/fOiTKB/qKf1N+joWkAdM/c
D61UwzbLaJxmvGo3AiLY5AQ5/6+3GO6PKwUiTun3hLlzOBvKAioh6w4oaX9O1JI75EKDdMlrIhn0
4QaaIi7uuW0WhU+9Yzkld29V40+Efdp630/CPZqcN80fnpBJYubju9knELhPCntBKPVH6qBN9dz4
NA3AS8Hl1wusnlSeNCP4bLA5q5gsdkhnsbqKOSwNl3sGQiZDCOaAEmLZb8NeD2y+xqQr9sHoLpMs
Lc5fQnlyxYi1/Orf/bY52rGML6JsHSNt8cAr4E9n16cAaw+chd/esUTN1QTWVJW30C5BgfC+ntj9
vh+asHr6vc/NH8qfghlTGxTQikZUgtGVjQTw9EXyl09c8Qk3g+jF92LobkOJ25NxSJYe6jg5X6Tw
sSs4RS5dou4UMIa51NcJNIfGwoatIATnCGXQBOvX3QDy4X1jXdL0ZrCeE/0t32V/fOfMRkvJD0p7
wMr89t/XC1mnUpEZ5kwuD4NsyziKW9SytE8OaColQ5dlfaWpKRYrdjeyBjM34wFktcKGFpe59svM
o5DDBDoYi0ORumzjLAaaHtNdRab4M6+xtsGgEwg4Vw21jPUll1Fd5z7ocmx9u+9iaKe97SjuM7rt
URuY3LeuPezf2akNuwPE7gfnKaKGlKVg9quFqvwhDiupqSrT/1+txUADKbazvishs0p1pjmllO3m
zxL6WC6t1lY/iGJZQi4QfHFKiR0JR4djSxwF54UIilEKLzYyZs2kNGkTugn02WECRDpYvS//jbTZ
Xmoj6m1QfQAoW4NyFp0HzPhjAsMhodrW7vAr8vxIRVKDiYoEofHFOPlp5mRyY2HFWTophDuEE3SQ
IFA8lXmBGcsrSFBquIOcr409BDwZsYYJ+eK3ef3jcSE5Az6ctZnNmQs4t2oejjCOFetgNG204A1J
RerPrZZcWZM5rYH+dwjQ/EanhlpbclDMG2MdSWtXyqq+HKmc+3xqxUeTe3YAhmHCk3aUyLqO/mJI
2mFxKO16itLi+m3fSy0ju1CJGJ4NR83cLdsipHgWBmE51aOH9c5YFeND37GIz6GVRkEiE+DImWDQ
XVqdM8ROtpePBFuobTU7xEx9GDIU5okVo1WmYHxuNsOsbWVRytdEqJwUvWhv7tfNhdsizAagwjnd
cGOe2BfPC6UHNevujvDBAZO0WRJ3ipdsq9r5ccKDFTp6t6YP6uHGjW0Z/OMN0h5IwWlxrjmtUJ5j
n9sVYpji/l9QGECMDhLCcRzdi8THDg3XWEletgVzyp2Avo9HGmRS7wZbvHgZk6D8NlO6cI/4g5TP
jdLFtJcKlwsgPTnwDyptXrlqTdtXSP3hEVdUMFhrczGqkzwN9+LSA+mI1BvAgFoVts1m1NdV4FV7
RoFq14A+yjIhzCL12fFYA/lyAljeDgGBEND3HwC3n8IK/CP5NwOg6ThnaV5sUD9BcrfTcXDUCY0b
ShvHcZCneSeYbk1xgJXLtJ4zTDx++HB/JQ4ldbQZ41Wp1EaBEy/rtyZ9d6HH67d5av2yPOYq8TdR
cqFZm41rkMnVsiS2szBGEM3tGlbzo4KCo2Uc97yV/XPdVciQIcNvaXzNZo7NyDpmJOImsbqGZ12N
aKEAwgsNiVieVMY4yblc8hmSIh/lktBoKbBJnSvbjqnEEdA3YgAlYcJ85CrI1FnZrbFYr7zmUwbp
1c34l8/GCyMhXyKEd/o/C5hgx34nEq4DOTZWCnT1lI9cU/PeUmgj77VBg5KkbAuQlGewUiQ1OZNi
H1AIqwosKUfh4KJ7s7mKkcBDU8khXC2Ug/NQjYe5/4IVRs3C8xM4HrfCAbFfWxgwwfZt+1opRkeU
ErEZUV1dClZOTwwdyIxP5dnPin0zsL1eSVpAEFoOydEPYg0dQwPBQinz0vKZxKBrTkC330J30XAE
GKADWRBCzITswHX0BxOzgtsFuofm5r7V621syK3gfpzLjrtQSVzi2o5kHmmUolI3/UMXltJrpkUI
xA7kmlkLFlbPzyDCYCWwv0W3rTvGsFm0GQkiPRbk7majhpC2HxTNJvf0+WNp4QsVxtE2yUcJ5pse
3rG6gNLH3LgSFvrYVt4poHIYBCyN9eWAq2/vsOU7Cnc48TXh2BfvqI6YNg+aWUNQ/hwj0JiHuNOr
Ot/MyQqDAsoJ1i8heS9wHBf6SC4+vrukWomWmmGF34mgcD0wWZ86FiSEJHco7/Hocz2MozYW6hsd
o8Rsav3UZ+ZetgMQajzP+Mjh4y0NNk4lBK3asMaK9OPuqPAA0NfdmQHbsiJLXhUCEeWjMgIZqZBz
X8bNStIVdn2Q1uGz+Jga13WsqoukhCx3KvDSck32WUdFqMEu6YYlgEXZJD+HVMFryhIZf0GpB5vN
olfyhsrbZPBlOGJIqcv589t2oECrbQFwotVMyvXjFqU4CJ8MOGNdSzQ+Aykh9um7/9lRi6RnZBLT
T15aZk0WSiF3B9Nk5gchL3dpGrduu47rNxThgWahpDZ0UdzD7DTagDCURl+2NEQYgAUbOXLyV01x
4Au9N+ED/Fi4nDqyPdjr118Ux2G5l5HvuMR6T6zewetbpcgKL968Sds57nFKzErqOhT6BmVW1nO0
qNVdOTuwiEpeCthw2czS1KdqtL5DqFn8KKl3tMRxOBe5A7yKIVC/J/qoYbHM8oSs66bTolbSy0gg
cSagQ5+ATMwwEW1Og2GwRWGxWMQSxh81L4CqQm6p7IJIx3LzLNs4fPLAjeh87uXwBlnnbAtryRUy
3juF39iuIdKFRoCY10DYhdTLa4qXUk3lyUX/QnHZdFQEZOtQ9OtAblckcvIHSnraXiVJ+8N2j5Ai
Dod8fnhnaF8rRz32jrLN9jxfd/ritk1murkzh+Hxvwl+S3wPt30dpf2tNnxPOR2NnmbJQrOp+Jr4
kOP1IUbd5nTErwxAuM0w+LbT6NLawkIdZLF43C1M4kNV0IJL0xaDhPTGFQj8lynMpos4mwuwbJ9G
MO3TYsAdOHiGUj/GMKH017cjP0lO4NLGd4Xh9h/iWSQpIidZ3YJTkf4Vdjq6CRP1hhoX5+gb4yXK
eX6BOWx9MC7U9eIdOnSNEpCrTHF8vCedxYxepxKn3EJOQq/nRlCTGGTBlBm4SQb2Z8DClh+0gciy
7oAtum1HzzpyAb0nbObibjlc3+7qW7llonclnM2fDqY1r3g1TXHcqxOn9uk12aREMnYEdGozkCU2
LpatkwuAB8bEc8f5+4TqfJz5Hp2S0+fEgGj1uQ4rdI7TUcWifMZjxzP+1xc0zhevTmX8TAH+oT/1
K00BWL25iRdIGJNYAbr4BHwdaypocf8bqTtSiPQJdHLVfJJKv43KZB/tweJMYwYD+fO+ukIrfjHM
t/VcwusnLbOL4AjHpQGFM/m+hiwGSgZnW8pZfp6Ra/6QjUTwrDHRtB8N/sL9v+O/Ofioc4s6DNXA
BkDz8OG2tjSKT7ma0qnP8ZeyYfIbaoJSk7ru6IqEPzM8PaLw1tC0ONTM149Hpu8YvN+Qb9xZHAVy
5AThzdwIaFSISe5BBjdS1blFWy0ati9xCeYPUhdPDPZaCeeoo8yqIsoi/MSft9C60Wjsy8so5R2F
yA8PVuP/GXelfSzQ0rCP3uAX3IdGzuHh1c0Qz3be2lzPJV0HPg/1pPtrlRWlsxtFqKna/ekam8rD
5hkbOJCWe1PBpQ1p1zs1BtnUSXxJKJs7a7IU1m14yGAQcMc5GYDTYVAzU3WRh2Fu0armJytos0Yh
Gz6AZOi6RA4jIzdDW747HqMgMfNZL05T79e5ycxCN20t4Wcymu4Yz7p5Gbq+W7drEE+y9BTPiqvE
PIilWkIH32JmXy+sUcpsln91RKQlJWmtyIPB2zLyiJQerEyBt5opH7nCy77+PP1NB717d+lxBXID
IvHz6qFHsewr0sJ7iFOZKnYdtVh1mjuVo/tH4JZEL3O/Vn04hGzXJOpGcEK6mjcSiJbYGyZfGVsG
qbsi7Tr29ZSZoI/L2WGAep4gTEfY12zKqqQtRmWxAxDVMPEfHEwnCzRsnHgUnFkjQQ3W1mdNw3nq
U0LQG8OWiNrANu1TvTRTi2uKnFJ8nUjiag4Cy/yBHZ9YCZQdg8QQAqzh+k7QZTk5TrHTjV/1415q
6oBHLWTviNkVYRffiwgAWAv1m7U7LDjAwEF7oZmc/qQBDA+X5djkeUSbrCq8HZ0ToThy+qHNfUjt
dcOmVZ9sp/ZOIL+HijXLqtaUOJpc7ZtjwiaHcB3CudVb5flRouDt2dS6doAUv9jefdw8vHZndGqe
oEcqPz+k+0IWqAdZnLPhgepOq/SpEwITB3Z33pivTOK83KO1PlH6wHec3ezaItPwT1o1O5xqnY0J
+vLp1MkwvtX9vS680QJNRAtGuVZOLkgiN+7o5x46ClDUTQnDa2iq7F1EPHSdvcnMCXfI6DFxIW8g
TYVRaGNha0e/GO0DNfCrEAHxxsNz3OlbcDBfLV5v5IIrAIgZYDP01ARbvJ8kIUFpdtzoELU0MHKC
2C9OZ2Qb+rS1pf81373TrbCCddzN1NTIwlzVuFNeZZe++qdiUAHpKykPQM7O6viIEMukabZAhyp4
2OZdpcBHXZaxOQ/h5uAclJAK8X3HrazBL1Fe4Vjo23+TFEunrbbfSQel5xzS+lUqCIgbIwyfEgll
tyv9oeUuSoqkpwlmYBw9scKsPfOoIWfe9I8omt77rex1wIuJe0cGQ0JHj8XDOY489OqusrblWLCW
ceHk+a2ocK5z0qwU1kxgD/RBqAChTiq+GVGmzrlA2GQqS4KGc0cbbaEb0Wocet32nUO5twb3Glr7
AysKNlCyc2RXjtoGF32L772IR7jDwgY9aiTS/bzTsq5pVX876xbK3lq3YDpiYP9m7QaPIDpApOL9
jEwzkDf56BLsXMSQlyaS1C2v02b09AiN4cG4V8T/pbKUYwdz2phLJ0Qyo7E1011FxcVuB8uIE7HW
tC57z3+sY4fCxPo0z3pwOc3tz9aNi1i1+4dG+CMULjZAcLlJTp+tF4bU2usUJxEEPEJUM6MzrA0O
lM6yk0ccZ41s0Kpgj7XBDoGdR/l95XwixibfHVZPgvXHoYAZrmkzbum1BFdd68l5YaCAyNexK0uj
SdEjn908BcguEZmXubgsXP1HC7RdUZ91a1l/jyH4Czbmu5GV07gMPvzZnOHAsun1LoxlTSSjRm8k
2Avu1hUT1hLhDCbU2H2/uUpxxi0Od5Ws/j8iz0ayVS7eI0NUworHfn2bDzbfEx3liZs215wZwrZ8
xgl6YC1T7hvYgj6N1cLS8DhSl8RBW3Z8mCbWDxr3/nI9E08PPmUnS12Y4/NvlptTNZp0Nlo0fTDt
FFplKejzIu4/BTk/EB3YmnGt675dnBnYTRGsDrh7iQJ1mCgwoaAvlYBNWiNchqbGEwh9dj4s5n/f
zbOhs4K8s3DfArpWABYLC1ig3ikoPRkYBgFJghtp040bgn66Op//twT/V89utxZ4SLvRWW7OXNo3
iUJlX7sWaDLpihwMgmylFLbMGw8VA5px2RHyxz6T+p8OrDkpDkMQ4QXdh9tCg77hfMSy5lQhugCn
gUyq2i9N4yOCa+d39QpS8/d6UFuRd4e4OFfCwVxoNN767TsRbxbDlV9XROTgxTqnP9ITLHTYFUAp
dWhgjdBVL9icSG+EgY/CtnjIykwNYNFacGXMBQNTBaCwUIMKG4a5WFZJ9iMw7uJYD82Nke9yyYUF
S038h7Vy3JHxxhBx/q/yDqMZA5FMt+A+j9cR7MttrKp+0C90RViZ/K4y6F8eqbf4cx+vEXACkBQG
7wmWCOwKaz8fzdpHB5AAu22fvOBNcOpl2GZmxLqnidFtcUyviKfJeILXiY69BJGAsK1Byc3Hu9jh
m6Fb/+lbmrZcs6pphsaJIHvQB9hIIHJVDifSD9S3jw44LKM5OCVBmhHIIPqVYWYxJJqqPTLfglYJ
sPLg4QHM3Y4sxtKl5FEteGUu++KFCjz405eOl6gN+Tphq6Y71cAyrU+urikQGT6pURC1udirwH2J
6IUZXSgY7b2ZwjNWaBnHrS3LL8m31UVEI1OLIVSFoeGLp6bwZfNsrJOkVUU9eke88gm3OqtcFUQs
Y+kp+D16VzAYgRHqK4qDamdsH6bpQMGfZ2OAgKqxHkI+i0jGt4IWJwivLOViWPFQKRakLsBgGFFo
MyUnLidUo/i3b7uhJFviqi7cDGIyy5pV2zbkB25vkxaHwkdyfkYzEHoeXW4yoRv/aDNe0+KXdadg
6f3B2DrEoGeSzuwk7BuinvC8C/G5N0nrgaMywHIuHVSP59iy3IYeXOm2o9n9sLEYq2Ag9/+Yc5vx
9NJQbzQE3Cm59dWgbICup9E0vXnFaLY6X9DkAs0Zv2gwt3NcTrGwDQQlZpiIzlxvw1q+X12aO259
hE19p6Oh5IxnGGhCJdOkiZcREpB+WWj7HlQ1EzLHikb0vpGu844r51wFYIea9jbo7MqtsmjboKZk
ZkTUjzME/85ORIVS/sK7SZq243QH46Nnr4UWe4PVVIdCj+j//ZWf+WaI2+jtDHRW2UxNDc6Fu7ZS
VBP5w1RMV+HBKksfzy6QLs6jv4sjoH9D6YuP8b+9Bh/qIZJnBMj9D5VB5dRplnhU56LlkzgrT1FE
jnS7+Mq20aQLR5cXWODnhiebyzr5qqPPEsnqMe1hwMxq47AoS4TV3xn4WG9mFXdeQVrafz3vCP3o
YtCUJgigNAe2GhqTQs3Zq6jJB2YsEIcpHKwNocrxPp8M0Ej48sqrtF9zXDsZ2u3P8F1siv0Stgce
uUSiF6GjHzqaonBCLnJjKnsX6/L2KAE2Zlv4XezNrOOAFUS0Sk5PBrJ8Q0TR/GvSi8rtRTPn2YY3
UnU7PKyVdbnYr3YmwJ/sOHdEkNYmcnBKtB5pc3HEvbaVffcqhMTV4KaZnXhe0r2YPR7tSgPUDeNz
3DxjUYY10RHAgZiV9NQIlrCRk/vy8pDw3TN01TZy9RngXKJwreJ+aO2iuplnWIxTPZlWQoOZJwne
h0j+H2hHEr8qCDq8h6HEYmgQzD/UMD3rKlErztjYm3vvNZu0ONN2BPLAqlzJioQw6enWuEV43KeW
D9IG2ZAOHiopmLnCr2hxND5HfOqyuElEhcXwY281CUBDZImHRYEH78W+IoKYiGKJTdww04kfexz/
nXFuwKIZ4/hDFlFeSlQuA22GkdPZ6dSTyZNyrUgNHmp8DKQiQPasPeNiyUKMye8q10bVej8CR3Rw
WAQ1AKlKsWkzkuoeNloVSRF9EV0pl6BMYyz3cl9Js6grVt/2Db2IzuqYtIl1M13Ljdo0HzBNmhNF
V7sKtMem8qx2JHS29RY+vXTmaziyuXo9SgDEbgCKO1gLgKvA7MdkIcmfptPTZZBH+vL9ItXntf9j
FoGcIW6cd3JEgsdarn3GP9w+CMBSi188V7SC4CdUDkJakhuDYs1J8pLhj4BslSl/u4CdtF/y+20U
JK3KACn1yX7ZEaDhQJu99/+aqMi7rTB4QewVYTwwp3KBNxTQ53VkHH5dUbBw+eCE2rw+uV3tNJAn
ToP+GWa7Sn3282x4cIYK1IE1M3rulXf0GvoslM6tF6tuh+kc5bILDjmq9xt9EfCyu9iL05r78VZD
s3t7P7N1Vnq2cOptPEALVPkgjNBQAZmJQu0AS7HElppzzj/KBQPElD8fs9QIbSHhmn/aB4vbUrD6
ATensUQRnz9G8M26zMaevzQCn9JMYa/slnQlM1e2sq7jg0hKZsT7V9qr5ZNtO+2juBLaSAqW8AX4
Vh+QWJr1BhSv6TRNa/VWvf8xG88NT7U3NiBp6euyXUkHlMFpj9rjjyOCSJECnGvKvnutNdiiXDlw
m9glJISYXlIa4t+w2+kW5W7wPxIXf/SDHMo82Sw+uRAf9DPjJSzCH5OlO3AFnT1P85LieL2oR/VK
gZzm8DiF42f4zFRRSo66JNgYom5jJZFTP5Ys40FuHHvI7cPnzE/7cBo+nc31ib89/1HB/h6436i8
nYcxGFKdDBcM/mkKYk/foOug5GObTkb7gQ0J8MLRPpq35oJYzyiL0fVBqfXlMsMSybmWjYNJ3ftO
MLY7s/gMHj05a420V2hWyS7psPQVg0XDIgin0zGUk88OwVC2c1K3mrKXSP+YDRvStiuEnwkl+y+p
pywyyjEUt2voW7t5954wsNVqjS6f3fKE0rGH6IaFTpdL0apqiqVtFOigJhbA+Qgwrmgvgdo0upg4
PhDg1RhQOGhW44UqKII6tgl4la4O0UzdRiCJyLRFr1znRM2Sm2Tuoati2u7YKpxu/Whanpgm7xtB
xkYo9Yg07khN0z6pIEUnc7sSwYrRoEMhLy+ry/D7di8zxA9PFEFWT8wW7PUJHfNpip75x8RGHUDZ
1npc5H2tgRSWhx0EWfU/F185VQu7usssyzbkwRXFm2YDxPHsPMyo/ICSjQblCq8Q2ALac2PWPa7v
xQZnZwuqx4pTzpoFTqMd4f0ctjUjmpJrrQTlvVmLfhvjhcsaJkus3h6WUA6yHOUcRNhsyVNud/rg
oZjxiUEznleCYQ8aOiIpvA+cIzt5OvkxajDLKbISrLbzIVz6DtB9aWjbj8ejFouspstNBIIs1HOF
6H7ToXKQ9/W6JbWQeCtgXN/BbL/1SpGYH9ziyOO3NXb1eLv/03CtZV1k3e4EEBJOp45duC6QGnt8
r01Pz3MFUpMahIQPm33s4b1fe5DU5rpdohIHNUcE8r7UKDmej7ILHCbSebik+xrT1rWyn/GyfnnV
37jN9+mxWPWlPt/DTVXR2LxHUAxdQnMLYbfEk0RP3W60xLTtWQEorpgDVy0DMeohZzpP2m6q9NKj
CvHelGRFi+medn3W9It6q4ioGjb/UvrUxqBF4JCEu8o8IooiXQJOuj7CTY3wMiGXb5rGORhTOY3j
Bsqvpo1sqIQSxfDX0PrctDkTupHah54zFzzqXCKNo0lLeadRpvwuQTqEV26VKgi0W3oYFZI4AY86
HghAAqEE8qBa7sallu1OWTiNqBg+YmcXUBlQ7yrIFGLzVpvelphajsnx52WR0pPkzP3/9caTW4cN
44T1UOwJRQLuPeI7PojvzsDX5TVVGl0hc+QngBqvbcGz5JEDQg5V8Gmg+MK8999LwUWn5Yo15Cnk
y6e+cAkOsMG9unAJKuNYpvlT5as2wJbVNGWG9aL45Io5hb/90eiaQ9ayEJ1lwoIV60b5mTDiNKtU
5PkmEPvL23iXQLOiS2ZGQvo4Sg0DD8CuL3eosiip1jeyn+sOazkQcysn0WC9f6k/l7ojx1SaxLdE
W1K5mnZK30JxlDF0/pMLk/21L2u3dsgEInqJOCEdWcZdoYtaJRWmvia4Y2Rn5d+l5pVTOBoI32NA
z2Q/ycJlx98iZvzPpHsrVRuDuXTYF1MmRYiSK70tOM3MbxgWbsGIyaCNDjbpPYo/SkGNfVx81nCd
a7T3g6KOVXYjzH6Pb4iPX9r6vULlgN4mvVTZK7jeQlWup9y2C55tsfdwlOjAVoRIk0ng4QgH+k2K
xCJh25dF/5Co780KOXNPpkCoX9/43cnUhDn+1q/1u2JoCqtYyzJB4fOBV1lOHSwJG5EV3wIsYRVz
oKIk2T0LVNV4FxT+oZ2kzLQt+CRiglVhjiurz50qPnGMrpBMJ96LvUEZCQbfDdXB3pVnsXf2mHom
03iLgpLWasIqkXIqP1kj2QswIV7gLdLQoxCOCT59VL2tS30dheZZK/E/yfXeFbgAuqJCnV1rU6NC
zVPuSqUw57xSH0vIsIJt+X7qfXKp/vrdTJqUdYjLmkF7gKS6+QFWSmRDurJ8H+XJdpFPGrv3qW98
oNUzGXtDUyWtXotFLgkfhZOi2xFyKKDUvDXz8k3WPjuZaIj9e4nxDNLIbBpfkzNgy60u49tzDZJu
ngzx7HAtdtKFr3jtYPZb/bZIYbFmbLE6eYRLe72vp8StajJOqKYbDGreITLHb/GciuGBNtLS0xfT
rO1kHG0TtWE+Z2MoVZCxVYNs38rVZoT30BdYhNIbCdhoK6NmmiBTJNeJ/+4NnFbDG1KmjLgECTTP
A0Jv7qHemQtKmyrx7ougVTK2XoORcGS62kA/HivVZi/ta1uAThiDngsYXyQEcNPMRZANqPmAXLDP
Dp7ek0Q9Vha/w3N+JEBtVQMKIFTic3b9ueMTD/kyZktCu0Xb8LHvy0RiA/BAG5QPS58qlEyiXaNi
St8kC24FmLnawbPFR0AT/OByudZFN/BNn2+GLWQhlyPkyGg+03CRRZyA3/wNBO5LZyV5uZOSYv55
pOq4xyhUWHjaUQOwXAu/UAodhUddaxLxqEBhRP3lFAB8G8silrvZ//1FflWSmtAngJDUj95KZbr2
mSHA8TonAz9FVsfIRDsMhGznx1fcLT1WkncSLe4vaacxhdASn4FEWI04lkwsm2IbyUGcQr9ocX6X
qY/DWBzxFCSqWw36lqXCFvTAXcnwF0MQdQlS7udKcA05/NhGdij7wIzPtsOooYGs9HYTlK9RJ1BJ
8Mrf7HBvcuRmTpDofuYVEJF3kyZGcGap/j4Zy1rxQ0lK8kuN1iHLvuZD9QcSD97Zn6Gpm9ko85Yv
OD9S2OXTMqrCOePvfT8gTcUAFfgsfyqOffDVFN1+TZZnWpALFCQhf0Zl6Tq4infgWjSGSnWQzgyy
smWJUkEPg9SR8nM0gXaap0YPcvh83XAWiPtc+YlgonR4amkfg2pprHWAjQ6Kl5vMmx9OHM3PKCvj
ed3T0nhKwR8KqCIIV3tCNapC/xIT3keyRm3eZRmjoz1HHTPuwCmvCfNxwPGvGlW4vsQdgaxxJsUU
q4efULR3nfxNtH0oiu7TchpnPNatyP9dxFE5J8nzj+WxFKNmuCRAr5dCrs85quts748SPK0ExkGl
ntXfxBLEjKsqW81bBDFi61qVixljnuAiQ74EQDRj6rq2lEFYEvJkQOXawQaT0qCVbWM4TauvYTtL
CeyRZsm7esbLefBD7cS3mCMnr6ZZMznfJQILsMvXjIDicuCTEB9MQd5TIV4mOw++CZBItlyPhvra
0IvUX3mQCpDb7G7iYS+wvfnzuLDSqlnCh8VChK3stPxRwex1XfFg9aqI9DscqDblivVYobot9bzR
ea+Gci57EzNosErMlE6BBvHLr3UX816POUTAhzeVh7Bjvc+cWHo4yV5NwHIGFmNXWhqrfhXNEYrS
BXSEm9gJXmfSSLYJIz4TXF4ZwdWwmgZ4/c+XRnsQ3dVJ1axf+3+EBxnEonIYw6sKVgSP/y6FNmZb
s75qLUel/Wthnno6XqONBDGDM3Cjoo09aS6KQU8oAeEy26YaOZiF+0Vsu/YFkTMts5+htMOeHnWV
Sy6Ao4ltdvxZrFEzEtEZZSGDkI2LBjFY+nT1wjzRheQO+9QM75pL6jNQ7xfV4IMc4UF3d7nvqH/C
Uuy0DWDAZtXtJHkOmE4dA1dY7590g9tHIrLJxKzwxqdMMLW3klEwuyDP9rGhjXs1Q+BakrUZWDmc
8PNWQLxhhq5zSLHDL4lj/NfWw/FdnHHwY6HIZFxXP7OGoKdmehHT7nSG94T1ofXzOoEqqS5g0tCd
bVo5UStNycqKH2iI5RoFVhD2bNLesGeQG9prg9+KBMjqc5bo7gW4elx13jVwRZ/8kOWLhroUz5KR
bZwLpvZi+MycCXRc5Wb9Qa7dkhy6HKliMGmKXDle1xi16x8A2uxy7EVWYymyyChs8LvXv3X+AzIn
d9tz0h7dVE5q5mh6l62hfeFJlWpn0Ef7ayFOmI7WP4KChl5xsBi5GBMR04sfggluMsp//hBTr86m
uYROSWIyXMw36mvgTjI9VPJhgioM0blKy7K8yOHkzrcRj5jdUT4fLPbvqk68kom8xZbsFoypYIqT
rvsFcOMeUy7mcRmKOSmVzcqNkFWEd9MMcFw2ct8tHpgxrgBtlNmvcNkywI4+JPDuSF9NVAAEIToT
xP08ErgbJWmTa/A50VOqGsHvHErdYSrxtU/lFPSnLjmczOPaKHzeTjZJEBQHXGEVQBCRiCY5UIcI
+OcVNnnLFYeC01qiD3P2uMUefbBDvFPXkINFO+H2Bv7UsSJRwuSUtCyXZpzSKoF3dfMWHlHolGnn
UfGpeMEJMHgBimlENx7n3e+luMq88JmJzbweY4OdJUNe0jlvDQ7GX/PlsmgM8N9cpCJFSX4WfqCp
GrrLkQ2lEmB+K61XmYzodOhroQVy3gIWA9fD7zrCPle985+Wk4kGFxfF2jJ0zWqNitDE+CG+yyvQ
UUAXOsyXVfgF81GDpdaZHmLnU5HF+66PBOKtD4rLCBl5M4rgpjIhR2cHfhIBQMLD6xgvAS5nkDGk
c79lWBq5kW0BF8wRfK4tp7kqrgOs0m5yiUwotX2A6uzgIyGotjKIS2XlY58H9vwDlx1dVwOF0TnQ
Z04+/RTqOyWS7rTUM/K0VapB+do1tccfTKM44Bd+38kr9KBOv9Z6EduyR5puT+2hOI2aduYd7BsV
2SwheRk140dwwj9/a1pTpiyyxUsTzjYJsspCbuaUgPHVb26KhauWjShW4hjRjKJo352nxGQwrxoL
X/04e6271Y5cUGPGx/ZMzrhszLm1Wt8hde9n/tUnKtHnA0ngI+gOO14hwp9JovkAVtecEF0vaZTU
ILjDrJ6IQT1rerVuZ6kL+PyPYO+A/edUcL0j709eeD4Jxb6cIZ3CZWKQzCg0xXK9tt7+aZqROY7H
w+Z6h69lWqyljYXY5MosIyzlS4VHjr2qJzukj56yCff11PbeU2FNPOZVlLz+xzc6+IwTJpO6jMcS
3yOoyPGaQH49uNEAoDo1lLJf5fi5w+5lOjvXQzKc3h2rfzmX4k4LTTEKuCpQxddwSUoBd3fwMjvx
t4kUEQj4FV7GeSC7qXSEOd0bGdFODaeSJ2NJhWKcZw1ircHdaC9e6eLuVmVSM+/jVXr48SqGQMSK
QQJ8yBg+UcJrVcds0BHZbPpPaOE7pL2MXSFuZ+RzCoXhFcuYMncOFhMInshLoiR4KG2xvfRe9AnI
V0f6qaUO87Hqq4u/ebBVDWNip2s3I/BTZ1RmaF6NichJnvIhnm9xAnwFTsAsfSOR2/CUw10UigqW
wOMIP62b04/wJCv5tyS4TVfYfifeJMxBSyFiIOIkYdjNHhiuLJNA591OAOj1Lm6VQ7JYdx0Ias+d
FwW0zeNfSNMU9gQttEye1lyJxv3bNxc5RLClIOgx5lvI2XMB/L+7cyaKG9dORzdIEkR+IspuCGEb
DeDVNqTFXruOq/5tsElPAr2NMmVwMpAExPwP3ytl3oMd/VFLOU79H+KQ3B1+ekJuMU/GGIh/InsD
0jI33SO0lwZagFlDk5aUnFHUIcgX+9c6lXpjPwhL//jV8EiAaaym23a/Dw6L5U3lF7lCi1O2lKi8
uMAvpEkDCAsuRLQ2zBmww4zqumJpELKAHNCmeC3ZLdedT7IuQxrZecZQihKFcag3hDmbS62ZExQn
cvKonIBdjzjJJCLLGXsqdPmZRWQvqRGIMqPSS3Oe0v4bUzr1lDpTsz+M9GbPvwP8QMN2Qkwqjxhz
L7q+jsMShn7t/AStOTrWT9Rnt6wlUz6kvYLgoM4hnunGDa+740IAytldrLoK17O5TRXVCYNZqQFc
zGTmIL5Yvm7m+OB3xX2UiC8NuEGkha2Exmr8V2rTQEq+hWu1hZYH4BaPVAo4g/P6vmT4w7STfjhC
CgLrwl/Tse3TgudbgDUNB7sdUBB9n9xbb+y9KSdJETOOUvPPCdJm36ivtOACMp/6Mgaba+HWQWru
CynqFQ1Y6Q07hfuygj5lMuDBcqAWZFn8Ey2LKoK/exeKmwEzVD9+XKdULvrdTZTJXoHyhS54YWKN
Zj4Va/Aj7P2PrqBZRXn6zsggwvPOaR+VoLTIMdlMPimYg5cy+45BjNn9JCYm5ukueCUqkI2ipznn
8K1OQx0ftMduX7C7oz2Z1panWLI+78vRfE0ibfXK/Id4MhOcwViZskWTRO4Z40nWHaVSbwYfLfVj
RuWdz2gYe1RVbEAqmNYCkdL14FoOfuyRBIP9r8WMDumvaV5FNQImDBbuDsypjO99Z6pWLyUl43AE
Y1ZZ/zjwhZ+Wx1M35TaiWNAKsmZbhQyzEzzE1lxe5Tyv2PwB/mj60YoYIx3a0rmmuxwFL+KYrqeA
JTH8Oj1PYlrNRuvxQGW94cGi5cQhypcIR5aq+CSoh9vK6p2IhQUrYlfm2rpTbqu5zcMpZVSvVmKl
qSWxKjH2XWtT2dokJJDnaTtmoCBuarQt4zSVsBqEjQj5abBWmJnJmQLRj5XpzMi+DYN4Iizxda03
4zg9CsmoVoP8s3MC/rzZXmb/LkGlZbJXhUAop/7184p0xcLpCeR2tSQbkJrc/9jLFvT6TrwSTDc5
p4Z7Tq/A22rdq1D6b+TxkeSa2kQYmRDBXsbOPtMfkZO5TilfIe4HRzmsfxS2TGGsIhe2Dag2T6EE
fEl0r21nqNCRPCc5cd2aJjFZ9sJP2nRqle7uYlVhNs1LNBr556JIgvIduX18V4btz9YtXfbmaU5w
xr8Z5ZGaPsPkt1/xd5h+QtiXnozQ84IdQ+Nhz45V2DoR8yqrE7f3KtGzPURbQuOOg2a39I3ka6AS
RdPyoQsou6r+qfTaimfQlrcbLlENseEU5HSI0d+KrZ6HlQDioFxIXbQB/b/kPyGIYMxVI/D/DRry
/V8SrIM/WBYEXz8CqCOpX+N3ad0/YrIxVlh45XKj408fzwceSkpU5mv0BKCYnoTjMYxej3wQ1DfL
JfLZeHT0PQqeKcjc8mddf4t8Ot0V4N+/j79EZnsuNCHTyfRrfmlS6TwiNB8zYeNudvemkGXO2JOt
XsrZIpiCzIV1x+cPHMnTNaVZsQAOswQ2PL6BoQa+apAY/3ixkcLnLMPtCOv0khySLVIfp7Cxw8FV
b/f4maItMa9NCfIfEVfllw5fNuphwJrqvGTbUWhnd8A93c3k4Mm+UOoL8GNzlF/UwDcUjR69/sOh
eT3JVzpqHBR93+9ktEa1QZCa8rRfP0e+IdWwsWgq1fV7oJXfSgmZRBJpa7lbSThuNJt5iuyO/r5o
BcsdJaTpw3SbCCCPl4Lse7Zz7o0AtVA6f9RzrzMbg0xQzdc98NeUWdUHklKG2rq+kBpcc/2cM1XI
flrdyhpeT5Cbl9LM7F7YsC/vhf+ovCtRJHnP2M48bQ8OZ5DUfdyHb4erHMXnFaDH4X0L3H5vSKUf
v3F2b+G+ewW+alTDPayIZDblBTJgJoiHxzdwn6M33hRecW2KnxFCf3bMB/GmQ3k7WXmlViRQXWDz
YxHF4btqZgzeEHtfzSuTVkFztr9GIV5TuMltHsqf140pE0g0PbLHOoVVcgayAUA490wYa9hu5IcL
1zPa33ChsHNW57e+X2M0OkCMlLDoQmigICxOo7r7Vm79sHsDVzSn+Tg9WvdKNdA3O3S8yICi3/O5
oUveTg0/esWIx6P3kGoN1HAycteSI6wFb6iFWSDEhUq/cgd38wfwrJA3OBNATnwLDrlRxsV0bNde
FrkYv/MNDCclNkwpcEweU2UbkJLOWzlTWyciTE3+mtZUnuHjY9XSgDPCgGk9rl8Fn5CBLnwrZOcM
KXKBwS9cu1xyDuOQ16O7TiFXj3Wko9hjxoNG2W/biYNyFYGSCG3+nyjxjfraly9biwxzL5kby2vD
9Mz0r7tVAwt8qw//BhKexY5hXJ6+7xNX645JZ/bDWGbFZo0Js+4XugYKF5fp1EL6ZAofoElbz8bP
kL5cMQdERfFtKNabJyondbVJrACofPE+iqX4fLdUXolJ21S/OTo6iCSp2OhBooqUhXVoPkUrNHMX
ksl/c51nUmDEFuMQ0GRrdNHs65vVq8XjJxBKWnPHSCDQ0uii+H1kXVNcg5PmgUKa13pD484C2DuM
D5ve5h32k2UrB31f8+q0+P4BB+8zxy564qRimj7UHIXJRH6xq8M/GS4z1cc0somWOYSbvvvzi335
wfdwdKkjpsfXzeDL5+D135U7VRWmXxQu6cTVUEfCr22VU4K5Hu+OckZXcvHB1iGUVvsoh5MhcmWG
NOgNHcvXqE6dDbIU5qC2Cupe30Y1DADKUv0DTYu7gIADxHi3VgxhxsPoE/CSv2u+v4ZVUBBcTj6f
bx4fPXDjPQ9XnGXGS7smoeD/9NiBNKh7ltx6N4BhPcJ5Vg6hdFM/pAXR0LQ2biAAvscgO2YYQ1pg
xDyNgLuoJeQuUoKZgUvsm1R701JLlIJHuZTuWJdrmhyhVBgnwZtsSCtaLD6wdcUxv2iSxL2wGCDO
5dJ5O8rSTzBd0ZO35yG9aP9Fx8v3P5cMz7ciUfmgd3LnbN9YTIwsVUcJHK4Epw5kTYLxAp2TXyiN
xhxrKJBSPaMt9CmchGSIcTuXsNVAHgClC60k8bgBCfcG0MmPYnVMiRSWgW+Zl0GSTcc73juitEEz
QA41OmbS58NjMsWGuvPRsekc24zOz74fpzlDcLwY3jEa+nJQfUXc35uMNJ5M2aopTQFJ0lcrYHxR
CkA16wtLuoj9UEDIFpuEWVIEwaaYmabB04ALrfmcb1KtanfeRhsUfUKP5zq4s7cC3bsvbC5IE7NA
1j4TRefza8XhO3wWqml+dRehDnUJXzMUdIAldyeld1tIaxp0x0tDnt07HekaHaWkeb3GBxSklLGZ
WDOn+J4nDp0F/ZFZ5hK8jF9jI7ZiNjQKQpnTD6w4ypbWurzW5dxbRlhJpJPi17sZzKKVmB8fi32g
zYYIABVAZooj86kEun2TSoDoGXS57TnL9t9/dWeC5oOin+xf3z2F2bdL/pqFLfeKSIKVfU1FquJu
3JJmDup4u4fckeVC7wTovZqy+JemqN9zZaXod7pCYl1PtSAcD/DwddCthKMKYLb5rqE9984vOqEW
7G7UM7ldNNrR0wOQk9kgVN5tduSqwaYWuLM4SAYugh18EoNfmDf3w7fn8udloodujBJFRqKGqtoE
/t1hjE4ADsmlvcg9mwMciTOy4VpZU15c1byHRicNryqmF5uGsoq2Qh3yt0yAvbwSEvaIBD6tyTB/
yYLgBtBOh87+nbLLZk05mOiMgJNPRx74CQtkBJE8Ur1yjd9PeFnj3EcaZ5S+GAzWUTxjKxnWNaMl
8jh5TyJlqshkAnw8lwyf/F8gtL6adS60LB46QFrGm52wQoSKi9NcXIW4nt5e4maDNsTuR2MgvB/9
Hhti6IC+HlPyBp+N1K4xHNBVAcqotyxciMJ5haxMK4nszpSGflgGCE1I9cwRE/dWGTLGXiBRJMkp
pUsTYoeQEv+gw5Gq2UZDEkxQBfw33/SuyK/fehP0mbbSVHXgoDr6IzdQWcgLSbED5yHIeXyOOKe+
ebkcm9//D7P2AuWJJ5a4PoAvH+toOfKDngh+3jyXAfl13KdUG1kBM5H2cRoDUTCuU0sKPp1310N6
Z2TImgD0eVSILQSOtpn9H9tSDD3s4+E7t64WoLvRoCufEgCtFIZHMotmZbAA34XBV67JS7nGXbU8
ZLFyQSrahtp7uY3+VcFeJbJcqdq4zQ9SLMKFqA8Y3PEFyWaSCRNbaWRkipMyuttlgRBf/Rp70tHp
eZOOdSuqPVYQQXz4TFyJc5uxfGLFzyXha8c+Evj/ph8SjchjhvUREwXgT1kySAL/WpSY2FMlpPoB
b088Yxc4B+C/DTJbl+ttl7VuNkNtr4Vvxtj4QuFXB3Ft2o9W9K5JGHjQd4fIf4z0nYqUv2lK/zWm
stCy0wr+oGSgZlRLGsgc57pQdlAG/mPwe+v95UEezePItTsyifye3XviPwOfwXYj8+jVwVL+pBtq
IC48vD0MjyktugycvGRJBxxALlU1P05QkhfYWIQ12rxRdkCuYoBCZ+G2NTA/P8o63cSIJ5kdvM5i
KBK91wKcK51Fg0SkU+829BHXjUNHjlrHBFug4jKozBbCZX+YVAZ2swL7cEK2JnKuuI9gvd6CBaJi
PhDlXzmVO86poQmJJUZqGCC5cAvWrAuD2XPkgHCbS77jZggXghKYHb5lbpKfxP1wcsOESGkyqZ/5
AZ6934YovaPJdUK0PJ49iGiPrRgwgo60C0sE7ciLQlRQttRJVl7JypAqXOCu9qUL9/UbqfCuZBUI
bgvjCZ3N7o5qRW2IMX18zEUo4ziDUdgzga3FgVMG1B70XaudcBbF1ob7Mv85bcnmAUISBiCd6Iea
XNaCkK2vYj0cpavYsE2/FYrW9NJZ/OskCSF6IQSsHN9qlx5aT30PO7+u2fg+2nv1ml0fhp3tG7HK
Pk757cgtuYhYJzjZPWfvhWz5klIuF+0NjxToK6rTy1uNY1WQznUui3qDBvcDdRchewc99myafRTu
O3DHxTqGTGAkJwEa7S721Z7D61AS6NWJHwAuZr1Gebqz/wokta8Ilpbn4ePRDG+tMKiyglbTfyBk
+LOKQkU2V6hg7/5TH7S4iG89oCJENZ8PNPdCple4eQ6kspGnefYzfP74sqHc6JDh0IEL9aKPvlR1
woJsv7352y2dfCCXyKpt9IGgr4qXGgh7Ye7QGwwl3vqmI99NT2MOg+w08uEymwWT4hth0z6RKac0
LIr0981bj4yKV0EEdwSN7pT7VFr6LGLWTVFcA5HlO0yWjPzOR1T1CyrpHHkffWpRnKGWt4U5uC8N
ClZvlZUd271HFhTW97L/xuuCiS1kLZQEfCdqhJO5FlMr5E+q98EopVlLy1wYzyYYbjH5Sf8zRVbA
ImeHh8vwXgzNLz2qhMgwW3dR8Qrf6rO0wt2dk6Je9qJCpZMfNJCSt9PopfkAhSLjtFM6TEXK03Ld
vBaXkFCF5vI4vHxPYIIuuJXX1SdOBkTXOA7UTeWHV4+LJrsD2pg+LYUZw3kyTzFgqz2sJ6h9yATs
UqGlV6dchn8BxLnkAkHM3ROvYVULvo72HXOSm/PwvTjvjBdfJr4yDH6o1bRcddNq44b/jvvf7Iuv
vSyI9J6H9fg3xXaKXNNLI9iHnAQiS62w+13ALulYmlXqjU5MucDO6Igz9XinAx7TrYJxUH52efhs
jojy1PhqAmvcEO8xHIuGv7fCH3DqFjwGBEWGV4Xiqhs2yfLO0pM/f8UbMusLtQ5QMvj5NGyqncPd
zNS4CZEgCj1t041eqYeGy8moyHK3/5Gr2d6UDHxWfguJA/SJVpJl1i3xDPewKZkI6alT+xnOu2wd
X7eK2XlOKgxRnk4IwhdkeP800c69/NftD0Zqrt8fcODqC4S5c+N9oL22ABU8V/Va94pIyj0/eGcm
5ZDClSl672KjfCzOjVQDl0ugUprddI6lQkpat34N9I0s6JQ8FCcdlRbCFdfCz845NWGNW1Nq7nhv
1EtwR8a1DH+gxB5Y/5f7ngh0HnIqdgfMq3BzX0/dBn+EKgKLyjHYDQmqRXwhFo53ZGu9DS2iNLGO
XmU7g+lsHw+BE5fUFJrvVFTDGV667C2okYQ2SGwmBFNxi1F7anZ/BBv+ZRod9Go0xp4hgeGyqbkR
h8Yz0VZKGHM9plOqzMUNHE1ikprESiH0PHlhyunn23qMQrXKnRajPojdzh73d9ycVq4h2A54JtJz
YU6rnzKU/ATwTUnkLVYqUPOnZ/wunD5/nI9nEYB1gg/cTkIHcpuOEVzqLAAKazn8szro/1F2Pvrr
j1uuO/4xgfIqGGClpA3wzRkADZ73F12ntFHCDDpvAV5T36njZxMqcChzt+ygoJIybY30fin023RA
2XiBNfPrp6oFQyyrEIYzf/zh/17p/y+X3L4ek1W1aRERHxSWwALkGH7VDhLBw8wxa3Ii4E7P9xNj
8PISL8Ieff2VsuB2xjmnlbnGae2cXfPrEM9eXnpsML62v0dhryvwum33CqQCxWkbtORz0+43r8WG
BInVV/9BfVn692TPvylq+F1vIGgLv777ZsPeNhLrg9I2ePMBZ7NsW8r14zG5SviwpgrkRoa5wx6D
vBtJlKha1AcISURMXwzcerXR3R+JsMfOSgwETpFnWjGcNHtyqigXCV3CqIMbfOYagYhG8XVwmm3a
+R5Nqf2Q47v71xbMFce6Q3dNolWYBU3G/xx9FFrBAMBf0bvRm7C9l2P7K4I+WYRMtI2ZDsENfL9P
66UrsPTSqqcefZVjK/cYUfi7fTZR/TLfaCGPEM/weMVoL/+HTo8qBGeun8G3Ahrb2y8UhGc48Wag
vCLoEAR/kBZXq9/9zkI5oseMkVqYn6OYaH/IN/P/T66vxhmywDwFWlovDuVMFJttBKjgP3uoPkq6
P226bzcd+PTlzGx2HppRJvbf2AY8j6cL7dw6OdajT8SPFbPIBy5cB7QOudLd1da3XtC8AhmYWygb
54IDdKTHAvww5/yc/cTqkuAFaCPuGtN3ipPun6fzBYAgerxtV2yNf0GsYN72TrNzrs1fMY9dvx6v
uxKBxErth9nP5Lhva6arpSZUOAaaniPKOqbxtMBpvTYtgJ6Lviat3YZEVYxwFm4LGJEW9KpxA/Yp
YqkWR86xgQGEvgv0Mc+yU2B0WP1z1gdxwzPFqsYS8avHmn93K1M6zlOpaOmhzCrZVOO+VI11g8v1
BhQIStI6Ujz6esCO9IdAMzi2U1SD3h7A0kfy+A7NN1lUyjBF6wuGDQnfzRXiilFBmmBbZOIWdxWq
68XIs3htfXuTWqj7vkA4VX53LoYCNoki0K6wIgL8XimOvKTe8AXbDW5NaJVPICcmrRq2OjWUOw3A
7Z49uR1s4OMeoLCnCPgsDjyqX7rFYczFysjbLs/i+i9DsH19j9ByrdVX4O/byNGUULdZ5vqpJo3m
bFraz39JKgVbSsJudYQi4FXjckv4xvMZoXEfre/kas9nf75R40BEPyrNG0ubAMGQZWqtd5ygszx5
cl2xlUtg0Ag8pfS5wAklc67Fmd3ETlokhDoosF3WicfYPJQyGzWvPt4shQnIStMlNH5O6WmSVXo3
5JF8Ds9eLMr+jcdsR9Q7it1UrX8tsjMxEKO3oUfIUUaNJDGav+aJkZ1zA0q5qMQWV3kmVhzZwvRH
4ObJmE1RWQTfGqlg7CFbObVyjNqyxDXWYan4Pk3dIyhXd0IEq3dhCdJe1jGFaudbXmM8onRblgXh
A+EPme/PYIP+ZYiHxDRJcn84TlEgazrRFBtVR4Ue0hDUhcmPNQI2AGu5iN/XL+zDU1qooCU+VuLN
sfsOxoz+reI4Tt6D0scPvdtqjM6Qqq6OkOPemfkS/XHf+WzyDuEv7uFl9QCL6ILedKTDyPrGoyns
y9Fogl+PDx1F3k1HX4jn7TW2rmhB/AHOGiWkpKacajt4KfH3Mn6n0MD7CZS+TWObSCzsb0dwi7As
rLkTj4ALbor58R57vSQRxMxoc52vKJr/AkFtWxLQUaJM121y8qxh0xYN/muKrVnYIyTcnKpe1XS2
BfkY+EykJYWXzUJaop3KerzX5rReR2ykfBAgRZEyyq5WppQaQmKfcd7khNZf80mBP6B0zfaoLwHm
NNABQ3Ythudntj5/CK0pwsze+JMm0tnx6z2LI0XfBKf4L3P2tbUbxQ4kjQ6hoQtrhzhG4cRn4967
ShAceO8ZRlpEZXOTZ9Eq25NSbrIfPK/lB8cVJEEKagG1pBANoA7jPqctndaMIpoKoZ9UKc+YqDI+
Coi8FfpoFe68PMMACekgY1wrVnB40u1Wnkf+46BN8J9zB2ZhUcotgwJ+CV0As7Meaf8Zl5zDVPpp
RFcWzSzOg0HzO/7V6y5b9QRyFm3RrrTnu/c9Acq4Kkl3VA+asMC8jawPMznHUY17eBHBgLp8T67o
+rg04I5EIEcbtA9Y+GVKeSPUIxcKlTNNSGfpI5QzLEQZ1Mnv7f7q6eVJvUSPQmU4mwB6QQah0971
+m1+rOfN59KYU8QciNW8PxLD77HB9+RWPoe1bdpgjrt5uPx9wBeySy+7vtwUiuB+v3nh1C0hgvjY
q+T4fF6YZ8JlsU7Zg7A73rSj0H8+VF9BQDCiif7wt7eC5U/ra5pM423TJYpThGvvAoWgrKe3I5K9
Wexh7acWgSUGITEf9JrTuBTGUx8+9s0jq1h1vKGV1RNJ5aFP1d8nVIJo2hOdX/fdY6owCC62NnZh
N6b54WojZamtdt+d7fmuFTSOhC5wjvJa0gvv6iQpIZbJ9TaweAn/VsZGiOb1kZIOIA3082uvOqxq
s4FfOh/n5ncEZv+qJorgnzElbbgh1zsq3NlXWX8AVqFU/Xk3CH2DbiK4Pbs902/DEIVyvbtMccKr
pHM1eBjroH8I2a5xcQW44nmMeg+iFqz/tCmxVYge7Ba1a5zrZU+vwPw4y63vnXr+LTsfBhEwR7rG
iWmr1Do23u4FYC9eGDPEZ5YED0xhMALLWOEE2AaxzqWMWR7Gym9KhbmKTIJQoW9OgSL+cVQqeSIm
/5TDwI8piiqxZx8scVT78MSoXK/beU5pdqePdJdEV5PwXKM7SmwlcacA2wY5tvE/tmBryNu+xMY8
f4RNjZq9onVjvpOebYRdJftYFTCkbSkzW8wwdd34xZXbN+Q66KxW+O1JxG6NWinBCvEQsiHCYlwx
c3AzSy827cUVHYi3btRzDBhN2blb1RsJQHRN3Lm8c8DoC7mM1Mma+I6YNcFwBXPDmr3rGSmrt3SY
Md/OTw11H+RjT94AFgaSg5LvDwTexunmhPEMwcvTbbUxXHBt/dCwXyR2X+L2hgQF/nZnFcv2/b6B
3MDxOezTJNv0PrIb3lhbMXAMYAGvzWOBRisJr80swwwrhLvgef8G806OIIyvuqtwSeYkuWx5KL9V
Ib9fCtvEiMfc/h22z6fEEzW4eM0XMOor5WBJGkzWEzNkPqcRpFf0O45IPWlj/1iQtRMpMsqYx/iL
VLyWKjTgyAxpFQSAkJtPRD2cGAb4huC8TwM2pzWGvOg/AhqzeIVBn4ECTa7zdqYb0hzcEtS89u9c
xkPF9mgju992L6J5KNxlzPj1MmpFwZTZfuDiPO2dvDyuDoX3M2X31d4fXnLpi6E8/J4dogWiUaB8
cR//v7zT2jD1cHL/ep0enPvps++YLIIrDyHqg5DsVQlHwYeMhKd/h8aOLqeKD5dc9gR9IyFt+biu
GbKNkLxsoNOUx6zsODc32CxG3oiOzn1s4/lKaIO/JBav8C7hrdRVwIeM/dwiHranW9mHOji0muOb
SePzpkPsyQMXH4YknDay9gKWxYDG8VDGU9exApNRXkrhTOVjiuKrv+XVGHnzoxvpoo1LHEWYyV3q
/M97LHZ4irWkqsenvQDf9BaGstvfqrwq1LZNL9N1OWdaktIv3MA9wg5IfpwojtKHHIfFh0tyopvq
g5jWoeqaN1R0+pTemHeoB8sDvLJdp0OjCc/2dLjRdQuf6ggmo896QfPfbRvaqm+8d+LBV+v3oYKd
jzgQSKL//NqfX6tzws1NdGxpjugAmAt6stAWEpUzqVWYjLtoh9d+qF+rp8xlgT1bFtNxYXTIrjeH
ab0aynAKj2I1ef9CpT+FfadFZjtbMASOXs0oi+XhF5yY2a5kD0uKFY+jJngS6/wGufh2abJBqkZm
ONkuYx+ZLRSf2qM4cjC/R9eEmAD9GkEfJEcjuT3TL3M3IPR1PcgWPh3E0Kx59UGFcgCmqzEq5dFF
dB5tEFzuzEm/WSOdtY/cPGZQyoyC9yHofEqD/PTGEc0kOuSzIMVIYgoZiLp28zDoh785KYY51dQN
TaJb3bzglHvN4IQXw1a95360VnaM7Un4x0rsMK40+EAakrQvr+CrYArNcrNw6+apj2gKRXXUsE0g
4brwNjewjHY0zLujO957nmXWc6OT2plNpiM0wJUeRtC+nhVwGFb3yOCnEAuY8pTET/AkILqZ70te
i2pycGjD5X37UReP2Xlqm4+n05DdpLVPjifojTZu7WPTjLLII2GMjJb8aLS0MMsdfejbkBFfhHTW
QgAe/X9qOg6fCTrHACFeJyulCi4dWM8f8FLtRhqmIjLXCIqrb2t6XNsnCGkAIW4StIKjri0Z4bnU
0U7BtvifT1gmyeYt/PeXj8kWRs8Mg/j5hD6m7cJLZFjlFO5ZwFwImjeFMAuJPKdpZ36kiJbMNn5Q
rmHZ8KEwjvH/Jx3Avl4qrprUiS4Qv9W2UPNDKDoteAgwqtcKoPXBejA7tcu5bDGDk5T/xaPBPL0N
01Lq50QDUKLzxBQIuPyTm8ERVRCpFVNLvYyAxTDVA/pY+secG0+BHtLE1fbsH97EE4qaaZiOXvGV
vGo0IcqQnmyqn+If6Nhbabwl2jeKEF7jJ0Im+iR6WeboaVXPDwhySMUDyVvZPrYBzzQMDYjcixHw
Zrh8Be1hrjn3kUhWB2Mtyy2GPMbVycA5azH2bsEbN6pysf9k+C4yBisenm0M8DpRJzPpCM0NlJas
MB64RnFxFAsMt7ejNEo5DaHu1sJYLzMXvK6KPaPAPc9mjQYMMwy/kkt8+M4/Vv8GBECrWIDlQ0YZ
Tg+Soisn4XQBU0GZKAkQNsiCyeVvtxa7VWOfWCtj7PyOgLiOu7tzduZxoxQTfi4ssxRm+fT1hPlm
LVSMo01R8Mvapd7AthpSGZU7EUfnKGIE6fEtO66toF/EhE4B5YKRAt1Mbf0S04VNsg6rw0W50CSv
NPMFvabBvXTC2fqSilPX3aRny6DLkItmOTy0RUBYd9NF9OKebKmgvOqxCIQrlxsyua+mDxBVRU7r
tQWmlwqXk6I6I45sMwIIKsXH/jT5oz+H8YayeQ7fc7R4dEtqTw27ek7IcoW1wZ9Smm/g1E/Lj1j9
iQhAnj56tKkbZ6iuid2jAyKU+lHxKRrZnlRxlFTX6lcP3g2kQTNxZNYwdGTkBk3vfmNXoLCfBLJ2
fCYBKZVaS1vpKbPHglbGjI9b40jt7/k12V8RisNSQJXhiyjRShdh76qidoO5ORxWsFKwiGPntIkG
EXD7zHnr+CC2CFqQq8Jd3nXhxa5rGPAwrNvzAOPC0BP3osa5z8tU0AGw4XOgw3zT7URVZwx29fO5
9gV1VjNwbYVniz5+/7PVshQ6Ps7+yGVM4KygteesfwdqLklHYId8rj8tccJXD1/jM29ZLtbu0Jc7
NO1fA8bFLn8XVli6dZFM9z6oGnKWuopZNGBC8PmHub9dk9ThVKQ7dKhj74VdpYjbVPi8nmbIBPcY
iTnceD8G2jNMlVDNEwp8FjCBsBHhgX3U3ZfAm8pYnY3zZTkLNzcf/eiBT7k6D1Q7dS0OUBf97bj3
86IsubHTK4iXATHve4LnVpDf7kuMFX+E7DqnOcfxhPZ9OJuryYQURLkO414pfXYmW/gQjRuzoQa4
g8eeWAnMHTZnOM47nklx7jssFU/yyf5ATDnhiy/xL9LfYY7NHuOl260wmnMafVAxoZAygu7Vr+Ro
6omYImrrZHLInMAYyybWIpvUJkNfOm949BuyD4KLLhbx69OXcMibdCvlWOpEcuqGBXh4b3IaKIHt
kBVrhIvqj3GApFIcxa0LThdvFGXccT+CJGupwbdKtBAsLdK4Tm6HZGBVHslIpVgSp2yJCN5Fvwob
jyQti9vdac9IMILyjTWtkLtkF6pOc0/BhshbwtMTFWG3B7UyDekPofMaP74GSjFcMCmqmkkJzpBu
ilOYNqdFB4OGwbmYBJRr9jbU9QAaRg2mRyMaM3ydKSTfELvMKc8ePSw835cBNOleR1gjmOuSODpp
cA4QkrReBbo3/eGw7t66gvgqO96Y4KevvoYrxhvd+dleCgl4MNMBynpGGtup7rWTDhLAGeWxoQIS
unvOBtOIFsaliY/efX48OewdePhZ30uyUAzLhlwOErNcKcrzWSX/E/jhSmB8YWn9u6azhtArIUL5
D4dCNicc2/5Q8MLECHcT6yTL3cI+mziMTJ+/GBzE5oJXqnOONYhRI01k+przDmUJI6BX5Jwj3xoB
y8YP+myPT68rUzcUzqSpBwww4AJ8Z/QG2o7sqi9GLj5P3+uESGZdLYVkmwDtgdTGUSTfr1yZ1rLU
Qma62H03yCCDNLlmCq2KEEgSoeKngMHgE9Lp5bj9erNAXd10EaQthOWMEnQksQdF2zXMiPmcg+qI
6kROABUmccTvK6CLgDDoDFBXqRnzda+bZXRjDNGr6ufbRHy0pf2N8IFGhwabLpBMyvnPqF5WOAHJ
3KuPtDtEDwtYK2LPl5gvmZH/He8TIf34bKVNTsgB+/N00pC2qQ/r3VTa+EPgpanWKgL9Ho82GguU
1mT2lDTDnuWnmxtoBTy3KirCpl6shPE4nDcUHvtJ7yDYOAiGGsifmUptqLXeV4ui4Nj20S6dGWeR
A9Q55dvEjhdrtrD4bx4Mvk+KIwRZVOlXpEzZMVCI5j9s8HlR1D/YAnruTzhoh7RpO1y+VO+zzdwT
SYxb7US2Z7cnYluJATX7WuoB/Y1h1xYg9nleGukBYNhSnbdqlVbg+yz0HHF4VAxUnELYFBF6lQsn
tgFT7PYMfOnUHzhzJJwiKHHrmObdfpLOUmkwwDQbb9ydNYVW13waeQO4M2ObCtFgJNuNZDGJL/OM
2akq3qgGilb46yHE/2zdC6GogHTaFZhqg8u5jk43rYzZ2pPrppl3QtIH+7+lmIgZFPD48L6ji6W+
yAa07HmJ0caUsf2r/1ThYynqXFl7FYk8HvZSB+PGNm+arZ42V01SrvW8UtY7QGvTxYHFp+X/OvSg
87RJxCoce1elEpOiCjv6sGjZCbiub17gR7lTlJL8u8uvsiYBN7OrWcekaW2J7oMCYUx6RPsUZ5sR
cjwWdb1eCXOEJ7JbeWQQJHRBxB0eCKDtcn45QTMsHLMZXbiu5zBV+yJ7GxWqsJ9+icNlPaQmK2Tg
xNl6n4eYpOrwfo6LXmFGl/T196vvcJVDb7gmwoEFiwRedScGbH5An1dsS2XHgecSHB8BC6/XEZvy
4zz0lgpBuH15HFEexp5mY8fMFRXw+fJLxBUoW7PpcZTPdysQhs5D/Khh/EANTW3U2fMKzJwoFwVQ
L6i3MNNTxp7wbRrQ2C7rcCSjkoSbt9t/Mih7ka5GBtH4Wai9oyIm917j/eKnoU0bbxqHPYRhnlT9
ZMMzxLwicNoO67PC9zsmuwYVXAMZHcu8/zkkZcpuj1uGpX2oTaQYd3d6qSeqUYtltKBbKxPlHyrl
ZcoJJ8pjEa+3/8RqtnJIJ8BhpD+uv52w6sW84ZHbuTUlY7RGUYxldk3xBnaWKxrc7RgCEeYC+qGP
QY7kjwsCDgKVYrLsiYgOmb1o9wdkiufxRHVoVThKImzmfrYadJJpLBr8p7crH4XBmV1Utkfxki17
PN1cVNM0yzjQDiZ1a/cF03aDbO1XF8r2BG5eKQRZI5WAkcthG84bO/ulId5c3VLPmQsFc+7+kNWv
mGiskRG6ew/vAiChsjbbRUp1Fvw/1Ro3AmJQQHDPnTqpw1gJs0he796Gqj3QPd5cGd24e+X2uIYy
rRzKWvAjC6N0RCTxCpz2nnXNbQzeFlTch9CDu1/NGg4QrozgeqLKW5WWSd8xcC10Zc5xlWvjXSZq
MkLciRNAAWi+MCAoPZASYDEFMqpvlBn08kvaSG+ya6J9nCaBbZnoWY2FzpaLeLjlD+o0L1VIEPoc
Wybu26e8FVUlqaurGbAIe5Kzjtt6tGpYS29ONfmsyZSa8+Y0Ah8AiQ86yewdukNEx7E8v0CCbY2G
mmT9P/EWnetEYkA/yKzgxyVlpGM0pAd4/Wwzqu7SvGcUoNlm4YhQQVRIVidKFqy1QLqbQp8TBHFC
Ilo1nkae6s53QrmyFyOmSgb3qDWuDNREi9+bplbagRdIM6JN03yAeVAjkxHOqzu3QyuStHEFunXj
oDOxEgGQ1RiU1oTsZHSRayLn87cPDR+1iTbg/cXKEPCo+tx5+GQVCEBO+8AviOj9klWaUsPn6DUQ
Dky0elmI5LjKyq5NAdgWlzBZAu/DLHXjfYkgDL3uGmarV+5sUuU91u96udkzgarYXE47hU72GK7h
pSk1goKCQ0G8r6vU612jzmQ/oLfYbyu5Dkh2xXV6CHJxLOrMyzqclUcxgJGaSWsz5cLAhAWyFcIU
9/oDdCS6gntNIB6ymttDxhN9r66DceXGWSAUcgS16t59wO9T4BJ5gw95HnctJcS0L9XHC9Vi2GSl
qdDAPEdS8bj7qb1+Iyv21FI2thRgUIbW/PAS9a3ohsP3rb7q57/J89OANH3VxaEv7MI9Dvwh/JSb
9uvDsANtNjmX4Cp8rm9+kdxBmqk+AeoLCtKQM5IpUnd4nv5mycrpQ2qwJ3BnqhcwORGp60E3Z1gZ
pYTLthV8Lxn21wjolGni3V5KaV9TvaAshgP37t+D5KB946TooPvY+sw4iOllzm1legFhHxXAHBW7
2mx8Xm2pDLarKHp0LJ7ssIluKdiVeN+/z4GsfBK3RrYgQ6HI5K/ZDRXb0deSzspkpJi1D9RVK/ci
+OKW3axvyMKyA4ODOdWe29OhjuzXMrE6BbQwM8k/4Befd/M9U/oHQZPwRHGfvnAZc3q/pXb4Jsev
cs9EnZZwelCmkKQfz5NcWq4H8eytaPKFcoQUM4+0j18ds0ExjWHSkC9QpN2pgqkdLNZdzlL3/Ag6
nHcMHncdKhBZdiPOIT4KcvRqf6x4Tx8Q/h6DnnnsQWCu8pI4/k0yfbMFfTC9+fijcvdc5XhMDd5f
XenEcSHnlZC2GBo5oEmYaf/axPVToT97lr37J5cGGeuGN1prjzjwTPFb4Cm0DZMOp9HbcarXrftV
LDnT3zkV208IdrRMftW6wqgPMRgaEw0ae/TU44lpL29v8XQAb31Borrwi+baaIFyKOjYxjYuyvrX
wnjwGCjQDj52XZAVkN5hXOMB11vcex4+7ouOXJp2QzXo01cg4CM0ZbBF/qaZq7W2ixaACO9yXTiC
A6/MYW55NwLo6Id59R7Sc/iLOLqsSzZj+zBJYClXaftzUuZVTeKpAITPmLwacyuvK0CU2P1MkXW3
P0ldkpELM2xvRuFl/CWx6Img0+XZ7wUKSLWDKKVAKwsiGLPK1R4GDuQaPK35MEUpXYK/CUjV3oYM
zz5h4LZkdMW9f525zglIKoAtGTB2IBAOrN6tHIPMNszk9F1tlImN3qhQPkE2rLKyfvyFCfMhOW2m
Wl09baAvIDv7ME8ZjizSqn4rpIxveXGESzo832Wf1SzY+JpMFony+iq4dWZwUBVJnBwYairdN4Qr
Z7RzyfFi9D47ifRg5mQQZYB3pLKtcYbO9i+hwWqOVpqdFJtVxempIIrYHOPTRJNlJIWZTiHFcqvI
N9ILQzP/rg0Jg5sSrVrpcXQCe6Z2QljEA/zMizezfzORafDROBgl7xuMEHKP+cYMLc+dwKHuBfJw
wmnhGnXtxLQyLeOdMHGH7Q+QsCZ/u/lki03Xc39cCYRcQ+hZZ2ae8nXLLxJ2qOqxjVtqUl3P7jDn
sLMHs9CjwCytm+NgOYaQCxkscMCEH6fRyKl2fLrzj3Kbf9JAG2kRVoOgZdsPxFonQCiFF7sMDLNY
HNEuJqi5URo4LuoVe4fWMp0V5d9WDo4Cf/99y4qjiumcjw68wg0X42i2pOVzRmuZwB4oleFTPJ6U
LgKZm6NlbtU5tUPHk0dWqHHX26nk0x8gIL4B8XJNbUdWQgmn+OOZRTlfZhJ9gJjpxKFuRa0EsLxH
IX8u5cDzOKHOwW6pXSz2yEx7DUjPOxC9ZKqnDgvvxbmqU1Vyy9nKuiv8d+CJknBHWzimOVBnAjIW
5VZV2izjyZkiibyRuWdmVeOYrm2dRO9XuHcXDtkHyUo1OZweN4fXhswNZzXzVIUqUnXbI34IiMHU
letez6jQzM/74V5QAdYCzIchOD9pLOYc9bwcHtPWT/P+OZFfBqSTyKd7bzwWVxJsn5zFgcK0wxwH
Wt4vBgfNk0e8fhbQODwoDEVkCiFeR3Wb4mwyhSLk2Iq7kDoMIB6iBXOC4KTYxSDDlZ85HsMtWRWz
koOyfB40mROYha6JHxvfgn88Ed6HbY1UUvDe8eH9YmreuzWzjm4Sp2kIiP4Kt4sbo8s+i799AH1x
Rn6OFMPGldam5b3qtA1WV6VxLcLQSNTI4nljGgoy5LnSrMiRgRCefGHBlYob7T5wJ4wFrUq308HR
d7bUdz7k1omVj4LA5i8LgS+r67dSU2FHqEEflA1VzQVmQjuvphEt1HWDF1uXWYHUh3KUC5YT9FlT
fUc0AsVG2UQlE3CyOd1rl4u+G6NdcJE8NMUAB4jlkLJ95tTl8jon5JS1vd9XtisarcAJxCdiDaSJ
t+I0WxK6JU9YrOkgPAQ1mWNPw2lSZXmgC0MeTXyqq/fWNxX48L1v28uPlkVNK0rT+WzR76dHOsZv
/AGmb+D9Dt5aSwrmN9oQaqSYMMbBcB2ugemrHuhtv2vgu9fzrZcKJLfGETRmQKCjSPHnKfW5qEna
X3NO7RpgdkUL5EYQYkFQ4Wxemh2Yika1nne1nfvARR8nwEvtqNDrfuRVKIWh9QEHHMTlR3CAkpvX
fgEgiCmjMTkmSzn3kd9oEyZRPQ2sUd4ldt7bZW64Ko0zLMeB6ADNAHhvdbhcFqbtDDxoKbu8Ezfk
fpPXwgLwBjPwJ+Ws1PP6SCV/qx5K8EEEms274xIWB5BxTBIHqQhaqmQlxxvKsPYDGDgxsiv3DF26
e+vDVscfVwrx/2RiqPFHYn/uaMTmaOj2w4cvRNcQD44l1IczHDnyWBZ0ZhDOMFD7s65sZctU3tT+
yH8zT9+MAURf0/3G7pbfFq6XL/AgTo2IOX742LHl9y88WAV7PeWQFExd1V6m9Asr/GB7ET2tV7Rz
/74dycx+eJCXTD8MlndcTfL4/g9jcpG65rX7833wHKXl8a2n5b1YS+ukUSc2IuiWXcS//ONilPZR
OBA1JJrtIjAxPbYpKDVl4Cr6vjYoVfbZODDi4mlQc1b4eXkK7Qbl7jBwygfdV7u9ffRncrF8kRd5
Xfs4tcG8j4MChmoE+Kpl2Wud5dPzeaSaHiKKksDe41RrPc8orZKJDI8LP4CKZvPY8kiWs4Wlgyj1
bD87H345Gq4xUX5KuUDICqXF80vpZGsvvv8kj7NzyhBFYrqjEmzflRfZjR0MWth2Ek38u8XfZYbA
+RkGR2bzTdazyBpeiRi193PUzlWVAQIAX515hTuE/65U1F12zGy1AwVpyD3d/EUoSw2Nzn7ZjWxt
qo01PW/XNh+gJCGvYNNzXPv5deLRz1NXBeDJfg1nWoWXIDqX6XsXpWsek/HTldT9g8O4L7E00p+U
VAtrPTmHekB7NlTtOX9kkm3bW4c55MEe4L/y80FeBr3KeVxPmyohTICFhUwB3c8y7mHkP1l+H2ZA
NSmTX2NhL69h9wovDUtpN3EJcMIvbHRZNxYylb2rnelsOOUekrwG2TehRUkLd1UEe/F+JeXlzCwE
H9KEwg97dXZZP0Rbx8F4tVATydJizIodXBSbWuKUZvENffURMg1NwIurnvB0qd+DIWw34A5tVcKN
7mBS2ij1O7h54/c85TQbwwDmB6x3d3EYIy9Uay+vAE+UsXAmCO2wahDn5kAA4rFO6rGWpkpvUMuq
w1Yo8Qyj4t8VJ/edrsHyZ6Am/L/cDR2bALJhvRmQQgEXqaFCR07ayTrp1zlyj/ZK+oAv18uzrm8d
NrHH+8Korub6l511m2WATFRXqChVefE4BXIcvFPPlOcRYALa8pi5StO7m4gg4kvtWZCn3JNhknvS
WdQXkLJ/HiBKS7lhdsdTfwKCe0D4GH8Wy1T9iqrNlvhAkIcZ82aXJILQPiX+XtuDvziLeIUe1ozj
dgNB5MyE67fr+q5yuOttOzlvx7T5MpMJ4Uug1aBbYGfGOKqccQES6uY3RHV6XKazXX/7/ufyGFCu
C2T4AjOSLDHsSITLx7CZM5KGCrGI27ryjHtr2gmKzfmk/AMWP4W2hq1ThjcsE2zwP4Cqwbypp3/8
kR7JCcbXKkO1/e0Pdg1ey72EPBxDRYkTkBNf0pnPVUb7KICoswRQOLTRWlzfaNo92nGMe9wakyiF
EUpAF0loxpw7kDzwXzNV8wWuLEaaiPWVz2NRhFtYYCQS9MVeH21ern64Dm1Fb2Re0xY6TsGGXuQ7
u8BYMWCzbnbOQN1g6d0be5fXl5GADN6z9sX8Z8lpDPzg8VTTuDjMjiyD+Qyoo04e0CZE32DW2Qic
MNS0PF393lCgDyg58QZLC3CtYwWvsyBj4z39UyLYngn+E1Fi8sLO4D2xAuSvcvsTLAA2JeSM3pCX
XdwTfD1F302kQa9qSRDK5tGFRVYMw6UkHfdhXeBATYsicRfCSVL3DFFYq09rxp/7dbhVXwXxhPBt
tc4vlVASJnGENc7mRAqXX34OvuqVRjStBEnxrTKzmrGtQQ0NU6eczsrpLZ8mgV+pFqdQjWFwGz1h
xUA28315ks+kj1YmSuyu5PSQThBI2diu8qcGdVUK7dVZ1gksvbm1uPbA1Stetj8uhDAdRkKMq3A3
e12l10vPHyduqW+MAcNEu8YChmDIiLfUzc1glR8VCJCRuHNGFYFbBEl9DSOFaa+VjJT6cyh4Fcti
ayVuTwAlgIFbDdU7VvJpOd+rroYVYDvrmzODAt5kSH09FEAaLZYA9aF1bCEwoISjrj3Wz3jV+DiR
D3xTGxK7zhRLb0bLMkICVqMISttWSJhiokrRcguFQDQJdyJAHvJ9pKQeTNue0PfpkECVmvJOcwQz
LF8nI5IvgIapoFMMy6HButfsscz7KBVgZDOqzvFO70850k+4EUvRAF4yH+JPyK4OwgGf3jCsCSCb
KaqO80baK8saJiYLuj0ba7UQvg0BfqPUaS/GRymwFd2JNf2l4NjNx4ywKPwa2E0JskwGUeucEk2E
ZYS/RxWXoL2vUeVcBwtdY0eGJjpOzgOqnvFay79SIlw/f7n0h7IYpq4pSo3njad/c1aexPIss5d4
kK390DgF4igMOYzGIsFD+BCIufXLLxyZrzIOFjyEls4ZxyGzwNI4uHkKytt78SMr80uBiXg0JF3H
41kwm/8VKDbn95pM0RLk0pYM4FhZ6XSVh/h1f0YwBxzs/BfzpbidypPteingpOnPIXX/yxFe9L68
tS0k5BYHXIR7C4JU9Wb83yREaf4g6XPUvV15Ql8wsz+aod3hxNpdDn1tle5Anq6RGQ0weM4akoad
Wjsi8ZQdrfO9yMKDvjqXwdzLAxlAt272SA3uD++u4crxfEUuhJ1JlA5qsmSwzi7R3x4aEQ5fQ1n1
seiyUKIYp/GUjFHQuSjVkfBJ3J8fpPtG0ejleWurWQXBYRsFZuEAazak7VJSIyvh5pI5bipGEtOX
4pd6i9H/0q4UTypfoxj1cJuXGImyav3aEHsgSXj5TIFLbvAYcEv7quimIH0k3bNsxyR3HOVshVTi
6/94HEdFK/GdlXe7Jwv6LRjwyR7p1M5+Erouo19HWUxvpaPQGC4iaxYkS6Co96gaTafz8NzRQbth
mnDdchTs0PDzCMotffNw0Tf/J2QTGtUrVS/XhlNRUPoT0IMGVI8xfn2YGNXmE/u47+ST3pFdsl+d
iD+4fsecN9zMnWudea4J2Fcs2u4hu6xfQu72XyFdEjDr9RYyYShUfg4Bwnfwfy9QhMTJYJBE5jIB
lRDa7WCM2GfUdNfqdtkeGrgAzQT6Ixlv2nIc4v0E+Ig7K4NHl1IGWV/IgnF8MN4fwcpmTJH8Ldb7
Ti95RPrvygsoRUN7ySOgSI99zNchwhrYv3KdYJL4y9bawPcPIEvciK77x8fCxjjHn1KmFsPE8v2P
MX8nRoSSpiBlutC7GKRE0+3Oa2DVsmsF4HBsKCQRX5EsnS5eKv19xva9C/IAbwPG6DP4L5Y+bMop
pgMTYasdY6+IU8Lm5XxbcoVCMe/pxC4tDwXlGqea+dT/yB2RxpywEVTimiLSPxXOfj7BiRRAz3Bx
3UhlrtgpV7LersFMhLxas1JXthXUDCLgsaHrGXfQiOXlE3irg7COLbRLfvFZF8Zbb2dAncxsmmX8
b5XYZBsdVCbf32nU4q8+hYHzW2RjXBgKdB0bNm6ZppVuJEJgWJRCfgOJb/YaluhQtBTLNU3cZ/jq
rF7DlR3VzREh6Y9Nkk6M12+6ENPicyZJoPJEeY6318iKIW3oDafIss6HRloFtwWMjDsQpcbhK9wk
41MB99Fbe4VyulJGOoTxR9NLTwdM4+R//+QrAHdNwS3By9eidzgDmSVDP+brO5jrfKyDBqW4uUgS
YZtHlX7YYMS/V2L15Q7/EGtwFCSGzf+pCwCehyuA1o//Yjpblsp1IhH1e8n59vp9kBVcWtL0l77L
A95bRCqnVYbtz1ZMVDMtUH08ACos34wz4wmW+mA99f8W2wWIS/IDEnoccvyws17Gqu+c04vu0KXR
91sK7Q+/q6jV8K9yVrthaSgRoF3zwkTIoPWH5iMsYZoLbWFxkpfILjbVOy0qqWDEVgtEW0yLrnA9
5taGlP7E5APIQeUi1rmXEBd1tVt9tHdxnhSkfeOF8Uv0Rz98QbYJPiHL+7OzaL3fO9yC7HkPHbVu
pb3LSS+aHtufBYtQlgUgWEwoNgewcxZQevpfDJncD1D1X7cZxvUJeItwulC/ZJX45d8vJOvx7Sfu
mLUFOpBkVKaX4Jb5y4H9LZFNVqiGzC2oF0U8SgwwNpZOUZL8UsM4IzQucICLcSlIIAACTnaKTR30
/6ycQbFonjF7Gin4q6e1HXVF3ELP3noNhpPD8K1HOH5KgYLN4q7CtRBLahihcSus2hMgpA0whR58
QUDWPYHl8wrYQbs3BqED/mm1Rg4Fj5vavCNZsQlIz5nyPBylH27nKrB5IHtI9xp/gqfGwZJqqIGU
tYfZKLynEB3SY37/R9KdvpUPNpSYfHwAYmkd0O+yvT/m4egYSTetfyprLkDwD+wOQhbEcO8F21vr
sl3yFHhoUeoPwvO3YpXnX1jL6rGA7OGDucph3sjoYqB3Vco0Y0UcIzZE34n2d4rQm9fWEGLWeyU7
b2Pu+6iz7ast35hU/q6v8N7OFHobFqeGg69cQ4y6wdjEUXhoyualX8A9PG5Z2RuGre98HArQbuH6
bz15/eiPuWYxUlbTxYSSwsraRyFXRp/ebm9n0rniL3biguHLLjnhJoGM2p9JlXD5Fe6Uq1kym0AK
8ckjhdnpIOHt4F6nTbTN5pu4VzVfl2P01UTcWdNS9hh9IyNLr8nVEhev5ZDqmMSHnrNDKvG0mulR
kF7cKXvjqIpcLsg7qeBYnFADtr4+pRI+oVTtjjrhUNMDe7ekCXf85OsrBIBUrxLsd92qV2zwM4rY
xJjMeTygxXiPeU5ASYerFkd2rIzarz4MKOUYwuqt2iT66R2AyRvifWP7+Uc6fNrbhfQGdvgzCxoQ
wb6I07LbrTICdhVuPhssfpe0Y4mUpa7IHbx6mejJLg7FBnqnE7qV6EHdqYSmzZkeB/oK3KBO2Pzg
FN0thzcxp9m905ranIp77jsAUuxz3TcuHdFEJEdrvJfkQE3oc0jsaT6GGTjIjBGliPB7hNWxW1nh
+YWAnDMBF8P+FmCyVFD3emMAiBF8KO4a4ZGg9uAESN9hXdc3Ap6ZhziFYpaNW8x2UxP1sJ5u9cuE
BCVl2+3lkdCj19nMMxzS6NHUyvyP8W2OlzuIsAtluEi1Wnr5w0if9h2M9vPtURnly2I7om6Auf2z
3RXTMOk188D9qNFjZ5db0q0U57xeItd7TI+QLDdaLBwkQ15KTpL/9SdkJwL1dKJFcvJ02g8m9iqb
03Ip5Dyfi+0NBlHuXxbbWOn7kBmATvUOr3YJLNy0OJD7Ih62iSQI1aquhJkJZKSomnELaYDPgzlQ
uYwi1UYG/ow8yB415uF5bCmfccdtOJ3iYx0KTTa6Lxb9DyREg5d0SJMUnXzL3JUDgkzuTWQJ5nVu
TaoUxho1zxT0CSVxhDUPmV34svExym1l/D/Brv4zTqm9zW4vI8E0fHabFYQ77rC32k0KRcdRk7m9
7CfjEF5XAXpk+C1n8ptqWo1uZglOHKi8AvG6alv2OX6VPPCKjIgJBl+BnPyx+IFDsAlIOoMSFz6E
0dwrs7qEoN2UjLGsz+eycHHG4rDN3S9UrwHT6zKGR11wWH1XWOtqO/dJUsRbqK4GZnA66x/diSKF
+Qos5cA5zhdAve7uZFRiZ01UJGP1aP+b4DbX6NVZIug6UL/TvlAl4dr8+8x4mGl3ISIlE3TAuP/q
PMKCUiyluwoX6MDN8MrsnPNuEnmGlP5ceQIpUtk38nnxK+cEpG6fHOnEzN5DqF9hQSe5Ao3FjBCh
iI4l7BCE09npK0KqsrPDjbcxQ2cvpOciw6fX+36msr5gUvvtSLMah3D3OvX/wlA9Ov8IrssGDJhp
D7crPs2HrRMCRGCxcyp5uuhwx+Bx6A5X/1nAoohT6GPCq9rWH3QX7KM77pgPpCgb8x6DJLOKWGqR
DSxjjCAvPcEVoJdFuIAEtXQETMpgJq5WN0Y1zjJVjERp0OudGbw74J7I8jXAhYoPo4WhYBsNQm/2
8zsvax9GdPX7Mx5FGQlEe/NQKbXJFwrkfQaFfFBCBpTIx5t/mXXkESjvCsX5rugtZrwb4L9JFEwC
XGHOa4iqy/e8cpTBxUQk4wnZg/6TTYE9VGaS6cq9z7LE+psJZQVNSZWtTOkHx58BkzoGr2ZgsgI2
YJTp/gz+UyMfsXKzf9qg9cTSS+s3sfJfZqme8y4sdK5LSVndarLpxIYykN202WlaRxB31IHAbgYg
9N7GBY9DIDPGGwOrabpE8f/v6eAfCS9puL7UhAQAj/EzpT8A/X+nyVD1igQUZ1WMcLs7jcIa/uNZ
DVqODPstZ7E+FjEcjWNrHPuZkShm072Dz+W47wqXQ9QHha0gUtl+cawHLqRaRXnIZtHIiLNz4czK
zLTTZmb976DrRYsPJ+quZYXm7I7NavG9mD6D6YSgcjyE5r4uS6bX86AuYmS10e+lB4V3uCIIjIqB
vcTdL18DQxboIwk5BencIawbRxwzgs9ThSlW5XHA2rKNbjeNn1Z+t9XPHTrOWMHgIO4jBSh2fFmn
Q9OUuAH5H60hVJTYtH8CsqS0LJbHc2V5ysV6sJJgbBQxEip94yOox3mSC8a9RVCf6zZf154zGMU2
ANOHWCtfnuDIUmqgl/gSWUq+tjE0mx6SHYRpWBMV5cgaouLBvA+LnuAgfcg8IN7lXxLtzY26gCD2
nfjZKO+MJOjevKyszksdwq+36J9TI8Vq0WkgKNY8OTZ3tkok4iVz1D806sbP2cg0t9QhW0IVSjgS
EzuJNgQFtjacJEVq8YLVQXa2qXrdaftLt1kNW7dFWMfCnqPEEqjUIS1vHQMtUSQLg2JC50S5uQMQ
KIyKJWmgE/3i7cOAZr0XKecEW6wj5gOy2n13R9ulaj3fR86feVV+cc6iPn+CJPMW30gfoXuw6i46
d6Vzjjw6HGzvNXPrcqonlGt56WSETTzk/Wgqwd9ttVafhhxoDfjR08/bbIkko/5YHTTnwWKn1asq
je/iPq0T+R7qOA4uksH+xpQ75MSDICV1mZhHVDukU482k92qWcaDXnGO3xXJ5bmjA5BxILi772yQ
wNWHJqnMcwISIwCsPXRA9MzgtqrCnxg+kKdkl4NdPuI+NKC8zX3b2Nkv9/X/Bu6qeyOukvw2Qft8
e4+8wkeDCVssLcd88aso1niEqAo4KyIUy7Ov3GonLxbEfbs16xLayey/5xxXLqrfb9ne6E1iHWkV
MOB4hsQ6dApKq+5lM9KkWw7mqcvkKYl2pe2g8zTtLTFScA8006lIZReC2fU/hpbxCJd3XHJjduqL
Hp4x70Dl06D2zK9BBGx0EeBD/4yjHehePl3QELVSGmRxG3fp2Q9/54T3gdU3oWY21Qy6VsNTl42j
Fp9AVGX722ZrXWLbc3L8ncyxSm10M1TDhAgckiMf4ubkbZVmK4D1/62O3jDM4T7TiOyCK+Mwf6gm
g7QwKbq6lXthKq9jeHF4B6HfahaWCJCjMg6NFXepqXBaEAMEfB/mUuQP6qHuhJN6HFMgrVUTutMe
BTPtVTDrHGE1TNPRhi/CMhS1S723WwD9w2cQTX0dgiDN1MGIXfr6ogji/RU2hhsEbFYQPpSfUzWH
L73JHsCUA/Af5dfkFOLcBWT70ayEdmR7c0Rwmc2j2j2zk/4FggYRqrjUvXo/zE5C2QUp0eS/JNPH
cgijch/7PyepNBe0llFkDp0EHzYMh3FYNNcr9x9xNRhVN2t5Gb+SsMMWkRatxA7l8heczXdCyfR2
4HTtjQIdT3jTrYzFZYQ9Yt8L6t03cPeY/f/3R78xxj6f4OR8lgPJ+Wf+Y1fnkXnjR9oEyHx0UpA+
cl2v8OQzPnBs7Bw7NHfOvjl/IplPsdeeo9m32r+9r6ZMh5bK5hGpfXOKAz6C5QKTuZOACqu6tsuV
DgzZRoPjamH1YL0EsQJ62QaYF9cFuR2wLdKzfLlLJNMRUuGoTbdcxVMywCP04RRLnH5cZms8pAPG
nEuxSdk0hEC4GL5M+eN43Jqjku+36HhJ8vJ8Id+V/5389KTimaO2h5UsFnLn/w+wVkyEdSK5S0Vb
riFvVTuYLit/4hHOJ1qtSTkNAmUDAfyB+TGixWRW35BTPCjoRaYkt/3d4abHvPqgR2tk8aIcd6G6
TByQ1c+sbyvhneN32IlC0Ao24+JeGj2ZpUv6G2x6OM7KMXnyN8aYYBi+9GbTkKdZZetq7lbPWmD1
/OLK5q9e0kmmSzUqulnNQpcDBiP+TMJfhupZgJMmzae2soRz2tA2G6Zk4IjKB5LST9WZWTkfBTCP
JQ/xtYhaeFbT2afMUu6Xshl6YO9SeHhetPm2Jw+9zoxFsma6zNIXI7/82WDhOU8QBqH+apXTfc7y
5DY+hMFd9MWsa04nJjnequcWi4d7NElNXOFhh5f97dErQCQ0ZnpAc2sgS/PSAC4aJngSM56f2rBg
FSbB81FinuFfR8ip6+drettCrlOW7bsjAOlxpwM8LCq1XODk+ugsONL55AM8AX1tIDRCQVpaJ+DC
1k+xZSZppkzl7dT+Ws7ARxPVe1KhHnxh0JgtdFLZyXhK3zueNcbOZSlDhtKWNnVEtUVjjHvwe73A
rZkr2h4yfreGSnxDu7nKOxVvOU19WqE/I+Rh7NEFFobNSXTD6kOewrm5IFsfpKeGZBUQBmFVtRDd
yoYpZ1uR0mI1UdTB76My2dNs682kN5IgMu/P2w1P4hHDUAQKM/jvcPeUPa8kPq003XwqLe6w0i04
lOqXFV1QnZoYIHsaCoePAY8usLb/dMW5dMFPqEe9dPh+IGn4oSengJ8qLKyjWURuosQarGV1kBja
+eHIVzVWTv6IyDSAD5+BPrYgsgVUkB1UEaAGOnSRXBzbkQm10OaVAbb80Rc6yez2jtcZiu/AmLCi
V0thxd8mXyAu+cvCFO4Kr8zIYaVD/2n092WGc63P1dDaWeHfUVRijc/Eg8NG+1kDCy00lobLtkbA
sOwMVAv66A6q6qd3Mr4JZ8AMDpMMtEsEOJZBIv3wSVlE/JNgLipRNxwrdMtG/skfGnIHXUAKwG/o
gg9wsTCoV7Ohudigv1Nm/uFZGiG2+eXsFzoj1RlyUkuaeUnCl8IJnm5uM8gP0lNm1wGSKBwL+nHV
4EVJ2mlYNWBDBWrZljwjjoXUlRBppk/h4QS2PVwX8VZXDp6PfBNcBxuxuihpMO/VtsPiLmNA1Djk
zehVUrknMByazjJ+UP0ghHSd9lR9MqA+lPWtNHCxifeul6hWNsz3PwSMf1C0g9Gw4XuIJOJMhW8t
2uiv2n4ExTr8QDYdpYAMbIz3gvqFtP6d6sT7VcO4ge8RS+HEsl2QzbQJqn/nLyVUqOZEJOtgz589
p3tIFZ7H8BWXtFoI+CKqmtwlkWeCH4hhcPUBjEryhPcPTGpbw/JEUxSijmhRs7MphEOOe6MS4sVO
iuh71ngGAyu9fpTZ3D4HLSUR8gs25+1iu3XeF9fgFOyDCKVVhE1Zem2PlRrhMY9YVwEWwpii5bQm
aX8bHrDzSF8Zc1z/0B86iEOakAMOT1G8l+V0keujk3sifqrEzrd7VwVpPQxTws1BaIcBS2woXjRt
4GMRKZjUIb+HjcQO0Jm3veJZd0KOE3OTp3jLwqH9LXU3GZ9sE7Uj3QdtDnGZJ9R07crAFTXZvBWy
gCFYEdtfXTzxfrPGgcx8tNhymdnQ12/+lEKJ0D2t9rVJPIeo8uuglLxDprOVeiqxyC1aqFz7anJr
cvGH+5+h1pkiVD9YGuVWRVBmBhH1N+97IWkQ4E2dT1RUQSj4c5oZa+hwlKjTCI3i5MgpbHt4XNvW
o8AG2XW65aoVMAtAu/f75PMcSPSryke/BxFyXn+trMv1W7hmA8i/AwvtDOklREfAzHrNsSyaoykC
k59yb25EnREAz9pxb9Q5ndmQKPgXv/uOnmH8EhCe2rFVaptDhZdiIeWnYMNdqwwMrRFDmAcEfH6S
ZOvp/GNJ4O18M0DcausVSIb4DxAhBa9NiLGi0QxhoxvS4N04OdbLMiEoze3g9kDSSkgJsf5mYNup
1cXoeBc3AgnpVN+P7rmbeHWggkEEQ4KdhBuhvg3oie/isvMN/QVsS0ExqlRoMPpUrhJDmtCrHF8z
FToL45f8Au21YrED/xKUWzOUbWbaz9tLJxU605cNxPxXrNogRAwcAeNp86PHOQWlvD0qKhR4RmJI
Z7VCfN2mSeK0a1+0WjUABMZLyjXUadoEx+WUEJ+1l5QfWVtKNpmXK9/HzvvySG+ds6zfwAiz0dB2
22DSfc7Pwdk77wW8vgh9bGGZ6fQ5Ql1oaKVaMyD/n7QHdy6rVygJJgUfn1b/4Wqzh1LIP7GkIddm
ye2z5aWcG6eQaCdletzKMcEMcdNqKPaCGre5RIxoSrDbmGuE7Bp/qcOi2aif7Ses+9vDz40obmhL
Bc0uWJ/w+MlIGTHRUHLh0HmQb38HYqkddYVbcHvczaVCzHJXiHTTccHbkVoaWyqvtTq9Om3jWI2w
xsrDEutV6OE/fxAaePnMLPP/XC1v7/gJrtfGOLxU46dpx5gmQyCQnSSJUP2Zg7/VXKXgHphymNJc
Ek5GgbYamDVJUVF/s5eTdp97u2pfDGtb7wUnF9F9jXWISdezXV7BLZMZhrcvDvxGzGKKuhRCpQzg
/z8RGPxY8TUeHtV0mRhRWQMZ3nlare9kvOPrCMeXQgryBQvbjOVIkeJzPcpFzfaOeGS91OBGkF4X
hq6aBtsUvTTlRzSk93h5gkoe5azyStpYBx95+6aEWnUCwPs8wjCZ1SUOkz2YGZmuUPhkDTWUS5Yv
wSW5GHgeXiEQNFEHBvoOhuwM8qFXb5y/J7xDvQO0oyyfXQrLS56jaYyjLTGqPSLlT4SN7B2UvtEn
W+VVR5f0OWcdqAmrydgjSMyeJjkumwxnHNmf/v9Drko4LqLAruB4wYw+MOQPtyyIRCSaIZX7J49g
joOJ4CayJ5+AA9QID+MiPOnsxLSYdXEM50LzucQfcU7f/4QGufleZX+Sl9CvpgYWsBZeQVPNR4PS
QveELt7kZYLM7biSVjjM/aeW2U11d7VYFSn94lbAHsKWXT6AFVOBjqRP0+kyPPtoKKdNBYaIBLzL
k4RsHgdIt49erB3n33YsqNiNpPhfYgzLIxfnkEfxOoi4QFc2F5q72dgcIm6nUNKY/6VdoHq5IDTI
QnlaU9PjQz2YniZ9BbqkCKE5bG9DZIxqH4xe5Z/dhW+XB35kHV0wQNgyq0/zeC3UqYnjje1kKVQu
zm/+yZq5VNe8E3XxVURkRiCiOwW9Hnyi68bnWjNXQcsxEkIW5E3l0RhyAmBsTRe6yh1S+vciYFax
WfrYChZHlJFtysgkv5XCA6eBm1lW2JEETUlpazEcXjJeFR1NHnCFBMKgzxNOdDGsQhrSy3m5pD4L
dMHa7TbIAK+faK09dgmSaNQq2oeeH58fme1AMXJmQJBtguia4BpEx+otnQS46SnIa4ZXKAvKAa2q
GkI3Fale+TafnQjuKev/HQ10O7lGSi+DlqUs3iNrii1Gcj+WcuvwifK/ZtYfZHhU8rgEYwRM6+kO
hk69EhAGdQsVGp7+yEhrCria3BCvWJqcmdYFzsKDf83V+eHX4rpBbUQfw6+F8pWQop2hQEgwUXKH
hWNbKSHuZW5K4bs/Ner9snpyPQ+dOL+oq8GQVUwbaOZvi3JhWze4v0OB/kP8GP1z/An2Dhtc77je
0plFlJ7S8yFabNOSwoupWpExKnRxtDe2a8CyB5Puyz3F5RgmHpDRs2KHhGVOBVg0JwHzZhazdPvg
CYlwKXQO0vPWpmFV6ZI4SFogYa+9Aq4grIBZGdyJsMLg6zOev9PVO5QEWAttiSpkvA08TsF0Uy/A
PteCVlBVjQj9e23T2nZ1e+L2gGlrWAEe2l4k+2vbsuGL2k5YB2UjL9fN/JIlv+TSd9r3diNSJFZF
8+20z+91dhMSQIuHc9RCjmuKP9RfNvLR2DVn/F0+Cgf+Oi0II91AYY/uK35MX5tqW48B5fMzH4yM
ZSR7cFcjdiA6+qEaucqhztTOkmGiVxlmaYl0zgRT+xhbBTCVasuQAHSLFseBBqFT6tOsWJysby54
MbXMCQmGF7JwhtBkPBFtD8ZksI6fE89cTBS7C1VCvtZKE8ex11NdGWtPREnQ6RQGT7c+jIw8tZMs
MF2zmwl9arpeKWeD78pjR7hjLX5z5Hy2nvP4F8ZLF7z9qIXOjkJCpd0+jsOTyyMaQghh4ZDNAoAJ
2MJB5os9DRSC7qaSYyt7xo0sDCwiBJPks5LWW1rGdc68J9DuI7VXgPjrWBK9Q43aLKgcoA2uLW25
XzSgwXqh0NN6RDAH1kNsyxnesioux/6hwJ4P7m0OsHEcVgf2s7nSypko7YxoGT2kRN+MA8n9Qk4B
0dcf2eCJqnwzhcWEcUDMfclf/w0pdN2IGaIZA9id5zHo+yr6Ry3jmcCoA6P6eNYnDh2e4b1mh6sl
JFrmemM4f+plBvSHUtCUR3CEGCZDEKO2rnLd0nhXMOpRFJu3Nf4DUveavmNww7YCHlizwyHSpJuy
Pao+tVMuL0DdqXJIaOVlgQKiNei+o2LQsZY1Tx0jzZ48YvIWp8xx5jVWduJb7J0JrTZH0a/d7wL0
2Mu10dfr+7CXWbC8NXs06OyH/xa24zaVIWIbMnEvu0U6+JSIJNhncXr5YmPL7P69lhLcy+k4SWYk
/utPrBr3hIGPwmnP3EeUWicf/XmS5rWEwhF2K1xOXJU2zAt8JwvW5v7ueSy6I57FDopgdvAi6OmB
bnZIqlyCaGbbBMR2uqUSEHU+jQboUiIfCaXaUArNUdNlkhm91Set8cc51ZiIexvxmt3on/DolQz2
jcKsbjs9BNQKYu8I7p5D2d16ldquDhmIItQA41f/lKbnSK79I4nVFq7MjOFWDB0BSRINTEnDNCzX
TNFBDpYk1FnjRI05aFclLp15TXs8G4UN/Mo0TG6qsR+F+hDAVH7a2Rkul2QwMeEjWdd65+rUH0M+
9OHgzPsrxKzWOVMpxt+DEGBb4qb/2m2UTLWdZ+mhyj3bwPgHN8ZqLL/JijLrjOELRTiF59VCg0mk
o5bKUMia7sP0PdzcQrLOh3bh/o4dL2Q3fvM0ip6r7y9G5+EYZcWfom+l9dOVV79znDltlOVL7wY3
xchcbwjm9AnL+7WATGgjT7eH+s128OVuMlQES5ftCUXEOLd2sew+op6JQqYbWMclfawbfQ+fqDks
GbhoTKR5Ld1aMzTnf6BSjyo4gfuQ+aeKce+o/iBmdbtaO2ve/2UD/R5DQ2HuixlfYJjUBZcKJVkj
QWqzhRnSoHS2fZWIIQum/9Wng8dr/PzJ9ioDsVbgweI0lX8gJD+IPttD+wjvmhWvkT5ywDT9Is69
XYLVAW4UNob25KX2dA28xTCuujplkOeXmX+ncX56WsTiDlxPtcpLQPK4ewWv6zmCHBxgrWfb8EeW
RyNZIk95pCGt8nwkoPm6/2BeoIiD+k/b8pY9n2bwUtZID5vpdajqhT1UwuKjQgeWuSq6KoZSoKHn
JioIlmxorRDlPcdrrsHKEXf8Bw4qu4TviowhX17yt9LZD/a66FQ6LHPis5MrT30hBHR3Y9o1ZNHy
VWkN1lPti/yf3rzMO8htNDBAe6fLwpx+lnQtMhFo4ciVTTi0pX8MgAmpHG9hwCh7IFWHdOTZ93H4
apg1Fh70rSLS7B8rV12+kcYiuovyhCig88rJX6zYl6jFcUljn8+kILNvOErVksIUGOc171mjQzd8
oym0VEIA/BOI9OLlcSl1oNCGe4TcRZqogZa6xlWjVDb/iEcVxzIFg0Mx3fWRP5giVEvYdzDDaMNH
6H7x6WSfpnHoCoHBCI61nR+RIkDw1hEdedWvtfWYdqdIxzcCE050LyTxjpotgrGXyDzSlehJKdlH
oXnB2By3r5rl/m4UFYFu/YCA/qyCG/1hmXhNwotcmDErAJ2S5z9qbXN7HxOcuBtPCMiLgMO05kBH
NdNUe5KdL2ORflNP3hz0dc3zjJtAGrfQNoKmpFw0iFacy7+VYKXDjOWu//MsaGEcu5zqGU57bjGR
t+gBcEtFIC/KzFD/dyIqtoatOqnEu+THMFgLxDT/5s2w26PNX21u3TZykH4Lxh1m7K4n5b5b98+h
2+jD7huVwVekpdWHLLc8MVJaP/kbw7kFJiI1wtBkFySUkQksx9tiB32ceyJ5tLmysaHaCfQoL0bv
oKRf331rHx5mM0NRI6uiQ2ILj5h+0ITt2g4YjDlgBpT2bhh1hT4Y45Xyii6z/doHtRqwVtTLTHZb
2IR16kekwgho5ahLQeprsYhBBBLcb7wLTQLEHvn1tVBvLRHcQdVJmBKh6VsRamF3Y4RfGyliXtuT
Dio2wAA0vF85UMEazCy8Pn5yXnD2hJkTITtqG26k4trieCBi0ZBB6BC0B+i/jJ49jf2uQ+AKx88f
rqhe1Ff4lXebCVUVr43WySgl6W0CCxI86dIROFnnzy1zlinrEsLnAgJ7weT6p2H1LhF8jAZ3icpO
1zbMrTlar7ThPsq4U/vj7/NtMvY98zV4bJCKJJ9UORSywLa8taVfNqI48uDE5PjqJoaahj8zdUTh
qXGIQxkTM91U3pe/og/VupnJdL44kzHTzGK5GKosNGpSnKjRFkeOV2MgiitndEzGqZJnKzH3nHBQ
XT75PeouZPMLLQXu/BxArzUeuQjuYWHSeti8oZcOB66GeOk6DmdyShKHMreym3Gxpw362G/IbmBu
xFxJ7vFgl4TcHkJz2/1Yn0rfDsXE04DCaguf1s9y2EGfsMQEd7mQ2KmkFszj+JRRakOHafIp1F08
U/L+UMcgqfqClMwRajIiXkydadyHy9oHj7HmLgkGTz5yugxYQZ0SGFX6brydB2K4QB385yjK5FAQ
r8ZI++szhVUB8skNgiTB1aGKZ9Tw0aKpONVA8aZSWyezF5SKOJSXADEA4JUnvJdf3DQ7xBJc7l3L
1gwpTw6g8wXw+6k6JRmfJM94BwJeO8o1Oo0xkXsLETDI4BL5wdYQZNo9u527OMumpXG/pXRQRcsU
IL5Jr2CDQ9JgX287LmEI24eLeB2IWbOqaL7iYVzbyVWcMKfoIegH8fQrxEyVGa0nScoEGAYBIGZj
FEj6+Lb9GjdbUTkY8nXqMvzZehor2gwhgt2G2L/E5ZhjNZDBZG8KHB4znscX3thT8y5EN0WeyiT6
gC/crGM1srydsVqjZ2DvuNKATlhOyd/o8Yh1hWALGP/3bapsITmMOuOI9Ii6RLXRw61WzN806Chy
bcwK6qHyRAWH+wSulE//T+mXtcJGLPCtqVcEdNnztRTELHuJgyvNfu/LeW3X0aq5FFFKpKh56eyJ
E6fhbgYtdKYQz2bYTNCp5cZ8+Fa+F+pPqBNByn2n7feR/Lz6elJZ0cTv2ym1up7PUohpxtJexhau
/dyUrMEFjrYNnY6tGtvuc79Ax2ewuDk4DU4VZ5tFPxm1LKR0b+KsLmCfTfiCCKM84vlXYXE9eMQo
BOXYUt2lMV5KQA+qdH5WqshGjm9y5/c/gROcPYPtiwc+Aov/ME+3920pz8uHLGluUXae/shWTb4l
UAk6jqQjsKe44rWF5SXTfx0DmKX9kJ/szLR+uHKKc2q5yCmfbSkps3DzQz03Vz7+yJteJuOppLwS
ETAhhnH37V4dSi0TNVCAq2vTC2H9UhDYHODCuCzZ9QNy1rWucOXp6zNZsuEC4e9NGr7+CGCBfxyk
pXQhusuafgtDWcDIskXYIb6b5YFaDH+Wip4TyJommymTYWBfvs3ocmdwvRCRFkdpAd1mzyuy39Tl
79bfHPweGO6/VEhaEn8+VRE0WzdVadnZL1mWy/AhqB7+qhox/A8CaoIg8Bp7LiGbeUa9mQLzI4yF
uAuPlw0a5kagZuJddlt0DmrGZey+E11egsxNLFuKzBMShPY8vSNBThUCheQicgPlKOlSN7xDjkB2
pgDv9b5d59+F9X2bmsysPrjfgGF9XT8+btn5t22wMrgDi0rULs4uFXmFlkhnzgGaRbGkhSjOulzI
S6tyuf02YcLC4U1gF9rmuyiiTaOpPHW00ULc+0swsLSxhVRVlF/Gw5qy8ZVQ8SW6djcjgQQlMNDg
RzEafPG1AZ8lIZhOxuGkYv0AYlrKGdZWMq2uv94nQuF84l0EqjaieNlHFdGv20Yhwat2oxiuZbGE
wYKNMq0m1dqg/wq8R/JXfhkku2neWc1HdY2zEbQveAoK0tznT+6/nmsBZDh0R1TnLHzvxRSKrkdO
6JcwnLlopqt6JAwG+E9GKk6NAYR2XJ/QI2y4QH6cgPZ0+8tBxKwKwPGO+MWdLnt9r5X1OlDSzYSR
dtRioTyUubH/J3ju9vR9O4YDLpamqO5zdI1UBra0cM/jRW9ONwM1S0xk/xcNaE6hbigORsFaZ7S6
VRiouzYMdvN3UuLJne1jyc2cuC3hNUjV+zLqTcnsnmNdAdttcwu/c3ObJWrrko7yUhDfcteX8mhZ
ALTXDJz9Gf1h0b1o5NsJ/H9TQXgOmVSS5/6zSuMllVdzE24oLrg5cHgpRB7/u8e3kdSjIjXNrzsd
DfsrqW472Zv1NU6A6xm/O/HGUdA40O+EPYYIXqzkW0AfpFDzI1s3jj/K8ivMByGdp35bcQgAbqeT
ZiIvYKOFIrgH6af54CNTgXl0M0PdxXe8WOb2CBb5b/jH0Ij/UE1auc833VmADHmwb5sOkkW4b/nl
oBDY/oV5/3PjWTHhiJJ9SRG5Pb2ZR+7hptNVa+rp4AT0gWbKsa5KS+p79vhVUCR0GNlCdy9xI/jr
3Vw0l6lXWaoWaHYiqRKcHQSXxx61fAfHFdc0HUEvB5Xub5mQRXekUSw1C8Eo7Cd5rCVQDnJPn6OX
fZZ95Bz/3a29wqyiEpUtSB40sZB8WLSo/KsJBsmJIvU/AmnFvZsg06VEy04jX/51aUP84tMUzyE8
x6uvMki5Ua1uqF12YlIml4TMsWShFhTHwrx1l/ZXfafsAtzXisOa2r4Kn/sCDhqv/nNRtRMMxrv4
QZ5q7sU7wE7tX9wHNVuDVX/0pfBRP7KYGoGVxfIGOgKt9gXS7f9eWtlY4Ycr299vEU2Ww+a4vHFp
0I5TOxayQ+GQoJ2fy4B34sgCPuke+PdG5sJZfQx/sZeHae6PswWal5P6nUH5MIPZ2m9wF/v+oXc0
GqqlOXPO8D9+kWjXhFWeAVFZ8UJPXUMC7u2vqA4H5ztEdK20QP1tWpv1D4VgHjMIg9LttL8UE8bz
7bvzKSCvrpRTIDZiJxjNzkZS6tzVNJ2Z2ZzX2FS7UL04qtrZZxNdVwtRU+A138HLzo3bKznY1uT5
S7vZNW8y71OHs74WeLj7+N6UKCbOuZutOwRq0rrfUYrwjHnCC1uV8s3YhTj/mpuBv7NcnoLWjPkp
K0J6J9LWWsvzpybYmqGFhTyHaESc6xSzzjKaNy9AVwkeRgvBQMsEqoxIE3IxwqXOlt/uxcHfTaCb
2JGT51dgIHAyI8vK0vLBrhuU1Lr1y3Gq2lL/V+4mzsjDWnnySvKYbc0NaBXMnrcdbapzcG1AG0fV
1fDaVBZgQMZNHDQsz8vSphWKbiHpDE/lHp3m91bhtpl9x32SL53C3Vp3erCp5MdbqGYiZC8zw59R
JxntZzKIzypKsjapwZ6dK5x7soLIoYCfB8mJLkwvIKnF9C/eAVfQCeOVJaHwhsBHShlLrF7Af+dJ
wQqYASdHQTdO3k1eBsBrJRencCYcKkXxbH9W9UHXPSBLOAcdHeporal6CbBOLHk9MxE4/oEFyJ46
+1Fsac+/CRBDGZDCS1fzTkgvcmKSfg81uBgUJKKQup7ruV3C5aASvg7N7M0q2KYZEVOp327xyhW0
1AcQmOg4vGgGeShjX7k/4ZrV7TD+LApqAoI+WSkpCFUMIm4F40JFj7aOzFpn/QB2Wj9Wxj5MN8cJ
lyZy09o38XzKYGKFMAbY1FWG95IlLNarYsqmfMh8v2nzryY0CqZJDdHY7O2YZ7Fvcn/rsykEbkGr
4tbPwsgHQaGUF69xw3tjln1fdaL4rs43AboAB6qvvC99wBFzu4iF/pitn4TYh5YlcAPONpjeeDAM
Z6iEAY5wYFQ8EyNuR6c6tDAGYS21ui3s1uspQ9qPmsLj99dbjMC093YXVkkkdEAwgJarVVO9i5wD
hi0gRinthow3AbQ6C8T4H77jXq99rLLZGNjy0lmzN8EB79gsEtvAeMHImGcRmR4W7ud8fRPFyuib
YzXEEydTr08Hujq7u9cONJu5kCCKjzqBHXLt/KWa+AmCkm7BeFnrScxfTdoQntpKNWqCtWb40+2D
2l/v1C9Vfjm1tNjtoEvre4MI1q/KJF6FSSkZeOvJxQv3xUmnmLx128a0LvjGaqhZwB1Cs7nqCX2N
S0Cq8JPgpjjSoCFGRSG1BEERj4FerrVERmqQClaQyx/0ua4QdrSdxBC295Z8K5PCxv91qm9Wco6/
zpd+hLyQV4kpicDyVFx0CPkwWFGtx+oSzkRkzwQNWLxahMaFubzbcEIQc3D9VOfH+3dN+Yqc7Vmb
SwgMcry6pWNVLDSd9lxW9e0s/ZGwVaA5XEaeACVxvM1T63FB1BCY1hRSdsSlVp8CIbHugaThRRyz
99AMLgcIwgxxKsbbEQvLY0seYT1NaoZaTT0u2Mv+BZn2gL1cemcaBNwvtA0kaEEPSlyR+KTmxg+A
vBf9JAveJpmsXjRwIZXGuuwSwyMF9Y5x7J1XD7SlXw2SWyF7WZ6Wbk8NqFxZDITZV6N7SJEOUIQ2
YoEIqaTcxdWF4e5alUOwubY1ik3EIVdYl+Pv2ZMRHt52ZwbcgolAqba+3CJxZASu81lDFYAg/r4C
bn7HLqJMu3KmINPM1iWXGapuuxghNmnTiUDdNDOQhJJfk9mgszU6wvRvdjdIsXXiwdy0uo0x1oZb
IHNIFsUmCb6hskSPjxdQp+NpCOIYbBCUDPi2wb9esDafkg0oNOmWTvnpHxGjXJJ5t1ZT6O0+jmJu
eyuJyweLEGFAkinRv2AElLvZS2W3wPGBdfL4SfQt001NW1x/taeBuCNN8FnFXyLr+UTGeINIoDlO
NyFrL9QAgO7CEHkwu+LN+8+28Em1/JzwnUCXZDLA3eFCtW7mRScy0vj4VFdzUpkqzfl7nwRfyrZK
ql6o3ijexQ4tsRS6Bu4ffvVvv/Kg78WHK1Qq9YfiY+s4j208FNg4PraTGfUuPQSG0410KDd33b94
X6qpmXjnSPyDHSkkPX+F4Fo09m3RgiOf3Bp9XmkSGwPVjjnG+5Nqpy2Zr7ylNHvBginKg1YSG3Ys
TKXWHmYvjjzavNKLpYAUkcwn/ZQyjdARs41U1oILSe63VAdS8IRT8HPho0lO4bw76PmJfIovJv8k
29XGWzl6mB+D0F0m3+29D+Z5MsMt88PVAJ3ib7QL8zFugb7JTnzfXFky88tHQ/6gh7+fM1c59nFV
mhwO6+z2TCYgL7uEx58NtTvXikxODTnqIeiMej6KfyYnqfLfHd+phfb6d/iBVuOrMKR9OLxgAbEc
t2VxEimKeSh3qslMQlFUHvLTKu4Lp6MrOM1TxFyLNgrAF5ODwtpF8jnG32OR4lRql+seSxSNzUmf
+ina/RAW57p3WcVU6K/f35hV+gSw0IhIpb1RE1ETZmwezy0pNcFvBejuOInRFKbhY42rl/exUAW0
Jx2GYjpU3J0bu2tiDHaLRrYpB/yPejSv1NAck45WuCOSVpNl0upW7ctfh+G/O8dPngXtZzZvjYMs
jvcTqNSACWCiSlMhXKHLLUP0dcwLARmCORGWsEkkFiJxiTVGl0LlmMBn523AUNVwbQk5AnJrIlmL
Tb6IgOPurCHvYxYWxa2gldxk12SCHwUhHcOLSkTw8rlqhIWl9Ybu7kg51Dmq4ScKtNZjuaC4L8bg
ybw6Oy1ye5ACkm6hhNKFKmMFgesdREi3o6q5d4VUdjTdhh4R/er1OE+oNgFwgso+rJo4pdRt7SC0
wbTJq+rP5rvXcQDVoXSZwqGr2YofkVZYLfTqhFqK8vn/ri7yLeIPWlh1D1gOKzrHFTVRLp9uiqlL
YVaGyr3Zny8Gzl/gRNgf/FRYTmO+dl/ptFXOViv4nY95rsJgLF5zNavGin9Vmnqz8J2A6drDRhYo
EdDpaFDD+4nNnXCyxEmgS365qClVaTZHs0MQLVJfoJPsr9r91+x0amVdOYTvxciiSUkOOSx4rRgn
Kv4/z0iI7re+UTBbwDYIGfgkLQ/W0qzx+un/aSKW3fHkFGW91YQOPQSG8Qf15OdrePO1wVHHs5Q1
6ihHnHkgslV9xr/C6vfZyfJzDBwGbVMuGcCpOTXRkw/1BsAZeCmOzpHbRBJ+diVNr/qJpEUIuwak
8HAmZVUqp8IUO+jWwWoiOuQ+32/QZ5q3c1K+PwKNxRzK4jayJizfS37gpYWsK1XA71uoKhkxCTRd
24E2z/VmnbeBRYZyAMFy7kMexj4etaN/M5w2UPqUrz6UKuWh1Um6FvY6DtZRns74K7tJK8ek04Aa
j1MaTDaIjXS9hSnW7GifzUlhMPpOP5T0bKIvpnwdWt5pWuxpCS2EifNQ01rmINS6VPS6STmHNBwK
2aVp4G10hHRlsjDAcWN/XlqBiJ6mq2beN4MVxV6PcavhWlZJkmMlrdtTnfUH3+o1cU92sucVJAn5
mb5fsqVaJ8vxIuTOo2UXoQoP3V1lKssp+4HWmCPb1HWxJW68IuS9ja9waN7JpPdHQqDFwi3TerOH
VM0nKJKC+kU06SRERf/kH2Mk6C/xlpX2CtTRPqMPzGJz0b7gQOKnYLvyKoaWy7Fk3BgLTeYy/evz
FlTdmBDf6kBP/BjY11iTkm62mdFMVLwyRTZ+X+bFKljExHCKiYUTEPkTbVcdkOze63AU+XpJCVlU
FbThWP8yEOfD57Xb7zGHmJFbH+xm5B21vmQke3pdKN5IVRn7cSCdD8ZMlH/w+dQTIFYotFnYPUkU
UMpBwJywP6WQt2sSV2CL0ZqTmeExR4EYNaerAG7UvSAW+Za9eXBx1zbrOdEBJ9CPdeocOxTfZQ/c
Je7j+gYnR6SEzKQCrVMiiDOhhPEhzd5ilTCOckkwJO5tZj+c4JMRoO0czjFumcixSKVYJyHCUKCu
JZsmCsZlj5KQngPqQpEwdZ8iu1v75kaNONWT2AVO5aSmM+hgT7bpQ6ZaeP/b792OpYOM55R816R3
lSRvHERy1d+wszO7noGdRkWUrNhhoJoH/RDs0aNkpyPPFzf+8OI8c7jWp6+9reWc3BQq4Vy9VKah
7puWghCIoYTw85y1HZzvHLNGrAdJ0rML7HLj4c5M1/pq7/+hKb3CxcGuLzg0fTOgspQ6gh2GtNyr
0nV0a3wpPFQdK4/BLLj1zhPFvgqD/zUEWA0Tx1/EgDDXklg6GYW4gl4hwgjHC2tgEjPzYfRNqEG7
SC6jVJI6XOwKpbh2xhc934SddeCLgUHrvHdYWJ1wVWEtFhowEsR23jyACOfIr8V5FBMdVcZDYJCP
lfj1DJ4cacxjVkEWay0i9SiC6KIlCCHNUao9pO3w/OcmX1KEA99uYD+nw9H/t5zEednzlCyfql+f
P+PFJqYCk7n5hQppeva63R3rELLJtwUmpt0SL8z29Qaqe0TkboCCjvWz0ve/6H57XQwvdLF4Q0kr
awNqngS2owD8BesL7RRM0mN1GMaTFE2u9z9rEMZQre45Y9mHLFRqfGgzRSWO9Ya+zf5F6wzAXxoC
u1eUPf5L+270/uCUYNvhCv57aujU48j0Kj3gIY6XdeZuGdXR1OaHT4SebH0vxmbTVM8weUxaffVg
K/KNCDoqgzga/NDnThe791tmU6rPbOhpN8SxpyMYsTHkDegZKHix+oufMjcSpmIzhnLBxxHI4Jrk
jxSMgZamL41zK9b2FTacXMTuI0GtLUrRYoR2qHFXrSF4rBdPKg9+3MfvdNkDAUrsORWrDuIT8MTi
82od7TF9N86PvJBvLEIPqgtr1DdUX9g+w/GUjPShLORUUxR9reHkw0YoPWjGVC2qhDMXhufLVrwE
0f3zYMKpUZJEDoYvQta0kTLF4FVW809KiEAqlQImVa+KXrJM32ut/HRJrDEhNwToMUWSqCUakteZ
+7iyYSLR50fZ+PHz9m0dDrNNUeLU1dZzD+45vM9V6ZW/GpR0mNgePPWSi58px4vY1w98FAHrUX0/
+Rvfry8rp0vATzpxsjFMoJDLh+0xA7J7B5Kp/5fFguXJKYTH6cK9ZH5FoDAandLIDHX5m0/8uQJp
tnqfxkfBBxCvo7LoWCwxTsNB7IMkLrtkMMBznlRjw4tYCSsscqbfcNM1Akd5A9FaxMCdUn1AEf65
Yw+8CjNM3QBaxXcMKpHj/tewiSdJ5oXxaIE/XBzn1Vs65Vc61ClAK9dj2f4BDC0a0kkqs4Sz3glq
fjo0TV90uWo9Rt1maklAnaaAG7ej5FvBFz4zL8nyHQb1PNhP4opxK40FloEZREJEOHFf7rZ8E+GX
12OKf+WMggPkiKw6nx3IPVufclcS4mSyxbmowtH9PBxWr0u/954hA+16Wu9rzdMKL6w3gsQKhpu4
xd2YzcKdUvcoCkLdBhDQUMbaOr8J8pWTpMM+fXtViGTl1y1Uo2Vw5HLCyM0l3psbbEjxioazN6ta
e+lcQIVtV/jJDJt/IyCewNM7H2xXKn+VHII/4TWhRu/JlPTb73N6qJ8P1H27l5xTV6rESzRXhKLn
0T0uCa5ybUsXPDOMfaThWtjIDm+tHtvqPmBHGiKRY0Oj+spUvzN3hYIUNMbsa3ky3YvGCkMupWtQ
PDbduR74sSeqq+Q6yWkCFSlZO63l2pKFJG7/2W4hUuNz/xxWk5h+eShB7nYE4aCmghstdnjCybOq
mWc1pq9wQsUMirKjtHYB6aLyoXxQKnLP9aYEoZfFGPf9ovkY8GhOVC4jkMhhFZ7DVuXQsAwdH0PN
mRdWOJUv0SbaOJk/+ayK9vfcnplW9ZEtdvGNM3uUZE2vnad7UPltg4mBnu9ZFUy6LWEomIYsHIGu
XNmx3gJE4CGfbkVWObH92tcCrx9nzLnw/dSQaecSlPW5Q/Eiy5iXwfChAbrlj8r20LQ4VyvkFKss
Jx2QK5GmfLwT12D+T7WDmsu3fRrM+B1Cys5EqpaNUB/n7pYvJDM9Bxe291sec37B0OtjnJHP7kRm
xyQ9Tx3KA549TRZMxgvZhdwUSpo2MnP6jF3t4gzlBbinUlyZSQiuoe87HQOjJvRWEJIrXW8RsgGJ
OPUQoJ0P9auc76zPJoMu75qIL2gmjzrqUrtdBFMl09c3o/7keBg3Kdzg9k1LweMZ/o0TFQGfb3+G
+bUjly3gOK3m55hIP/2BaF+IXXyKDDUh77ZTxbN2y8xOCicyL5ujXmR7ZUjo/6go75XnSaAypQbU
FLTV/ati/F+fh9IezI/OKvX/34i5KQHkkzJzpz9wAUMQDd9WF5DAu4ZZwAQCJzEKtXnPO84FaNTr
MX4qKR2wSBvuJalpb6Y+W40iJ/pWW1lWzTTyLZCDaAlCTUlQ3UiXMkcGEtDNS1iXr8dtN2RsWk8Q
Fhlw7QQvtQJGrAGMO3Z94DGVYCChuOIGfDVsZYM4gIoAmj7ZqB4szyQWE0z9UepuPY7UkzQvqhrX
V11tvMj2Z+YygKU0NnkBLiGohyFm99Vj7wcfyTRTM7GqmNY4lPP81Z5d7FWUYUSXDgbllo1vcw37
2RvkergNpNbBoVAvW10VRYGB0JZrmJJsNrJapXXX3NwIQ5Wml1iRO9E/fvEAzscfkFnQTLNPAyYN
HsHgnEyPq4HTdEq8clo6QKmu3rcdRrzxmhOQRIsXzH7rWH1z1AJK3Iep98JTZvqWk6ITxCzsMEhE
7l9THQjmqScK0yWKEL1U2YDaUeOqbkx46tFNoRu7QNorMA3zlM2654dBtspWXWdKWG0zC42uwVQJ
dYkRByYkpggFmr3MuKcQq0BiOO8L5kznLGxdbcgBCxo0z3xn+QdIwjWUxvi0GmL2M2qzKP4Mmf4z
igJk0ZJKfXMdYzDtB2XOXJaH35B+re4jtRid1zeBjgDX/JQeT9NqeWtGG/30ogyTZqpPzyyWtZ2C
+TN/1TvYFkGJkYpN28fW4JUOzgesczbeAPsP1CP2mXW2Xc6iCN+QqzqkkeSh4sX6iHzaoD0PegHB
3h3kBvFQJf7lw9d4OVwhcbehnCuj/AcHGs630QZkKED5IGZGlENnDolf2u7HUzoIePgqAoyoOhNE
y8NmHdH1L+SAcwXnFLC+x9LYTN5euIC7D7NO88CdmvZzzp5TriRCcg9EBbYoBU6Z+AJbDzGNpwwT
Q7eK1bzvisiDUmiNc1lDnIgVg9nO2KfjLtCWWiYX3cKoVImblN5lOvPaMQwFAbfu0mHtj50nrOOZ
HXgu7lfPE7GUUULdSXTNLOMHiioA2Ci3IHmjte7LmwLYpwK3NlSnQ71RBF3LQo/jyV9tHiFXVO+E
Thhjuak0lTz4lbAvr+YFfXjS3TtBg0ANuuP4ESdaMMMOKNjIjLQxpdZ74Thxl2JR6E8osNxbAeel
TS8R/7XJIIb9ts+OGSG/jjMa1pXnbwjqOCJ2PeE3GuBYelusTZ6y6MTxYrbvyQNHffqrIftBRK6u
xnGphDKc8l6YNo+M5FaK3S7YktOtzBNb0/Hd/iczNehEFlzeJ44Zit2qHTbfrUXggWizrgEizuwJ
j7BP54M9zNRDOkCZLYyfY+HqPSeIswtPWEPBeQpWkCGqEY4nFSG21rZ4GBIqaDK51jQ+MIuBl8YW
CPt4NGjjXxn0qzUpjacRKcVS3HW2vkcwULM7gqC4WS/zqxQ1vdmbrRyKW3G+O3YedNAGkgGsvFfc
Vij/GxdNCC0OWuhP6Ob3n+YRhzfTtZxE8OIQhT2SVKyuZ4VoSYn2Nz/xupH5+6msaQZe2BxXwl1a
Bhl6eidxSHXil3BO0vR+SobOK/AQ15XwEYeB77VUZwIXhwIrPRcB0S6xez+dl+vQlcd+0W9uMcmu
hc6cDwrgYs5gx57sk4PTivhBZUPTwp4gaBZRRbF+fUQm1fr12tiyi5O1mHBljQFzlPHBSfAfnoRM
kh2Pm+3qVhxcfPcrX+Y5qNdPyvcs4KMCtTgHIWJoKBBrs2sRWO/YqFNvKPS4Ek70AMijQHyrUS/6
Z4Qa1KMdgZfYHOG9fWtvZZ0lDWPe7bo+ob8EiuUZhjQFyl5+lAoGQ/MRowyowk9cgSxjyfmUzITi
3uhVNIkItCiEAz52BrmQPkk5eAC4p1sYA4z6VEYcxUAqpwv8EgPUPbZCufRqAHhnTa6Koq+RSxf9
hhvDp9pNqw57oFIpw7wEsKx/DCAMoPWqXpvCFop2aUlJEgZVUZmhHM1aNtpOqL2V5A77r1GSqAXG
V0Nt428+Hm6HRjlWWOXyYI0Nia5VPSfwTvScvwUVM2c1mi8iPGSFSRLBHCv5EFRCxVrwL6kDL3CJ
sXojRrCisBDquFtc79Fi55r6V+sig/USrZ+myou7rLmPjWxcS4jJivp2/J2q2ZBcBYJ3CiJGCHGA
bwj924S2JdqkMPqpzYHvNFD/I4UOOmdd6RGJNyAI2zI+vy254fA6fCSQbO7giUeVEE++1cfW6x+5
CnviNhLmyWkfNjHZWzXYxDA2Kt+HzD/9SYZypqFQ773SbK5teuiOt/6rGWtJmEy6SxOfXr0suasa
U3QK3dmmNjKJa4luNGHogw8o/FJYsHz4QSDztracsr+0cIUQKkg/QkiySr9iU29zFPMZX/II6/vg
2ZrfUr2HtHKzC3dQVNXqgayyT/6rNgBOA/78dn6DCqWnk0R7ykAp9kEo4ThaMKYNK8mszzGeaOAr
0CB5+2xR9YMW4MlKwrMfoZZS6wExCuttuNgRhiQDZG+yMFzwMDfhozT3wNKvarpWGfJKJ173/8Yc
T9OfQmY8A4u0szRyldBvMJuyI+VKjcwpibJuto0YMYa5nqiZKDmK0LHtFIkJ2hUqnpGI0COh1cve
RvzQUC8ss//x/oljMjG2ysyvltyho+jc4JnJVuR258MMWFCXTARSpKgczMDDtSSYOJwwqkCUBbBi
JOiF9V4e+iWUHkgMzA2BRaT7GoACN0Yg9jXyZFJb6feLYKSLNe+wpXZRrtFqLM4cu3p/QsSXg8EH
9Q/3tbd/uUV+Kb4JHlJEtHLJBtgQ0gs/7mRWFGLpGraB7dPYBLW0YKhyxIdYijgD21F8jdEiD/Vk
oW8yhs2y+cqsCjLgybl0TpKBPEYypIqw8amtbhno/E1R3yXD68S8/h3j/Xb7Y3s1rDAGdyfq0zrH
UnrBZ52iUOYG2c5Jwkl0O5YvrRWmFXkVTtcD4mNvN9zPl0rMGW0uimSRs0QsL5jg+9GnHZG788KC
mZJvgiVY1aqg8h8U5zfqPeof1llJLatiud0DK/tslOIDrbjIIViHQjWcs49RcStkZwVP9Gaz3OyT
8tCSWUFhY1EmU2VLyWROLhMoglkMdImqYj1yXtJ+Tg8vYwIRN1WVsYfle+PJl07CfYj8skz0iGcn
kxEqevh3IXBm3QUNwhGxvKhcUjwbHcl6RN7FGZ/9f0/y3y/Q3Zxo/uHccCCfPfxcFOB/H14hyhgk
cyqbnD5tDn/4chlFpOl7+964VjMpmJM2/pwZEojdUZU9bacXv2vItRJ0DEp/MJTduONuRvwTrCSm
TMZKIw9iOXwV6DmD0DkuqQGdriVG8Izkx5ncC52D2vJMEvsHW1gd+McdQMULCX57zNvl/Q5hg6O1
7fVu5oOvQaNFn0jXW9Gcuudj+MKqTWZIFbdpyZKhSmSdbZ/Z2yGMUV+lcxASIif8Zyo1gI/KxOD6
ad/Qm86LkHJ/IpvDOt9KIayevxQLtUHDDxXw4uC12LOUGFKBN/GGxI9yBDKNlSFn5J3dngLrB8sB
BdMQ268LB2hna5m+0UCAfgBKwEPpOBQACOCT06howd60f1i4XUDqenA0R87iwlSJu871w6LOjjt2
GPwhTKbdltsElkeatiJvdElmlhu4syHqN71Mx2cGaqBKDMOqL0wJPHxzwud+Nq9fyCT3zd1pOhmF
Z9n7WR9/NAmOiCKJXKmhwuF82i49d+Af4d/9sYG1BjVExPMWOgc3aRBh9xcZ7iDiNOow9GtfwGWS
BlItCO7Bf/r/kZ+iyJ95qngRCL8rRWtKlD8e/VEupkBnpilB4f0pKE56V6Qu0QttVEvw0ciKXAJf
wpx9RmS/kMpcKshMoW1gwnyvOxk1I779Oy13PQ9lVPeiP6OAxkDVxoktv4dCkaZMB6oxzYeAU9/h
5v42NgJmnggbQuhoZGZX62wFji8NvFBBClaIuLyeHzWYajKzHLei+dXc7Q3Uj/D9e9WkpSC7UDcm
iRokzZFRosgOCUTcC66vwQCxvP6S5cWFsg7ohiOA2BRCA9UtMGHcTx7e43IuWDJiujf6hVH/GNQz
rOts1R9n8Z0UHiUhFQaA0uAUX6SEHTHUKxwEvmwlFk5g5Zi7N+7iyP68A3WpLNyuSZDocCspkydh
HaFVZAkbs2aZ7QvxRS8ycCJSRK98WXQeDyeneswdp6m//xmtcuk+FIBHvR+qITY+Gvl+irt66U67
04SPvyk3R96iFxPyCi3gE4I68pz+1ppJfJz/O85ARp0QrkaZwCmd2z2jKEPxdlHs8umq85jINDHL
GD2utaiCvA2oVw89C2Erhg6F/DBA8yN8dyqIidPBFsAtEeta0gIzbK8USMLuj4LMuVkn9yNQ6Ba1
hy9GR8zPQtbkDZK5QLss/O/TDuZLoP/DjMejhi089EJpw2AyEPdNPItHQ1VkxkUVMT9olOUbp6/V
+4UBOKIrjUQH0NIZGV9lXzVwIQhlZMzG7LHJDjUJf+kBIeZ4fb+/XAAAL7T7gDrKa0Dq5BfQlDdN
oYIbDupWOrNAokdNRm+e72Erf1C6RzpElHCLzCF7s7kogh7IaR11LEcneXW2eA0RTTW2/aUS6LCq
Bd6VxowSMjkYnI2Uyjy/fA9ljrhgzTp7OPBvgOAzPRvvIf/wrQN+y2pkrCmSO6gJF5qfGKvLgXyU
fMOxyC18yJi/cXNPT/2AWX2k7mhNcqz94D6Mk3+IrORTlUniF3X99fXxiiBcTFu5CGi8xV5BywHb
MucJkm0gCbaWjArOiRe1ZmpbEePP1xgJa/CSGh7hsqgObaxaY7k7kuF5OiTTPbXAJgGBw7/DkEzE
XW5GQ/c73u2r9SWcPc9OZIzjL9H5+iLyftPC43Xg7EiCKZ+Uc5/u5gqR/0pMGzXdWeyjgEmJD/HR
xmKNQomWBRRHLy72k3fZy/68Ro6I+QB12/ZADM6eRmg0OHioBvqNm3Vo1nz76eHSXpaHcFzKiBnv
CT3fs7JmjJI188oRn/rhwwKQeDUnDE+29kux7k3pTRpiMNxTeteUhC/S20c6aNzPm1ekNwOwwTXZ
Fj6/znlqRlQyl4wBLPYqKwU2YCHm6Zq3s1ftE9Jv4sAJD39P1+nFTxUK223+T28oHlybn3tMAOD/
V0ECLm7B68Gk56iq/wGApWvL4a5H5/LTX0/G3tE1Xc/Ngo4PtVoIEMXGqfTcrAGcedTPsZweQRe9
SgYa1kIth36Wr7YxkrhQD8iWkjv16yzUrFwTV9OByQTYE+/oyGK0TPvTetiqHV8Alt8Q9INQBE6C
hX1yJcVKbSyUvGkVSJM0JoAcfebDQTukD1DTDkFY1RqFdKMu210reYzQ2IzhhtB3pe9LoI9QFQUP
X7uMTKlb5tpqrIIPrKhJyBZH38fBUs8+v8ehwV5jIXIQGhrs9V/hPLayZyJ29iQ1O8o/zDJk8gvT
9KsjQlEbwCfufqcayNjnymcQbhrmulRtTgVwkSwd/sD6u1Wd8kG/5fc6PbR6/jfw7DHl2lFpHOBb
tjaK1GGhUdyvltKaJHgJWkKl9ghV+5K2aJ4WYUbLieMdpwPY7LIJxcQepJXabrhqskYDtd7suiK1
NDzoygpvx/urfCzsTtAJI1/ar0miXyN8nVDfcIkyO3rVbsx48UC8UvW4f+VCMvuawI7uIYHLbTXC
3s86oNwDWT6Ym8yo7qDjBrmFf9k1U5XPh8I5T+DBUe2rm03Dc4wobZz0omF7fspdxggO7p6GAfXL
H9fTHRtjZveyLPbO6aJNz+ZnGuZyswwO9UmO9o5YVv70KJrmjHnKBxawyu8C/VY7gh6hmnhRg0KQ
NyUpDHsm2GF8HvHqiw8FOQ4N3LOJ1XH727I8r6rnmuQKKEhP+o6tg7sDA+JC5RDuLYDh6N9cpHRH
iqjJVnwQsylHhpDvDZ4Qq78QGPZA/MQuTN+JayDq91ozNyvDARwJIf6voMqKIWHhqsEttRFd8Iew
r1MpUestfsvt0XCvVJLqB0S+PXLpOzkHI/ayEaW2DL0RebzkEGcSHUGdKh8IsIbTsmrXdbDmvUJa
HAG10+KfIVvYtlBYbR2QSa14hyJ1DNAqtQrGy3vi+XZpF+yQVfIvbjLDOJs60P82ljvsIdAoOKfj
M0eJpOYWKyWR9fNGajG/7767ftYmlMMii2wINtcoPmIoWKMBSsxyjnxhJP4MbIe4ImIgsA7CvQHN
xv5gGQgEJkELh0F0LwxM+APciykB+OG3dFX/lSb93mLvVfQuJzo8t4kXjblgq5iUdqP+iBTTNaaE
Tis0/OrhCewuC4DPVtdjYRuV0ks/Qf4PAD4g8j4fYVPyrC+sTJXuaqunBmsF2nDyILPorBallr1i
O6Dizm6FaKSADWkaEnL4sR9s+qlmN0LbdPFdxVNPnhdix9tH2SnAfUNJYphd1BE36gINr4cbgCnY
oh4QHLE93B5O+HX14jMig5oyxfLoNn4Y8bSb73+P006GsM5f8eNPT2iC6Ox3aBZ2As2F2v+fdCRT
XV5rR9h1HDAvO6FdMmJq4UKT6vbk0GtYQcqlGCVzY4rbWhiKPkfByhEKN048lOJdrSPL6Fzd6jix
GIrWDW/zhDpw1deUslwHHicU6WiCxTc4c3mmN5YXz9G3Jd019Ynrnqd9uaYra/RlgvpH4KopssY6
h5Yux/ZjKDtZCaEntXEbfAsNW13cgfscXkwD2q+EIYrDmELevsyCS5C4m9rxdGc0pqoZcNKQjXys
gjy2A5kLsvH1wzXqY8bb9MdRPmHdkMu5/y7TpC+kRiwoZl+DeWVW9ImdBR/EG3I0d6ETbONK18WJ
TuCKyKUVBE7fRXOefyYebWBsTDDWWLRiXb0UWtkS1gZh1mp45+BR/d6sbWRi9NSjiV56zQudYvgo
7+BPdapE2ESAjPoohDt62lybWTlc9Me+6YZIqeveqD4RVIQQIrYZtK7h1hh/jV2Hh2u1BX8Yu6mU
Q2nULh+rhTB6fE4AviU5PJHSAaiHR3SiCUjGQ7Vb5QIAGvVvx6J6lxwdWFoaYaxXlTZ70CABExDe
v4dCu5lVeug1U1COqyc2O2LA8jrI+G1hbbqHmYt+FatP4x/G0R011ydGz/a0DELXwJfcpuF8w66Z
37CbdKAJGnQPxPa7qLk9jVjO5BEFJ5d6KvJOfRQzgvkmBMZbHf0UUrIYNZP12Cu7LGE220+u5fsN
Kc7t3aUwu+6d+HDr+HzKjQhOKBWKtPAdVjUjMCBlXzVL08y+bKjWq/SSWo1QTWYb7ksWH6laE3Jw
mxpjZKq1eo5eVCu14pYSp7QqSIjiFk8WBZi4LwfyGn6uo21C+GGHG3o6tZCi9WQjckAXti002hTC
ZuEvSfXjwW3QRwqJig0AHa8wLfThoQTiIcs9KgrEtiDR8gI1/pU7khv6btpyquMgW3r9fPIMvStS
tGC3Fm4apFLPXcX58fEiRnwYMgZYswu3ebAUgfqm+mbxvcTHeFJOoWlCMUramb9X+2v6p41KGmKw
Aj2LPN53bO6OqF6h1BlHkM5hKki6z2hEwLJgy6L/ZO/4z2cxOvLIiAVxNIiKQUmu2leJL+GMCRNr
v0MjnvKZiAoioAsdotEEEdQp+rlG15q7UYgjWRPKTsFy4mvm8Zk7ANDCyqVfHmDFguIiWWLzSGd4
erdeByFq9TERA7NwXRoUxXvUqCxIicriZufFBThEr+gnOh3QQLmkbBgtqc54HIGzT/LJ2cJwU4xW
CGkRvz/9uiGam5gAwJU5XWa26+slDFnbjzTp9Nehzc8kCq5fQs1It3g39I30S+bgttDQ8P2q19zI
B9oE5DCuGRutvPBkRgeqs9YEEoS9csPiiS5RHXCalKydEg61CaXHvkhDQxcuHYqvpQ++gwerDJtJ
/C3GjDfoarT4lYm0GvCXgj3bnO01Kp7cgmL1ijCA5qxBHQqRp9m191j1pIyexor1aLVcKzTD5JT6
/qFLjbuw+CwcMQr9ddcboUn4IRYn446f0jO5YZKjr7REOZXP/CBjJVpDYTL8GhQhlN5PDiTTr4aY
IHTIvmlyDdaDrTkh9J3fvrDXAfKTLaFnqPRyZbTyR12aEJV87ge+ow/Y5GSRpzve9AYqX3UhJTYF
5PGu1BdD6BfdpZDqzQLpHoR2SHlKJEgZiDEIw9RkKAgotfpKnRG2ZYXbcMcqJKoVFVItNIE/rDfw
ID7qCPr+M2tsP/sw7XKLF3inJ3kc1O0f1FawSkaMNcy1/kwccpMhEZ1GVQYPeEoT7Dhsj8K11+Jl
Bo+rLBM+L1KjpWV+n6CvR2R0tbgh+iyLF5ehdC5SBb4rAawjfuGFEaptrIwlKF6B0LbdZn+u8P/9
UAONn2FpYtbFeBozMNb22Ko0q8Otjjfj+ZZwC2Q0qrW9YCrFVek/pBACSE3wz1feqpA11PW7hDAv
ybqCKEOgHWTOtOMaELJRA2hrkDxR8MZbXvhOjA/TOxU4VCSxmOrwtMXF1gvPiJAqZoR4AxlKE5o2
FOwSWuGIA6aIEvOFi6eFY2/4/Vlr+VVG3y+OnAwrmXlmFe75y/NgUA5QHQgI0EWqPqT6k4q7AEcf
pRWuT+PVKfT+dejk4q0PMqBifyWXzgyUj9U2m7rOJSwNhYSU+6klw1+uPaV2DJ1IbhMwXLrWDR8/
x10pn5ubKsuQ740EjPy8V+gE1b7T9W/9ThJJMWw+BcG5L+zikZu1JMYbn5ZoJkcbdLbizaPYJUuA
aRoMKuHck1qSvZw9L7QrNl4BWblBHQnic/b/QJiwACuLwIFlcRZAT8ZyPuwKXQfwS6QS/tJMuTJZ
SM8EOelysTZEgHKAdcnH1sh4dyyKcLNMH+YmX0zbzocavR47p1gs6YTLeUMfiMCdmwyMazo8GHJ+
Io5sE7/9VRD5cct2YcT/rLHDMiPKT2FbygIFJDd86sAwtCW2mD/yIuqevpeD8rNXuqkmQGw5iZtI
2lZdnIzR0fcE+U1nBMge9tYnIsm2RK88BtA635QFP4+QiozKsj2Q+gA6bITsppg4XR3zNn/ypXbD
iMq2Yv0h2ZGVHQbux3pFUFjJHbngrNgR7ZmnFYGoMM0tO76T7nlEK3QMb1It/+6a5S05jkqmNNpp
ddWfeDDkCIFqCnYnVgjcePKwjJVAnwEHOdXcri0UbnJvhP2vHJJFLekr7MDBHF+AasiZNUjm2L5W
NzgWsykePcX2fNfe3irrOgwizM+b54KKo1M4ndxB+G6cYehFIJuR+luwmt7qimnxE1mcYbL19hvZ
dcIwzz/AdMYVDzxELszi+IkTxgzvvxmiwubXRRlH22vREeXwn9z1buYnCtQT0oOZJiRkefXif1Pk
WEom3OWj/HC3NaKX2cSHY3vETTGGMzMQ6M07SlejMcV9vpH+7ko4ks8V9LfLoZVbc2XodMm0anoD
wE+REEtNHtxwKnRHF1izvEKKk3IdLAQpfpyd5Sc8HNj94tJaeh2VVfYmbsAIssTDN9thFV/roSjB
8Xy28y9zat1hu2nlalam0xG2cSMq6jchO3N9Wp6fETAgddlAQaR/2vUSuSAogzhv2alzjlMO8Jda
ZrVUESIGRfFv4p8XbpVCuxm5JNlCUrPsXm4ELa3eDs2pMbtRqkFf5acGSBz1WAo3QcQG9t7g9bjx
8xDY36ILNlgOHycWHcfjT03lTCEtym/YQ7SGBkCFRHDKgLDtbmRriQP+Yc23ongV/dtKJANtcEb0
hWquoBCPm+8ZaB1aKm2iZK9ACqkfhqliq87ZbD1cxAEllVId22/Ej5eMEFzkmvqm6wWx33axZNVJ
/CZuFMUuxuvJJCPEgC0d4oYtYpDpJceaXBOov/hCO8VaVsGjCfa7ENW0aiqePfouRmvtao1iy70R
Z/aNbdT7JgpVlL7+U50+ObEh/duLyLS4Lp6Z7+H9YANB70Zx0ZM8rr819DF8lIiZixi9rXcCtCfK
cBDschYjqUTVgAJxflpuNaN0Tc+o4iAHxldCVWpwOuAIuB8ECQZDp/eIHmqSAF9wFTnVKH97ndw2
vxwQflybUlLCoQkb1ZfH/IUDpeqNch+FkkoJqbictioDTn9NDEKQ1xxyZkZxa+qYECbh0KAUHhcL
si9L0wxXe+PyqsNAIlAkbo254EMtC+/aXhvL7mae7ee0onJRElKYEP2zdE2CDCZE9eL6HgWRZVmr
eKu8Kv++BveKZgjwh0VmFitb86Y/5ViWHLwitlKLXGXxCjOvoti1uxAFPGGwRVBeODdW0PJAu1+A
m9tuNOvzJ15U6PHFZ3DrKRx0dqecPxgM7rFeofOR1aYvCZYyXX5Ziw4KeZ5vWSmuVO9tk3yJusb1
/WqThcDARdWhf58Ez2b3ivxx0o7JJkBZ20dpAoS5oraMyyIWnHWeXPkpnK201RIgkQBCltpUL0fo
/XZdYFP2tKOdmu0mHBTRz4YqKORJtTkevjv9uMMa1TYdoUFSRfwO6N//7xJWH9lztKio3FX5DMKU
/ofxsd0g3H1cLDCBdM1N+YzoohDldAgkLDSSWRnEsZOAILyZS1vZqN4tR/Pv6JIhWGphGDXyfJRT
AvL8cmPNU5YrQxergsVywAFLsTgM0aHYngTsoIYuGM1OcErSzuePPOWdFfy5Jt3bCqNMrXXitu7D
4V35lQZu1ES53KxDtw022IowLJtpOMd2JU03gqXINck7QrcBUASauxYLC041M3W10knVHgXBWDni
auX2YhUfBWAdQ2Fdtb4KOBVnjQ42hOvGB5Y0R7PqHhrSTgDASsp/zsVoHaxgrw4Jwdt8u7klr7Rw
H8JAQnStSY4rUjVmwQy9/jdBk/ZTZRy/Cz478adUvmeQXuUXELDSceK2gdaftUXZLwNnNfM1qpDt
kqPwuByjkiiMEnwFifS3HW35mZyArFdeLGG/7OWm11aXzMu8o0t3cZL1/R7YB7XFsuGxkRi+lf00
QhlGElLLneLRLjuffW+nXog0ByGgj8jilbHbkH+WyJoZcCB1CLYhCBLvonwh6E3lXlz4913grVHP
LNuXN7S4liTxWgoccF+AmvgmdGPndvxL6W61g3an91hOF8qyEANVHd7be31XST3d4dCLbZIQIzw+
yph44xmXAQawDjs/z/BBX+ylHNqp0Ya8dIM/vtzvKENytYS6wvKb2GmV/n0bNH6wZHJ4fsmn/6Z+
1SLJbZdnni2reZH8jDmR0BgP3nfZRPMqSnmkOTXYhz5L4QmmLQCI5n8hs8areCz9NCbrB3ZCtES3
K+OEnkcCmqVyZ55fuGXH8hl1kwSJue7F8LGeqt9/8dhIC5F+jaf0EbyO0KUIBaUu38zhGdh41Tjw
Jka+FDGnp2jCqDF8q0KMCf23Cp2pCh4fmhdJwpeZP5mB3j1OT4GzLuQfcwTDshL1lsn6mnzjfQQF
VlR10bDX1EwM+QcZc81tvpPdcCRb98w4TDatCEUW8GwLB1Y2jt2cHbLysKF54bvmHIjnFTjh4t7y
/GItXd2FUPBBTYVpxVE7qrTW8eeqB9NYIQdkP4fc2ZuJs+1+PmAlf9KNnJMnqh+VRFxWFqdQBJPM
aLq9Uz8r6KBpksDSh42aw1cHMesvrYTl00dkbgBq7i+emyutgvVWJmObZdBxq8O7P+4M/6I2i76B
4scZvoq2eTX8keonT18UOi22HJTSaocVTFWnJDDlDTBGGNbwONNDwEdFnb+Q2VTwEn8vEv+nu8an
P1KaFrZ/iUolCxyoUal1e/7349vTW7R9ftYvLD+PgCKIVRrQ95RptaYU2jJvphoWeMJgPeT10QDm
vza/F2KORbdX1rpnm4Tecks7EHBGY4xv5kGa/ggdA3V7MDLSCUbE4Lqsnd+uW8hkEd47jtIcNcUN
p3PpnTAaxUYesBT7PiUBHcDo5P5P2qmu2rSuCR2AuVfXUsVQHxX9a4C7BsLxbyn5EdRr2RyOwtFP
eq9H5LU9Ysnn0eVyypVBEfJXLacCwMnMNVdo7QhfIbVqh+kXo4WagwGYOfB8SY5EMbsANXhUCj5S
zRwCTe4KuU9vdo855M5WsXKJvbGEaW9KoVAgNXhnCT+4lFffRoszXxGMMVFUSe9n6vwlqtpkjZ9t
/pe9Onidik2REUyKch19Poq0NKvRNviiIPXaUDxAOlHqvRBL3dHZRfUQfNRWIxsZxbuuhYWypVKz
y1O1J2+05n/S/Ih/vyKFv3XZ1RlRqFP1SsM/4FH4Mwq42Gj+8xIjjKB+uAu0OwX8CU2w+vaITPYG
/7dKwp7k1jK9eZ9vk75iYCAGME2ICv0t57q/akd6vlVTrRj/ecvtuOfNfhJcSbaIIewQhi+uc2Np
74i9JKdkPA6nskQ/ShQ3uMYZCJOqOrD4Xj9OEEQhlTb9+g71z1Iz26LIEON7+98n5jIO2S0tLQPq
Ut+jI7Q2hc5HsUDs/ZBg/5RjwvDsen+xE6ksxfmnqDYoF5iQ7vSUXZoeexlEZiRK12pZMdBhxoHh
va2P0Smp6qfhRJlFewhBJsz6XQqlyi6T3ZkCuQ1Hq16WvsqzeBU2tbJDTAIINSGwL3qtNOQ2yXMJ
g/CgyLVi0XTiZKla68n22YWrfpY5/ARsFXljeSi8ocQNAP0UcAK6GVFL6iQnT/swY98CZYnsVkmW
1sqw8PxawUeaVFG56utCOIwf7/PQsc5WVLHplRQb+GEP+IwIBHJdqUoI4/nvpGTH6M6tWWCm7Wna
hILpITswGCB2u9DpwKa3pTWxuK2nEBy4/V5WOWURcLFH77WmI04aw9KLScbhvt2F05U/CwBJmV0Z
/nGHv97SrJ1vT6l5pDoHT7M3qUfBJVSPG6pSXiID2C7lrYDJYbi5wp2B329jkxOy7b4HRYmHo+9Q
84v+gw7FRZlX4RdrDsT9REfZSNV62wpTX4kqDqVHcxQh+P8Htd5vMHxCmYpobVPPtDVFwdp8I0GL
Ol3qvd/zSEOe5+ZpTUkxhjeTOiQxArU1bNbZNJ7IBvp102do9HrTPOQUk6b2/9+57qbUqp8fBA2u
E3McmOGS1jwTrBPHUP891yueNN+YgKfiphK8lcM3UJWgw6Cec1B1VXMJCIrJJtWpDQ5KgpLZ7ope
Exzc4GHcGkUbOKzKqnO+0GuD6CaEIpqPlCNCDpglXgIBgslHCMsxc19pRuy/AtSpbLNU4xDTxrbK
5CswHF8FoF+elJS9fpBtVpM1MflNi4fzwrs6vf4HvyS1uVw+A66uXPd+y2n65AHERXZSa3dPykTp
boAT9m958KhlHwtU8oOsX7g44f0eBriIQvYEGjQ87wtnkcKa7zHy83GA+/E1Ua9jMIq5OBRVm6TZ
uoGTaRpQ5+gkgEN4t+ILG1Q0n7OUrDMGjhPV7JKv/ZTKgN8aiyiQhAdHDxufcIDuVVIlj3XfEF27
4be0EOpgHX2PR182K1VD4R+zQVyQWlIXxbwc5JWC648xapc6tibLmiDWwUP3q0brwmWamdAdOBzo
AD30Z/1L2rGWI8HV8UgLHJokIeS3Okri/JNXlRX3O16Iq1Zvb4km/WXIvuX4p/hNwB9KsSjFJbON
jjyuGMVtcRzInIbTMbKnYjKakLZealIMTijy04ZB3aymTYNQhALyZoLYtSZfNK5YCDi1Etr8IuXU
IqHR2AYlQfzAHSk6et/qpW6r7js+YJBXlZkTQV8UTHObbTmqOu9bzOC11Hs3YFDij3j/cDnhZL+X
7N9IL0Zrh3+FooiGcS+EPJ0w3SVipQ1Sa/AgQPT3tpKAzTDIImi6JZGgVNScqNCIKAJvzv9nhw6H
KIYvkCi/lWAy51WPtoPQJyUuPUz+yowptYC0HKGipI98i4yW4mhOU2ZQfJ6HcZ4oHNq4CSuiPZ6R
It4fm9kpYXQRwXksXa6kRJY74nDi9fXEGlbmIQAZAt15P5Oit7dFYIaB3dINbAMpSn6hDOAjpUhu
r1I5fIKsAoNYnzDo6/sc49vYD5m4uUHfgJWQ9ZiNAwqXip2iPpWYLapAiKOn+nSHHNzYxp9DK6wA
n2inVRzU3zimGj3ARa8TqZ8LL7b2A8LTRk31Ay5ufWsq7WTHpR1DNFgatjp8V+8E1H2ODn0eLOgw
v+N+GYrFwTPWNgS/Ne4xbAcHW3iZqslqS7HJfqJsUEigAIXqxI0l8Ng2MhQlB/sKR0wuwO5S6IJY
n5H16Victd8kWBiXFZmHLHmMKxsnoKo6+2cILiYbRJCEQqDo8vsIAMNaipi5QG8Pqehjg+wewzgk
VvyEYfPj4YOdGvjYcErA9EMjV730lcAZ+nc7hIa/996OcChaJM/gkWmRjwK7dtvosajS0FCUySif
rw4Qh25K9KJIRIV5lB67U+HaeyYP7fLGnNPAZHGDXVpIOFBbMFOVKxPJl2kh3C7KODB5e4NFdxru
QWnZGPQaO5VoaH2Drvsk6Psvp0rxl4VJ//lt3vfOZFHcJojTUPqyOIGfiQo16Kcf4T5YljQPNB/5
rkgRqhcggCNQ24szsOAzD4rzvXdXJj6GJEjyGZ/NHqSCyi/RMBXPdlaXUm75bi/b/HhuQSzRD0bw
OD4Bn7XeQlhwDbEF251kJIpnzkpPMDmMQvY9I9B707OeoboU/eWpsuj88bAR41D+fhB2Kh09EPOl
s7vCkpf2b8AslS4/Kptd8PSMCXqzFbJ7FsYh5rMrKO+gVO+ItwM0y5cuIZo4poQvttGJqk7YvSgJ
L4kppHGS/gaeozsZWcmR+NEk17OEBaqmUAxR3k3AQUb9jzQugcZPZp6KGePhh8PRoS8tUdkKMP81
BirpS+TD/43++rBDeiBO5lOl+Ihmeugs+zM4PeXbiGQBfAmclmpwp8ZYk9mEu3IGaITbvAyTBfLK
HJz+GGG7BEmoAvnIlNbGpP+JBMj5Wz7amg4RGXPR7sEfW4NXhSfHbRwsxwOjUC2jl0Zx39qBdUmp
WlpvYEIZrlR+UjYQ1lh9JED2QbnEEGV+MbsRg2anjdqlCfKMZRRkP4K+z2poImbYzDmdcnW7mOzB
6bHGxitZwh2wMz7HX2hbdju8UG4VyP73d9IYjSN5pVCgjuHbTXrNYdOuHZs14o125T1vRbXG/xOt
LJwkJoSRjcQh0Y9rP9z6agm8JlXzwIhElcGcz6iYPdIthyB4U0K5xqVbeIiMQhKuEV8m2gFbIt4s
gwUZvopHXZjs7ySoFuu8slgIFAEbCNOlCjNVEqgnKX+EvFjGXLv1XrkHja8/lVDcvV02UvzN4Wgo
wBOPJ3fIPFBg8lG+l/3AQwbcatpXd2rgndio9SwDejrky3nfJCC3cOZvzXDQhGm42CHzdm2HEMdM
k6QkzjxTy0FdJwx7lTtnLF9EiDKyQ0aItw5+LBrA4sP3r6gciemYUui1475CoeCxI5TbEZus7jtb
bpK/5b2ULoX2VG7sHFmJzzGQJs0EQeX3KbqYQpmoDxcKDL7VzLJIhidvZrNjK9kKhDBNS/ZoBE6l
Wpv3RKKECY1I0sZ8J5A4UbMCcUBxfMKh2ggPPLrhgXz5rkMNYFJsW6dATvAEKviEe6m/OlFH6PHC
r5Hk5Aon8SMqJ0qFZ4/2aLLuEZ2ewQUtK2zz3B/gf488HWh9viRpHaFvaXHATeKfFikdokQ28q9f
wE/gOoHlPVd9c/UTl3lWMb63+7hgra5VNvwyV/Ma29ZdiRIRcZ/sPfz2GUZBYLJNmlRsHDyKNCvm
vm3m6Javr00hsCaaJGoYpAiow2heKnnXrU05LiOH4krRcAUoRwt0GeiEwVN/A31IJ2bxhEh9jovy
jIi1C5Wji5sTaSLjkGwx4c8ExboOvdI8EJ+zRv9w/PDihWUlR4LztWbI8FHOq/HwOaFlzuI0iHbU
HV2uqhASd7P26UshnU1WE2nIcytJJ1Ditoqy5kXbsyphQDYIoDTTLM2N1zXAG19PSHf8EzIVSt+L
HGkl7P+GeGPWbTFyjGIHbQEnKSa1YsuiilH0uVZbaHKNyJ0RinklVK4CX5JW9xgMA2ciCy20XJ/o
EcoEbIdc2Hlhm8N6b1lTvCSQA++x0DLOF7QBP9TbcIFazVPSXrLbKYTG5WKP5xeU0t/56GgwX++Y
Hr6VJPU7efGBthkqhzkFzXleOK2h/MjAY7+oZCAF+6Y/q/ZfN4+Xy0FITjzSnW9pUls86x0Aw5A0
pDYUy5zLtmPdyEgC7Zty9J2fZ80CQUFda46b7gB8i1dnbWP2rD8Y7T0fzD7U7iicwct7tvtc8b/k
AVj1YPTS6X0SEoL3E+ndswgFx6eknFDnI0hfIrEvPfrA5xlNmkyMT0bAEFKaWm8AciamsT5zwZCE
3MUdBU2GQqudNg+qPxXHkG30C658BjP5dIjnfWPEOhH7RdkSzlP3ugtYiWKm4ORL/9IWlE33/3aI
DsNjklzfecNbSl4KCi1t5CXIlOLB9Hhr+Z5YFqkIeigKAS+kNZf4UG9P5p2p4Sg5EJ2STxR+PDx8
dpWPjsE8YnSzX++q9iXNnWkEweRDJUk+ztMCe7tO/av/xiOwpndvU1Ob461a312uqK2TD6z7XN0P
v8WYJtumB0mzu/yfyjr7D1fOCMNRl2fnvGDuCC107XpFKALRU4SjRXZF1UDeUyMLxdi6j04QVnrX
WNtqXybLTlVJ5TjXjG3NNNMQWIus3mkrmiCq1KrJQTjv4k04wXHO0Whvuttm7Q9yTXNlm3nfUpKj
NBZQkSvgHEWxVT59IQ4GbMXWGP7fqG25E4V9Re7dbtDwpp8AkeKO8jZZMSjVQFVqGTOxGnSdiDB2
EYElxzUpa5udYZ9JTWMrBYCALfcoUh5sBAQ5b4x5V1NIjjJgdKO7fOSUNJAhDDR563hamYfsrTFt
BM2IzeBX7zJF2xuiWwpb5X25lHCxfobBwlIKUsyU+D06Azwa+468Le6AusWWPSlxKxdRsNOjndZc
GdVq48dsbKY9zT6EnkTVukfCsgWCFgTUo5qVTbSbWfwMTJKJ9LeHOaZiH5Ps6XeUtK5pLprAGr0f
0Kv/Z0T1dVrL77cGebOl94DQKkDl8GZoS6VM6vPmG76wLbsL1E3le39VTWjtJeBSSD8L3Y4iPfxV
SDQIPJUKGhEWB+AsKrFg60h4f5YbAkZ7neSKzmY+4Q76YMCxPchQlOD+QwIahUcm4/fmjSmZh4PR
KTRZw55+8xWjqTUip5o0G4wnHevFGLMXnvO4mVYMME7ZbJBoTBiagC8YIFFtWzIxj0QgOArJvzOQ
YQnZWwLQyfMNqVr+wX2L+z6dnvvdPQXpa42PIpCvKvhFGTa06CAU1bWSaSW0fn48AQNYCM8cEmi8
acxvtja93vzz1YPm1qQYzW7BPrFRvhdesWW0PpOgM8YmiENc5wVtfVFn2GTeD9eHUaFBw/PfBouO
4fDnoNsUy5Jkh6Gh9p+naziPEEE1NqZMLXc7vmWI/Hn5cvXdbAcvnnT4dwNM25TSR+Dd7sslxmBl
3Y6czB4s8uNBSvJswfNVU45QPUGvdll7czPk/LCtJssKunE/qfem/oxmPt5WDVKgEANuYSEmMcaZ
mp1gEdHv8kURZD+Q3kaxAVOifDNEOWR4CnAMBUVRQq/7lPuhsU3gxnKYuEjUnDbnkz8TEYQVne0y
AyNB0d2wxJvVoaoFlwxOFgWLUXQuYAjL9Z6Xas3NDN1mIY8CVfCUTIw94LiVvFAINYsDTY6im4NK
XIo2bkSz8WODKDuqJKhDLqkCSxWiqZMOuQJ500X1OST18PeO6xJAd3FS9NHasetB0uzGr0yDPaWn
QxWQC2fUZ9rmwzkuPSSUAs847/zCqnm0k6zkMDlHNB8GBl3+9UKicvkMyYvKVXJGvWX0zECV68ws
wLNY6wRusonfl2rPQsztLL97LvnJjikRecSxY/5PCkUDO+vXr9nYXh494H6ltoCttalDMS8s5qLr
TnuNQnxaPlcBDoLAbyWnIrMVCm4QtxhWZAGY6BgmRpl3lf5QITKkwEFNeYRdblcKVMHCNIYTLWU+
Ga3L2zO5sUHXEUBu6UCeiBhm1FViHZUdjV7ZnTlBF/iXlm8E3riu7EV1+YB/UYia8/j/jwoiYOPF
bHmJq4JC4vO1vm4Hswf/7Ju+H9SyxIwd5dPAf+dDP7YD+/AHks2bwABlh3BRQwvZdwmlWFoJfFOd
MbybN+iWxs4HaJbBGB4FX184yzMja/0ebnypxhq16Bl0AViflJWpAgMpEVyxcsFJZvBxI19zgDpu
GMNs4iVQusd1rhFzWyg7/02nY7XMsLaxKC+fJ4Q3B3XjJ15moq24QisfOoyc5zbTPZxqWf2quaqr
NFV1wFhFanT4jtr5gdsA6XibggC0P/xgg4LmHE9rnF45OCj0xD1v22eEqaM0vVAOiaeovOS6ZhRU
PhMFvA5TtttqkycnocQu9Ucn2c7FU6r5RTiQFtLhICOJqOQNa42gSe0ANlXKWQ5OlP5/vknM4JTM
qUjPskFObEM+EY1TZh1wZ9D9X4v6bVYBOamhaUcSX8FbGGP7DUxnH4xF9jzdLcXjiVI/oQt/QWyG
r6WN0tVEtlsYxEZKv0We4C1m2BDrMQRzPifh5K9KuIuc9uMq8B0ME2JRQBcUdN+LN6xyzXZTxWKS
M22trrQ8rbCbEeZ4NCeIymylz6gqD/c4aU1y/R2wtQdu+wIN541sUyahSpLl2DAljeRj1uMXua2T
fbwAWI6oT0nZC4gaZegoespbMVX81nwbMkB5NGeUVwYZrnJSosnTt4aKQp8uQIgLNmPBCxAsqFhX
5LnO+GEnryfMvGuoeM9cAYquhXGaQ9pkMz6Mmr27hrzKVFb2zCfpVxu+o+HiMr8FsWAeDkms7im+
DPfiaLG98FBqRMe6Jx5muEn9E+SRUiAwl21MWFLciJcotB9vExFcL4C+tW2kIG5w6uDSQxiFv++b
LhQPoF0Dt8iqPkuso/j3sXrtTWXO6DCUGdNvn9XeteE8jBT6V+BZzKBTj1CxNb+0O5j6FfDJroHI
y46tDaU5woqqa3V/x9LzrNjvA3vfYettp+oyb7MRMpYz67aEaK+8FoECbL2RJ11PrHlKfNxKspvD
H8oMBGyOu3fhIUsCl+ph9cADouGcFIerBAscTFKD84i2Gv3yhFPvSbabMWxtfWUN/faYkZAIp2pH
n4kzFifFfkscYz0yte19oa05bcnzKQDSYJMy3XYEYceFmmcFo2Qc08Gdbqpo9D8AhB3My2STT6UO
Y/KwbyuKfC8x/BrQ6UHeB0R04nqXQ/i5Pd9b2DWbBMKZk0uhCklyP3bsb4BZ/RdltCSLdace/kEv
iz9lLAGxlQkriKF8j18DB0FA7a2JvtJWJdnjVckhiZmw/DyJUo4amEcKX3Ltn812Df91y49nJSPx
uKZJb/s9CYRAVzB2tD9iwo327b2j36P7vb7GO5M1GGu8b7m+fKdLU6LPOGIXezveV/yhWfyFLrou
iR57Ea0zdAtiklEf44huR3q014/2L5H+yEwSFdy+IQ4mwy5VLx9cUwFV0Syh4ejRLKdt295KllHZ
Q0jNknu4T7wi3r2DYecprkWRMYQh49exW71DpOpcG05rdZSqsJdXXPVc31QDpAV7uYO6+IAs8dLM
vW0os/nbaSvvQZY8KnP9Vli/73viu8FPgTryZuBUs5YERkPMI3gPTerze6ijtN3S8TKT90gM7Y26
wQwA8p8HyKkd4AH3mA6AVqxgcfOdvXLAJaLJfWoKDYphcGwmYPAy6BCvn1M4ly0bIMDra8moleXG
HAhVCdYbYadbBoXKPcDY1bnY/5Qd2OwPTX29iVmfyU5RaSmMjI6VOpVL/uOoDEbIDiDk5ViZ8bU1
dNd79/0431QxhiOrnwYg0q/v9Exp6NJ7iKWr/ki2YykzBk7p1h5wHLkYpf5AajF8yTmGT0UEAJpB
0JjyOrnr5VnlZKX1YMlLA38+o48ZOvPk+ExmSRZLnhGUNAjNbGBLrGHObDNld8YqeFlhM2MJXhAO
VovfeU3V1/GL09r+h4l+1dCzSo7IVzALkMzLIJNHq4aFZ9L6FaaAiKX4s1pChta4e/hxqtITmchC
W3LIsXwYrNwze53TR5gC8Or8xFDLvP2cjpHHV/oH0Vm1yln7dL7TChiOMA1/ABnZmogyrej6Hp9w
7kAGVDR7w++Sx6mFkDdpB7CzZfKdeXCKU6m4N8aVowA5CAuRYibpx7rqbLUHzrGeBb+PX+PAHSdD
bkbgphsfqCxjSho/es7G5+GuKRKj5GGVnUg0Gepj5rMGkg8aUFjVDXp9mXhnJNcoCQQHsznptVrc
6aQ6+GPfkrJgwreT5f/3MbSANxI6rLIZQ0DlmyZpbvzx1fI2jFoEqCMGiWwR02r7d1LQ38acXIAJ
xPa7Itlik2BGou1A6f2Q2CwrALY2rO/HLSrA4FSoPUv0Tw3m86vTNZwxrZNnNvvykmrPLMcir81N
TPndNj0w/Oyt3OItipiPQUtz4Wyepp13sD6ozOT9c0I6a9c9ydARCk8fA6Uoh5JB7i6R74B9dt9a
/tZ+S80XWQjQ4ZGphA11nbVTcSJBxiSNe99M20s/YLS53q0KF0oHupHwDmaqORpRsJ6BxdeBZuf4
9VZqc/PQQ9rECzVFYgRzrH6E6fMoMBmMWKanclBoD+H5RgAbh1H5NGBF17Mo8APWD8j8oUOYkpT3
hmX1ykst+idXSf4Qt8R+tcOYB8hPyvVwLilhpY6Rd9aNT+CSp8KgGldoScEMpzOpDpy6/UgR+ALG
pZ6OWanGXM7V7UtpEQRVAEpHIk644BsubWR2a5cQgZpfq/Cfs7UHQIe5OQ5MRg84lStldy9W/zuo
mkRvUw7/+BYRSTkzxCq2biDXN0aCN1mBnFFEZ0iI+Ze1lMo97QOSNTVyzVl0vzERe7n1Dmxsqqsp
9acq/3yRuEzVHZJaNRQGu4+CHRl1YuSJ+mzmcDJop8g1WqpzG64eiS6Z03kUpITnJsmZMQSKcAHC
0OQGFnqw+t+mK7fjjXKhRUYJJQo64Ie0MmKhibkSiwzw9zhu6RcsC1cG5Y4cqjsxzJR7/CIuACex
ybBQTaxanFfVEvS5DDh0G/XkU13H2xx6e762vir31ltpGaiNawSjwn7bjtITThkoCSfe7XR+qRVq
IV4TVXpO2uKYuG/eFE87eN8f8eQvAi2t8Ube5n4irbPPPWLivui0P0EV1OpU9P/FN6IXo8Qtl5Ct
L15iMXyniqphr39pfA/YIt7WJAXX977bP2SfSxIDEXUSGqMeV5wJ2u6aVQaCBOO52VLWGM2zmoEL
raAbYknmt6drb/YVairDMeE/emqH0ycoaO77xfcSyQUijqEvvI6Hxw03xy+o5n0wH17SSV/+6CJW
xb0ZYiNGSf2b7OGMtAIp8fcffhlO8uGlctkX2IUo3yREAAtNEiH7JItCcTY5fHUpIn72UVAKuNXD
Wf92BC2QPf7j7mov/goo+ZHpwZXcFXxet473BajmihNU5fugaUSFRJ8ulUFgEptMOw2LuOPnK44O
bHyhhIdYjD2LmsLFXmXhsrOIccgllWiGrUnVBy1LRo2IDNegVG5vogbyqlWw/Wwg1ydUnlxk9zJ9
BwempgC7nP3euTrkVsrAoQEH9I6OaFs+UOAugSL9d1dw/zg5uLVjwIrb7W9YsWNrgIoWkHh3v76x
zLtj7hwUaG5VOZpmm/kUoqHYo6nhEG5Wu4NeEM7DsFBSoA0OfsB6U1gEEbv6DPm3UnkY62I4u0Fr
XuEE20vsf/kb/6dhgVsIYHL1zYrfJ7JhHq2fPfVzWqOmCqRpPy0djBRsS9Lc7PkRkaOphnWi5nnK
yQDBreI9uXIy7yspYGUDfZBblFR9OluWTXJTw9tFLrVlIhaZwKob7Nv71lkx9vANrGzzLwYegYoz
qqRXKiUY3EPANGj7lAxt/HW+p5c+XfxrnRyhts5yJtgFN7OCgDvn11Y1aMSRXqaySUIy1ZnyUkYs
Oc5EMIn5ywo8qYJkgRxL5Op45geNN14JcQ6NS/RHE+GgaUZKeG53tqnGGwP+sEiYbACHPTcJoWEA
rtolSvqcWNeeXv/U6+f52tbR5Ie/egsb9SAkzM/6Uv/8QNZNQQEz31T6EimWSWD9AHx8KYfM3rhq
3rD+oiyFCeTGGtncqVW+SBdl3igERTMi+zQnx1dDVA0J4xdRYAI1xdbZYRSB8gH0fVIdjYDMCrG5
CkAKUidS7H808g049kn/spTqNMkZsfGm3Jf3TsVBiavYrg/ESB/0aM1ge/MFeR8mv8HEDMFwhFuR
9TE2+dmEKVwC0/DMROe6HXRJRKW/gMM6LegJMhT/RQXzAA2Xlv4FEg9a83Z6DK4zIxvg/4k3yTYA
c868EDHRztKUXTYsA5R38TWJ4w+yS8XfzwRu/4VsMJUtRECq1nQoq2tPVHUW9rEYbUKOhKUOdV1R
JgGGDiGU4fioXLj69xQoGngJCyO4ZIrgN4Mh2OGQGAOesznf0iSD1DcqNGLGGRzZ2Ftd5RVTY0lt
W1xsFPUfXlLZn7HnKd60sEKhMI2zv9428AEBgXEhT4hdDITgMn8ODS6wLRz7wiBTGc3BKDYrBhnf
idUkwyvmfrSencxm4H+N8phlFtISkEETlU1yrxrbzULvG44KPuYi3QpVvfqCpfY0hBWBgJI3DMsp
MQmgCwRfC33rhm+zwvQqWBdspty3DtO1OiL6T5i0/A4uQxcMnZDrOVYro3hq65K6aUPjznnyZqVB
uDIQxxEmNJYTp6Ym92eDLBMe5SOPue7WJxoLQYMHMStmjkQEQ704mgQX3buWu8p8zaoKEkQPNo1v
+a4wQ+E4lSESaa57YAstywFecYM5/uOLaKeqjsQJzNNj+m30+839jPkOrNlEKZuU5wojtMBmCE9w
GRFd5t+Lvqkpzx6pnxZq4QtS3lEW0c1pr3wl3xpIM1MhOEglAbyDkmBhSf9IwgU9liQp2Bt0BKlg
bqgD6A+6EyqxPoZgOsUZg0HJiVyqdqmRoRFhUsqSnZ+TsCXvA+WPIaUwBpa92sPvONR6ax1wGxHT
UNTN3rCaYm575ECc/9d+T2aYL97dQXWj0OT+vSLGt6pt/gDNXBQzxysMjMV/0poZBk562WaSA7Ho
2w3/ANMi98RP2UXnDR+XAEHpPV7F0tRkpVAkirBXL+4Zzh11wpKYuPK1FDRsWmsIX9k1AklwqZCq
+WZz9BcuIfK70FDWGoclnoTs8gmrDGmwjyEqMEI81OxRbI6mqRFD6M+NIvZ5N8LkKzPu9uOJKCTj
iUq8dJ7CwtTpCjdDv1xtM2Uo/i9rhylIK7N4S6mgQr+JPpil8XQXzwHcG4Bdebu0Q/Imy8IWv98D
dE0Ch78kpafH7aVwHkveUC99FUZC4qsAfh6Mmv80yG0OUaLrpiUvfQkO05ookY6CioOyIRj+5Y4f
2yk+kmMWB4B1bVmqyVCJlY9tZQlLN/NrnXddED/S/ZmHeSmvdkRLMTYjYlRqNMCDDux9+ZSW8gcS
jlcKQkIfLkS89zFyY/PCG72fqv+kiHrAiL/cqoJQcZeOmpJt1+Opclngrb/eKD+ztU/s3GM07H5c
RV5vGmbUFwCuRjjaXwBKdpd7qopUk0kuIcX3YiJDs506w8//0QYAK315M3kcLlSMrOwUfWn2s5PV
R6wwgGWe9Ux4AjV/TEaNLJlHnHQ+uBNdEMnWYw3QAJ1UGNMFS6lxsXEwBhQ8eceWIg8tDvmFipvW
/HRo6FFN+NDatqjN2mBxE/d9GwmmGhr2glJRr9NxXQjZK9eAWv8db+oIvouzOw7r2afffMI9HQSW
2GyRvSELKn0XDwg5kM6PkcMqf7OAMWYP7iw9EdgTGEdIsFggjti5zlP1Nznl7cGlwQgish0rOzHp
git8aMAekCOocdvfW4haJk+og8E2ykxfonjqWnjbEjjM1E8jk+YghsQ1U2kG062mKMBjKs0J4ZTD
Z07w7CHRgihde9rJgABwNBa5UBwMdmBwUIg6BxiWak0SgPxcrCBEGabS/a7HG5cSBa2Cz2NagDAj
5W2xy2XLOG+hnQqfvIUICPE/Uzh570T+noMTIUJarG+fZP8gvR9UdinywRVGetjyKUP8f+dQLViQ
hksmSorbYKYVX9zzHYntW7Qh/I7E6GIqx43V/Ww8Z9g9Zg5rGkGn3JsFEPwf3X6p8UuVdUDbD2Jq
xVOPF5oPbM/GzNCUaGpsx6z/Ov+eXit+hCLGefrSXH43XgsRIHxU6jGLjJfsBQ77LmEdDg7XgGN3
Leg5p2ColpAFEpQs2m2pGSFWYmHqLRkxzu0miOW9G1A4lV9nQxhHyxL9ql22x5wv9XirFNzp3r1Z
+J1NpnR7QufLCOOab6Q2m3jfp3OJidxAp0j/+2NQrU7y2IXGhyz6x1869bH1MEWqLjSGlfOHUAiD
n+8SwIXf8uML9RJsL8Ty8Y79blNmp1ySTxQG9hC/PTRYjPXNFAeuiVL9GMQNHfWXjbFMC/6t+fox
xZ0PdhxrZXnmZ2NrWxPtaYgZHFFx/tbTsceR8E78GjqbH3viOcPLvc+ubUjYEdVekZqRkoJA6MK/
4EDor4CXzFBvKJIr/8IFBMw0XGI7Dmy8u1H+IfJ0VVbFQ64Ny8EK4/aFkU+FmSgvgTnT6Tfd831f
Goyor2cDnICFIfnpFjnXVJBaqpZLKJOpOWyjx6od2Manh2SkKhUHSHj4Mexdg8Gg5+UiDYdop2r4
rkyD1cgKSgF2bGd2l6gMxadCx2ISvFaD/pwtEb7ex3nePLubAC4kRZD1CFsHLhIP6shQsUhMzxc9
vK4xFiI1sng0SycUpKL45faSJQCBaN/cbrF53/DH7Gnhl5zYz8BcV+Zb3Di0YFDnRpBxMkwTXoV3
kd3InJjD713EHksGhgoCB3zenkX4W5JuFwKIdm/iRn2LYPKrAKs+/Q/xuiAxrGyJN+QtgxaLYVXf
fykj+5Wu3VfoJZ96zpRZuOViNPFR2/YwaBszMsNkd3fAO9pxkYrsSA7al6v5iWE/kr4l1mEjbDEN
Nf7FseLP5e7f91i8LfshIRFHnlPgmsWYtawDcSozWl3KH0oVOwUXlZYs9vIacyWzFV/vlcVHwegO
fIukVJts+DSwNM39Sm+KQJFn1KIBG7pPJXsZvaig5XOWH0JwTOkK+ZeDIT1e6uY2tvCpvirUHtrc
xcjRNq1CuMxnagBprgzrSaa2hsFzNfEwuq/NE+HcVff1cZ/c9eLXvjXpZLTPXy9NGmI3LyP7aStp
cfx/prg8fn1QMld76hib7L1K5chEMuRJaSEAMRKvVw6Kp6pGNM6wJApIzNlWKqb01Wcng5iAt5zn
5YiBRUOexE7R3IFwQkV2oVB1QmudiWJazFAxS5MlIN53DWCqWzHKAGeqQtj273RkB/LLeArsmhjk
6RSgEG+q9Vzj3Kggm+Kxb0gcMPDkZ07HMy/v8/lGKP3EUU/9L7AwanNysBrQhjqxMNzg4pMELNT/
PyGEbtshXVJfz+Gt8E2zFapXziMf18bVShN6YEo2xl89AqPbSJ/vrcZ2EPNlrGP6exjPbvuWYGLV
5zUQ/QDP0MUP+IfWy4HS4lN8oHfJzRwM+UCH3mlJeG/yewYsUoWL7icy8CSx/uJtBHYHbR/j+YPF
oRfLTiDIk1t5RI4PJ9ww6sT5fUM3NoRF7vfe+D41/9wl5eb/NLWGQ52x6dWn0fn76pcRG0+sUIL8
wlmQWb9NkIptHpGkVLPM3BFViQZZXoclVlcXIbbfihQ+Mw4ReFF/spg55gUz/x2cL/P5ZK5RlCGR
FlP0ah4afIZ4aSmyYG8jjjaEtL+/pln6CEkG24yTt30kQMTmYGugU9HzJCknDhN3JP7BlnYP6XTL
95yzWkVZPhji+3r5y5m5IRL3353cS+mKMGKzAYcaZjv2WCUzpxtAFqV/SqQ45oaJEgJMaElKHcQ2
12YeIYmOg4AKk3QGwpX++66HD7p9PZUg/TMGrnhwSLZMnZi66RiCawDLwYd1ixQn7Uvogq7kow1w
hLZ3Qye0xixVpNKLB2d53Tz5lUgA4lt3hUAPBGsv35ysngu7pq2LvxnRvTZIQASF2zmve6hqZbH3
BlGlVRelLGXYudNVO/ExFya2Xe8KqOiVUffAQX3Z8Xx6dg6uYeTS50HulB18xbVCoEKu3tr/108C
gzzQzacAnr2fvPB2bLjozBVVyLY//zC1UgaJPicmC5EdGPqHBbYsWyg+Jng84v8Gwg+UhyerhxkU
h5FXjLXrpcGNpfCanNM2VNZuGGXR8oR4YfGjXPnIqaFOjUvCOyaJqldEeKnO7vs201b1267G2dDX
USLHSaRcwjc8uRG6WQT1GeXmDmkvnPwXrW1iuIPWd1NFQ2E5fjhkDzvKRfhn6cW5kX6nRms2mO3v
NhncEDg7br9aoQAj8boO+VMPlNWC8h0xS3HuSWBl3Gw9Qov76Y2UdD6xnIdh+pMH8X6kasmg6kQo
aselj2Ob3x0tdlHRPaqjIBU4/BszkBRTMJAgSzNKe1oTcBz0PTXQT2RN8YKGm+41eHWwMGIu8FWz
JW2svdtSfQzDQpqpnlKie22rDjUt4YbaKfGdlhahrmbr5xrNEOfG2Tpf1BT1f41Sh7tFBZ60KW6+
yhRJjbdVETUZMxTggWBQ8u+x3LU+5d14mSeC/Hiya5G+lbnPLDWdudjzzHzrJQtPfEg2A3b0xH/W
Xvvp0mHvfKU7TtwTZe8N7HZAPzkC9yjKxAkhmzDV+VuRTt3eHhTj/unY8tslNAz9piPt+gaBG+iP
uxsKrJMi6BkQMTaXNIHXiCj9HBffqRdWpG8Xxp3tP8LpCYoLozPES25sRfJedikRmxtLMlt/HbzK
MH4KBDlm/1q6GbSNbwYLtDsJAZJjQVyZ9x0Wo8ZHo96N+0ZOC5tIb2a/XOGuKVHuhiHYz6PMgGGZ
opdUgsJZDcRB49N7Kd6ybOhsWj5Ie6oKw/1h71meSe7bkP3KgPndG2p9flSJRyqWapJv65eFTglD
hy/7t1J2meUs93OwrV3cdbKnRZtSvbLrDAh11Qyovy9UKa6L8nGqs50p7wfKFLZO6ft7tkhWetNW
OPos2TZ5uCEbw3SVxJftdkuoGqvmZV9PKeQelNR1o0kgIYmhie72+hEsRNHp1UcLs7u8+Vpes2X4
8QqVhlZ49lAEiw7RUo86OxQaPun81KSdogmAdKyX7oz+/DJh+kAxfl/o/Oau38adQ5lCbnG3oxIc
3BKz5tAxYyfIl8TShEMtyBkrEBGeynD7ONxhuaBHYfTWc/VEcwUzGVyBN0LGqn0gOc5hc5igZHOI
n++1jSOBNyYWIUc1pe3VERRDYPOKFUfK4PMrhDKibhrWZBrbodyE85AwlwaKR9gBP758RTTWfyv4
J1TYh/js5beupt77pVFXkC5tmRqLAVFyI0hhyArIZkgiyEtkspqW8TNOC1mUVNqpAB3/JhTWAwVh
fxYKS4ai+A9H8c0PFjlaIMVF82rLK4pkp6W4yNpKsG19M23BzNvavOJGQVpa2grkWA/izOo/XSrt
16qXRt0S06RHjMEQTMCYEAZaS1SZK68VkInjqqbO8ZyPAQPoyosgOyYmBjwIB7eKTzz05zGohCXc
EyT2XTlGW4HX5Fw69ChWB21Nkuv8xVQWXvjYQvwzncSGUlcMkxJpn+SNxJAPhTwQuVZKSapuv8z6
6OectEUFdZ92vGPRTnXJGwwriIJnNk4lB3or02Elg3GAxCHryw9p5M86VCDV/LnZ9Rk/s5qNYqnz
2nHQ788dsDPGrJwQB6hyfvgLkUSjUXx44XMoRzA2YSVmjtHUwBkeoaPk3JxwHSS7z8IeJggx1a8G
ibo59AdJcvEM7OOIvZO0EPRDXcRVGZdsQ4o2bcv++51uqdmCiXuwfgxROwvcZPFYprZcaC4FOPCc
q16M3EnKrHocihEHqrTb8lSFC0ov/S0nUP2hXvCMaVIdqsDcWB6yMnFlEyIQYZUUxRWHbeIS9k6J
xijAhQMdJJXu1c1P0j/NBWCEwI2JrmajCVjLPSvkFIKVWPBjPKHFveuD7Xr4KVOdnnaLDjfd7vc/
WiR8qkXta3OtEQVkTq7fXNvPRZu4AVr3T2spuVCmW2P9SmR6ZWtqoW72O7f0btTergtB/ySqjIlQ
wv5BZ3g8N6vfK4wbADtRwVUFcw+0pRRIzeXBXWmqUqj5+XRujllm2vgNDoeTMPz03TQwOX5bxrVF
W/D98PGcbVKWI1aAuUhvgwSVdgekUK7EVhFdV+xeOAA4RqatHgzFtFl6IZ01NlSSCw5YXGzwMNkl
BGfxXEiBO40mbwW22qksoYx6nus2P9GDIYOB3BiCygWegTRzyNdbGPjhufa1wiThgDe2ESC91DuM
69NxZ1sMz2eBNkFFyRpAYwCZyijUjyGWeMeutNglbmH6XEZnnyqw9f5gq9lj8nS/vUru4lLOA2Zq
qdyrC12SMmJn/Pb9ITMzYTyshoqCu4MSdaWy8AnoyQCjCBndleyAOmobCql55MOVcFtNk0piHVjx
rUsWPH/aE8vYRrsTmxnzBWk0SIHKSBdhQ3lRFFVO6dv1I/8+d4nME+ya2aUwYXMXo5H+FYR7nSLL
7u80QrBLuK8SHhQ3m61Kue6HOMiAbMRgyS+1ZhsxUbsdMEijay9ebCp/kFb0pA1C923ixqjVxUKm
3u7pfMeKA4D2CcDL4lczUm0S3YuvladMCiWDmsERIn4Jqs6oVi7gneOlqGvXMmDKkUpJWF1YD8WA
ve1Bbz1yRtMECMYX9gUDuJ1nBS/m/YfAk6D7lgi0REYbpJcH1srvqN0cY8mcohGsAB8q5rSJa0N+
2vX69zO3u4dpfzajS5s22BDMUUrxvoHGGWFHXQKjyY897ZIJe0CMlacMsoJtWLwMXGEXYfkuOYKH
FhkrsLVOg+fdNsb7D/bUQ6lECFjT2IDGN6a8rr9GIKhBGWfajtGOw1IXpemvni1ov/fAHB3bFm0t
2vQZ6RE2WXj/J2o3z55HB6uzcab2MvCy8TsEuruxuyfY15Grw8twsF5UJKgJGa6HP5trpjWj5FUm
9RspkTfp92PdH4qJkztz4bp7OpcVKoODpNiLzPJc6+ElbWsxsDceP1eaDMt8PbBQJgTy1kSTcV1B
GjH1zEilIsxqr8C3IXS98MU2ObocOGmqvxdkXK0t6AH2/CYjwcQ4aO7yiHXpFPyWgY7ZXr41th2V
5UCUx352q3teO8h1NLyADbfjOT+cShY4h6hF/3wBDmC4xGr9SBZLZbECYjFOkfr2DoFhxxu0W3fj
Y3DSSiNqeJat19E3H029Yhptjf26HncXLMdhlBqUQX9CXw6g770YIkqbqUbO5+Ps+YsKRb+C9KD7
yr4iwoFgDVtLhRAWqitSNOg4J6AHN/xTmVQ49BXgnq6vFLAtBY6ELii9qoLU3YSLo/i7siV8bFgE
lxM7D0o7wqed7r26N8r35ntY3IxY4ueQyf2h54VeYnNcSW2iWv54sZkIDCdc+7tYmh3QEYpEsoYM
6sK4Vj+rMQRMkGid9X8VNnINRj7bmSa8M5VoSXoa0xtWzHUEDfSpeL16pwIgZExYSHGZ3dD8EvHq
8Vu276BJXm5pMirU2xWbDb9RhivnA7i+AjE7zbg0Dijdf2AobAipilRC3SxuJL28EkRNIulXo7+E
q1x9LnwHORJt9HOjkUvVtq11X1f+jvHvaT8/TTolfNIamqxSe2qpFTuVFAivmUuqSA2wT0Q3jOU9
VTsljdmUIfQSmS8bFWfIBbdNf89NiiKTB/KkYJyeyVnzytTU2q06CgJ+h/9s4jX1zDT2U94SFfRz
2i2MQI1JfM56ZDyqlZaQYSJmORZKIbBBnK4QnrhKmllQiErwJrlYbBfRQn7ZnspqY1WE1SNx0EX1
w1d4EXB3m1xLm2i1duTUHyLflOnFcdTj4vR0ONa53sER5TrJiWdtMWW1h/lbLaSGF3TU2RBNDrEP
/UEs6yVGpmxVVn2hpYtC9XUTn/EU8XTefX690I5Q/vi5TWVoIdugKV/i5T8NtrZVToYmYAGKcPID
XWiiNoojBqzy/JJCk/id4dhJtGUSnkp5zrlDC5SrtF+3STRhndsUWYpHub57SSfyhCRjqvNO1v6+
3H/pwMvrALhShOLG0IUo2zTGX7OdZD6USv/LLm/4htpT6xmll+E5UK1RlRRN/VA2/L8fTWZ5RJIU
m2qrByXx2IXNGUS+iEdgQrAIGj8VBlT/unz3Z1YYztf0IFwFQz6cT3RkGPel1unrxCa6MHRhJ4Zt
p3bw0ARVh2LM7lxhotSmTXuuiNB6qSIhX2RPyUM8CiZn+g/BoYftg2m8pHl0AILQyCvmjY1oQUDW
AHrwVEt1/abGG9YlaEkMJ5L3/P6b9ZwBmx6e5VmI3pxD0R7NooE/+4tsKO2VMkIT9YJmPbV+iAAF
k403ncjb0Odknebtj2k7GEmliKCTAeLwop69TIXuEFPnk+fA4Fi1/d95NH+XJwEhrELfwy61XQRd
bvnkiWIFRhfMFWkwugd3xIrNPUWtOxHFDDWfC8vGYNIkIIL0y6SfjDJUAgoS1orL38BMQR7lC1UV
lfw/uHJ2wAobpWtcSLImUCd3n2jTiYC68nz8CfWmLfiGza3vrWF2oHd1F5+R8Bp5OzGIm9hw73Lb
7HvaeRJ118SQFiLVBt8qRI44LsT4fXTEw75/gVHdOcpYUTb7DWpjNxKgCAW+CuVqwVCC3P9MRnAR
HCmJujom29AObAl4ZeqaMZd5ZDZA+xsAxaxwT/nFUxhKZxQKxkI2qgk+bysZOLqPZWiasc5bI+2p
lxYCtN0yhXGPFgKlIjgbV3QGQfQGQOrdWRaQYrbOUjfrevN51nkHTjaLHBTt1cl6//vAhlt4GcEk
26/jjPHGz4VNT8+SkpkRFGR8TQevlBfgoTVDajovRTOdNqkRBRqWX9zYnIKgPBAObZqBGL8wV2cQ
puv7GNIF9Dwg7emtrBLS/BdX5apoGFKJSfUJRxyEAq04N0FN6m1a2NuQ3M9z4k46v8fWOK809Xvu
GBqgWu/AqHRvove/TVZKmzZ3SHLWOFTISi0DytlpeQiK14O5bA2tmfBXAl3RXOVZBVJjyz+2opEi
gzQYl0VTK9vWrDihJA6RwgvBM7OvRSRJcyIYIiivgOa1/EGFGswd2PDXw/9mKPLSyK+8UMMVh0wU
hUOp2hnjgMh1TyN6eXxevWMbUF7xjruyGJKe8OJLsJ2P6lIK06B2BtJ/4ChbnXUmVMdCuzZRxACi
Lt9Ef30EiNxCPWDPp+hPvaIaB7e8b92Pv+F9SCwYCl21RqJhr/3X/dxvYzSZOh2avkvpsGhOrId2
3Txs3KrMJoxvweSKgrwYfxLWLmZ9ck9hIhu6KYQZiJUfcWKYyvf2BgL4LsyloCjDS7pB7dUZAhOX
J/rSC2Ob9NRilvsjI1vv8o+cBkqfLFTweWYKHM8TlD3NFymxTDDKTYzxsNvDgvZ+k8z8iueqglWH
ykUwYvs1p9q6T6U/dXu3dwDB2gjzVqhKwKCmcxXoJCfDVBhq1WXVzJhHX7sDWvDYVbN+h71tjsEA
vHddX+u434Fm8Ymw/0dk6Y7NnxbOtkfQ9RN6OXueJ4jaGqpKAi36Y69lTOrat4+7dZuJ+H8/JDHf
lPDttaDJOy3dz0FSCOxocwEw2dwkk80j13H2BU/TQaS5EBe12q0MmaZmMgowSEpNkCoavCnw9OlX
72pI6ZqSjqmD7CPe/EUCBKyMJG3RqiJS28UtLlrVYZATDk1NvMvBpxkbzFQVZ+/opBodGBEqSPPc
wzchZ7fy2GE+e64iR/xnx7tWxohjoPePeUqZT4GthJtra2FC7Bh42psuyxd6lv/H2W8yF+81Ow3/
YuQihSrr6vVszibx6nbWtClOH5WrdiNQGh1d5040ZYgDJQ2JPI9tZhDMIO34VE2lQxwgExBRCHRD
s5gbQCj1izpyvrupM/NReHNl5w8K42kGUhCehhROTtsspg6YQfgISGpwuQyMp+E64y8L20VR4Jk0
U6XZ8ijECGD09LJiXjBPmmcWJe6sw3ZJ+Te0YWVjBbE/b3jNbWMWHHGKa0DLC9gJHAh+8jM+8ePk
1G76U6o8EwVTMf0gtFfXP9ak0ltr6ZhzLC2fuwmTs0PeRnWF3VpTxWrgRiLeNzas+zdLD5BconCJ
+OHywdq+eQtrRJ4jrb3G1llEKHIouf7i22SaRBv5tI0bZGmFpxhIFXkG+eBYrme58r1uhboFuDSz
8QXvxStRgu3vYNk7EoPyiYJ1FmX23a7FOI/n03IBEA8b24m5bFGk4Q7lH0O1P8H/V/z8yHOFQnb1
7l5leHIW6vUK3imVzsR58Miki05R7k8o5auTLyZm5a0G5yPGNUSaaGQk6wWjqI/3NuOVM0zXsWxa
sZofTR420ACNkOHlnMC/3DxhBGfUZHi+Bxxmb4o4fELxdOjm/Sb62xcYlrxjpadTPLqg13VsBqTb
kg7uLW7ShhBIirZqVPESGevuOYdkjwcRrdDoDITRULvIFic0ocw9p3IjWgRFA+WH1yKE8V27dNor
DmoYxYgUaSERSM4CS0JTrDnRNUvWuTn4TfeIFQe5O5/LmB3x3oL5ewV7tqJX8wv29o1W8iBcNYUf
c2MlJe4HZyNQCKmZYOSXO3DwvxzRSJCcHZbi+j2kj7wFU38ZT8dsLeW60MP9dHdyfPvbbnjCVAiG
92FfeMqJpvgd0NMnDNYkGZ/OVuCxjnl4VibkYtij/hcPOxESjWT3CqLdC+gq/ZftfQJrG/DDJ/TD
9JGOOQO4PeaGLCOaY+aLDRNfb9b/gqCnCshqHp7YxLcMQzCWsWZCQRHz5S/lwY82FDdeLsnbec8j
UnPFDypELlTqpSZzz8Cb0yi8Jw7fzZTExKvP6KtchGEIXu0ie0QAY9mfZmiY3JzswoWTQQrT1BnQ
6D0/3oH/IK4cyJzuGk9HMEYUREgxcuYGbhLXuM5rNJeNKnUFJUiO7O/HN2XC972qJN5fHe6Irfrr
KvqabEbgaBRp0Ui81RpJMgjG3Ylr9eScR7cL9irbrjm1WyIpjefwT5Pmk/QD4G1ZXHGVAoZiBpxO
wwOB7Dxv2t9kKIMWB3mu2zqhx0J8ArWS3uwsgKMO1/PBdmQvhkZ+hzCRdj80pTDMqw2SDjuPCyS4
9mb0CkxW0LPbP7jqk2fX5A3osfGQPKvbynYaiShEuJjf+DEUJZfuuJ0e0FiUbaAvuJMDGWwPW/77
spOvEi6eYh17hJB4stIgEDbFiI2/SNozFfxY525kWvoyQs7Pgxu56rXc2Xem3hfcaAHxsZbtNvU5
H3Qoe/aQSb4lnikNR3Hfxr1aHo8Yn5ufuQSSMDp5eu9sdVCEL6vV1uQC3Pi6UsIY/Wf3BTKcNS2W
sXY90eN77gNasxBplgW0bp8asY5P0nNR01lDzW4+uJn5kzYiD3JtSmpgddIvyWMVZfoBPy08zN1x
Jw4dgyYvrWX3s4g/kJc9w2NQqHw2xYOz+eJYwfs6m9UZO3iYs8cjLBtL5xm/Wh9kx556UWNUkSH6
saFnZWX0YaUuH/ODev2EoofdtHnleI7SgHuGSy4vawdpCWdNDp0ZeAKJiVgB3vHgftLDN6RqTJ40
+H21d+LZ03tvguP6Xncxl1gVcBeDwRce9iFR2Pnupj5uvtkJ3/5G3MaGSMuaLlTspZxnVNJalza+
FHWg3n7C4n2tofsfffaimCAW+Bid24gwFiDyyt/hxVPAlmZ0q9BG1xVkA/wLT4mVrKny3n7/IIrN
2k9VV9B4b8I8s/KuwBDt0AjF9BxOhLLXggJkAuXsVaYGovZXI7IJh+zx+JmlqjBzbwoeVuoLCxeb
rx5Ld4GRBwrqW9eZz+7OvN70TdPqcJ7liYNokfUcgvWCaITKwjTzEa2xZtDf7F0d5IPWzZ6cHBtt
IArozv8w7G1EcHG69S2O7bbf/ubflC0DittrXYe6Nyq6yWBa1nMGZ8tUQS0SYNpvJ/vKZdIR/PO8
nsb53FegYyVWtx3CMdwX6i0nuPUkMhP2xslAv/oRMGZ28jhQltQpZRQyt19QXTDgYy+gdOW4qwJ7
jtSeawykIDw+XWAZTJvlYws9herjeg5ixquklhOiRwUetKx955Nff9Km9q87Q46puKweGn+d1gwF
4J73r51zJ4Wbw2innS3DeXqMovKuIyUgqtYeJAjk3vDLSnyI77/NynBsA/v1Y5DGujpCfKJB0wRq
xq232sDErR9vWYgCDl4Nv4fOSIhvx0tHysRhOYfjfRaQlPpkXDseOm8FZmvSURKFT9Qg0vdGG8N7
GP3U8u24mPCa68jtPEYiRLL9fKmOK0xkGS4+I6F8K9gCDvz1LUk9FtZncvt/YlMUa01w+qbMB6uJ
gXRpLuBjbpEK/TOV0nWENSgAKlG2dgufg8pY7Qvk0gIEJvucNtTO1b/NAUtLYJ6l3X3GdT/r00QB
hrXWMjCaLENk3q1p5Wvxm4IrCVicTjALpY0m4S/fHtsp2lVr0Wi354acP41wXI8xz4fvqERZro3Y
WuN33JreHDg06PFQQlrkKV2Fq9+z8PUM7wdmkc+3ZIO8JXkBH2BiqKyfIqs3N1qbsdshBrgpErnZ
2bQd5HgaXpvpdFw0NfP1UAmTP8vzGkfCy04NxzEvkQwxEtuSqO3r6a0MVEu/yOQvTUb50M3WFrQS
zmx6DNYrmDmMkiNdTDU0A8F0f8kPs16dIeYeADey5LHTxaNyBdehBCY4eGnl7mif+uOnVzxtdKBs
qrvCMiCNC3z0AwtZh7EjYfmfGFG3NBv7R5gqoaUZTYB/GABLiaFrjTRNY1t6kvrLQRfA5UAYXVIa
NPZhLqZWPgeqtfY2/+abhA7BwKUCASzVKunOlgcN+/wASRBKYqldI2AUjWLKAXG4gWYKGERK6iKR
pTJbZGrmgsxk0JmlBidTFgh+1x2L+0+EYWDelt/4JgcmpjEQJE6EpGf3wJPzCyr9NqXubkFszB0m
UyAr0AMhN7w5i4Y67xhmt8CpfznENfDQ43s38k/0uqpKzAlpOMvCiWqzn4pJuv8IWjCqHP7Kepir
7GB7zPrHQVtUO/IBRFZ1mPlaPyLNcfjrrUwXNemI40aLsAQdZJQjq2kiBjSGB7JCtFUIc23aqEm5
ddrRXY4WkOp0VtV/AYsaM4zO5D6qXJ/r+8j28GyKfL/IdgSqkMerCydokQvd7dEdPvBqhzDxHBdY
zEyQN+v6I0EuDovPjDxOUNxFT0wozjWidc0YF8aXNeP0Lba/zZwRrZwEAPXIO7MvhxYfYiO1BUMc
+2CVdAQxg8XScYwfLpcObnpoEGX/E9A0/KMO4jMOVAJM2UvuAZNOhOBn83cY1TWGqkD32HG3iwtS
sMmJXsTkcVTlenusiYvf9OuJ5ia0Pl898/vjHWnzTMBSk3EAdSsOeTSTFrOvFMaxkr3pMQrbOAz/
T6Gx9d1HcxHehUS991aTWUJAs3XPY8g4ghGaYsmx/BTZhbdNI3FjZFHlNfHF+DG69R7SP28+s3Hp
lRjTMx2By8nVQ80MEiNJ2Kjo+oHwp33v3xyx/tUtjVBYVaSV2q0AKp41RbWVhUaCTt80jHhrrigF
mKV0KkcfD2OxqarrnCyjv8CYtSl69as4Z6C8m27fxtjYg3+w+cCx4F5ExchZzWdiCPDYSrXChh7H
6u+ZOU3mK/g7WNHPwjhVyUlTeq93tw0pvpTu/pAdet5BEUzqgOF5+dPTyBbYsjiOvQPUD9N3mPUQ
v+JG3wlx9ZLwdvirDrn/HFXz+oGwFi4lLmzllaLjqQYt8GuXs2EgxERU9csbTiW5B+MfgJDFodjB
l60yzBJRJyklS449ybam32TjKKzkFBEDYl3+0yokka80/rk/jRZ+CkgiAC/707bt39nbqcHI8NBl
BJFUA1oGkbcNKTLqVib9Dof+VoYbHZu81HkQDNT2pnQa7MabStaGV5gbdsGpHK0+ARcSOXoP7Npy
fKYx1va9bGwWteQjRU/0PORipAz7rAJv2EshAHqH0SQKRG5S32b0vRLI5leASgfv0HAYo4gQW0/S
9g2hMnwTTb+YXH+IMzFpMbOmyfTpWV/8T3q3xyc0M8sq/+YfMKfEECEcC7n1jDdK0SWLarhyBnQz
3pZ9+o3wfZrj13tR14hZNS/51ftMJ4tUELnnVZ6eT6QZa/jXHfvMNwyVaGKoHkv4yE60fgWGSkHg
4ioz4OaV1eDYSvb/uOcNewTBrqeA87ZS+KgXzA3HHmQD62Q8EeRWXffaO7SAaDGt+7n+vvMn8FBs
3QI/ivJqh9oPTzdDsPNOoizRr669sLuZgRKE16TmbZlfNCoMQOEKEBPUnF0nUpbzPrmX0Ov0mrev
tlaFmvM/lzO6iBEfiMfvYOllrT9O9thxWIJHFxJQP4HgV1HDUYEwyQ06yIfLcGnLm0Nts3gx438j
Ac3qLoWSKqG5xxaGCUu4UYSY5jc0AW3TlMr29WvhGkCb8dxbkLo8hn8hfhVcMZY1dt7jFdxLF6zz
8Bz2C77POExU7SYQLLvJ72+NYqmNQoxEFJP9QK8RLs6rF7YtqPjGbbHX6DwMN5hOUcYPHF69hE21
s1GwtNq4IVx3YilpmZBqc/TPCHSLMz7cHQV+9ZDhObh9u+OrwG/lyjJA2PZq/eooP7CV+nRjNXwk
po3INTQxPoWxC5+y0IWW6miZpbgZIfs2l1kfs/b7SdX5ANbdHfhQ+VHYhc0icyHcIFZqEbrHqZ+3
dhlD99trB29/z0pJSIxrQyenOnfexhEKAUIgVvZ6xsTZ9loix0RxwmvgishZxIO/9yDb1aseWH5T
3VlK92Ersd3db/A0jMTr340KQWuZAqrgY0wp+UYBgDMX3WJgBzPPCtjrVP4r4RNmeb0FcdnzKOd0
3hF82FGzTfLnK3TU+nFFgjHNxuR6lKWdR6SuD5Llo1P6Jhvx+K/awDsUFOYKUrak4rsCN5FL86lu
LSFyJx8p9SYtK+AUbxtn1ACp3EhyjxVN7rRuSjrwvqnqQTWLAWQmKWMUiP1fzeg1ITM4vDW+cyjK
9WHQzrz/SAehOBfcS3q/Gj5AbNrfGjXuNJqgNxI9IDHQU1PAdSYWu/LqDkSufRJ9qDNrivD5cPHX
izZsUIj13Z6FQvGhRhf/a0agdCDTUWBQPBwkYzDhrRJ4JM+s3oo9/YvwMill0hYQoYgPLNa25zXL
lIGpuuej3DSFFw132k/u9jA2X/VB0Wc2aOpaunWr9IUE0KyhQcm3UV2w7S3PzVEaORJVthiY98Pr
HA9OLwGNgEGtBJWv69J+wh3ONDEHa9xTGmSjdw0qWssq3z5yBJN9L35+zhA6DZDESmZlFKLXvIjl
jBcCtkkqZ+1Iiz5np8mpkSAeGEYCxUqjyIcib2dty0oWTyGt6f3+Umlq1dvR08x2YjhgtmSWz/oN
S3RGNivkzNNuL+hGKHN69Qi7FtZ/ono6nctyELdExIji7MF1BpyMvhVHSTcMfYv6MhPNl1EaSCXe
H2TLko2vBx8Qz5lsJHBHALnVhCggsYxw2cYMzu9cuNQ1HXqXK+iEsg4qMlENBhs6zQaTq13ksQtn
pVMrerqPrrqYCja82NHksWXvluybtK29pRsF5kRmi9rMNcpN7zfRvFGbBIRY9GUHT7tiWFJ37A++
4RtOYdEflbmUwh66eMXuT2xVXbctcKIN09Vz20MMl9wDiZ0+Hi4WVruOoof8+m35WRci68VfCiPf
0wDwCJ0cW6bXwn9W6z+FYET3jzxMiM6KU2t66Zjl/RVT+g6ZSd5+Y8U+mKCc+gWA6azRJj98pNT9
xXnMgU8cuJtMyXzpicADI5bGfeXJpjiciUtCH2Hl0DKcKZhhwTe/+MUZAAIvE/ET87+9NRx3MgZe
uereGJeuSU+mlGx7PCdNJm/YdMrsxHhNhMl+Ity0mHP/OxOh/xPv4+9TzqdiJoKOlYIR/7irdM4c
jUPbmamFU8gIcPfjceMHOZxaxC+slPjUY9ggcPQsahXd0MtNC7MduLWCUdT7ItW2tHyUDar9Kv3Z
gj9YAFz0go+ledquPX6+3erpLir8tQCsJuTPP/wpxFTT+0/j8Lph7GmixFznvf50n5JQVnkFsZNc
isXn/LsU0yFKTivAzs4auqivHdLUW/TA4ci2zLvdLMybBhv1BtYvIqgvagRoUBR9uN/IfpiixoYB
IoipnmNI4jP1cSAYw0qohXxAnJfai2/CW9ssfslNfxg5WX+jCu5x45xh4acpZ5MpHuynzKpYI+pz
8DvsQEz1WP2nIBae8WeWOu8PNdqy3tJpmCpe/UyD6BwRWS0FUki9dXAj8XoVN0cvSGr1k36buDlm
KGr4eXi9s8Ne0TUfG1kofP8KUblw/qFARsxKlan3QQsISZBSpPZNAonhZENfij6bWgiIOQOHFoSJ
XmjtFNl3KrlRwg7x25zisCuXjvr+eOnJlK1hG0Eo1WtLlGg1C0zzl5QTmMscKORT7ZW4jAwFpQBN
D8v6zXokY8j7dKkgkNIvdSi+CZq3D70I6uWbNods1y7e4MaM0IT6YMxHIvYVttis7wzjsXzH2QyE
3m03qxKPrZTj/2igNhAqwMzORa4X1VWFc32+o/0ScMYUepNILSyNlGKrN+D2PMPks175Ej4zKy0G
w+9wTvaUOpAYnBctu335KqVkfkqtGKrd/Yi8CU95wHZYHJjL4NT/0GQpHUZv9QhCrsnJjtnYzC3E
8GHMoqjhk4pZI8urRHvYJeQXkiN+WCyqZ2/Vz3UflLtBRH4NdLAerhf/uFjsKIkJ09cAJhplJdl7
4fcXuyimU5xpC4kHe3NmBbN8NxGn92tRAHurxTtrvmbMt+4C8gNBuKPm4W2SiC+I7yHzHoumHZz4
BDtE0GvGUJ6s363jXWG1UXvJeHGpg7OY1fTIknu/DJwuYzmcZhB7CFe92FeK/QfoMZmyKdXOBQWf
A/IfBc+pUuwfLzCecQQgHOnP/UEdJ8X3b5KLwNQijD9cIU6sokFKUrjciPJe2MkKAW/qodla7Qz+
XxjYbkkZu7ADOYcjUWCv5hOW3IuqBHibZ4owbmp4RK3oqy19lkKr3w85yHtKmTxr4YqtAxlFV4MO
i7PlYMYp0VvkgIrJgt4Wrt6GVSX9RbGsLmPAbiCtvTusRnERtYW0Gu5k3K+z20LpI49K21XOflQD
FYQ79R58+uAYcg4O7BA1lxZ5Ep3Vo9bzxWwvKCd1OS/Ug9pNuyw71AZQVlr/5vrhBysE9q6xlfMY
JmTqKRzpybxB12++Teh+LMnubJY4Pwnbp/qA/4FYIPSXugvHwxA0Noe9Bi0JD1H9W02JB6gca8UN
pfMISNuF8h5YP9gna1HYJz4D+vZrUMs0iMlUzaSIsDcMg4pquWmtMcDVYzMdfz3ZRYUew+MSyl+8
N/twaAVom+DcBIcWuc5PhAf+/ZTWVCh0zpR27XvsgL915DMUEFYzFwpmrzFl0qTLLF8FdhMm4Tqx
4ieGSrKkys8dg8OSWotYlHDMkx8OcWndb5mJ6ccfojQbiNpDO4LKv/v3TqZMv2cTBGQCsds3UOJG
qCXfW4BI/rsnLPOKJXaPaMrfbs+QAoZLsoyhiAu4N/oWnl7LglEmtznCBmBRTuMP+hv4shcxO0PQ
viEOPWCGhV28QEYm19J+5/j8FClKDMAJxisdw7xiWDBNT8QsyPI/hHHNnYwqMW1tyJ6N9T9P5rv8
CXUYOlAcvuQTeQtt0vs+OFzlJmcbULtEIHKwa0UE0s6xrdsyhRCnAD/KQvQllMtafrBuuH//LdpR
+H/tsSbpyWwrbtnTFjE2widi/13tbxTEAxnT90dk1rg8tEs7pIjWJ7On/hK00+zZvvoRmDqoT/DA
3sSWftHK/PWKH/dS2aaWpVNWMqwEu+fMqMS7x1pJ7x6aql/OjmY8cv2aXn3/tH9T1GazMjVKtolR
FlFKuDk8SRC5+TaFCljYdjOXN62YfDrGo6uZ7ecT+mvYVsRqHcivX7qQjWPhAuK3PhLgyMixVZc0
WQ9FNefv9Iq0LlVqeUHy+79NdnMJx9InEIVORkNK9gmnExn6T8qhjpkowJAw7GvCD436LTZo4moa
wvWz0NgT9ZKYtAt9h6hm5iUA4M6MaIJcbUvxOlCvhtruvIl8t9EUUZh1Ga3mMPUbV10HWRHKhL+Y
cADp6nN3+u9Jr5VvQKmkQJPhfxr0qjCWd3prdrNvpcpY8/QgDOfAQwnKAk+ih+UL3y48Y7TUX+8k
3X+aH5bTuHmSZlGOUvi8YyttQcynQQWhwzBBzTZ3/UnC08VZ3oKmv7ZbQEmr4aqNoHspnVa/zx7K
f/D8EYljVv9sBlXeRN4piD663Za8QZHuEKJvxmgjgoYzVpevptmozFa993uiGJ2r8nwFCN0p+N3o
u604vSLR8LaiRVFCkudrUM0Asxci3fIwEmD/6OSYszU4nt2xpbfoe5G3WSTiFcw7PgE9mb5dkDvf
nyZk+ccGni9+DA4/fKUKKZzLP7AKzgKruNU9uHF7mnn3zRDZ8lBlRSv80oQZNb0TxpdWrvBQlYFd
icUX1FAyR0QVFjbNVl+N8fD187PGZg1bWCTnw1acer5LKhpBOiiFx7Qz5NFY5v18eTSTRM3H04c5
1TPfyj9OmV7e0E3+NYww+o3+3Hv25mImq6USUs9IyjE7ON5KoOBodwIzt7QOp0bKvOfcm+/n4zC8
j2OpppvGu2d03MC0m7+M01vMvv1VGeuYrdemNdJVphU/BdN87W88V8PH53xFl4e6S/E63yDOXfWq
G7Ec8Ir8PF4uUZK0nmpOYn960N0QUKo6v7O6Lnw0kgfgamWBiGxca297kmNCG3JE87yZZ/zCtOrU
tdKe7PCnRAyeajGo7Q2AqeFbLsTAsDefmbWkbMlfWNWD7fPS+XbHiLsYaGqTRUhG0J7wyPRozc7k
R4mxHcZ1JtdZqbarZ9g0T8jle4P3lI8N9SWyjvoSufEJZJ6thd39QGJ52dvPEHJh4xp0mHQBjixM
HC2eWTHX5zzM1H0uDcu3y81UVlLKGHGRdwiHAWAgwkrc5pHsYklR0DG88ErTthrYHbuectKUENm0
4DeQGJ13CtW8qivaJ3oyflLqqTmLW1ec9jU/tYtokFxGMr3DWqGhIjFL5uaVE6Y9arPnr28OmeSF
WXP6m3lFuspCTXrNxGQ3f1DdOaDiSKt/ayr1sGnFvRm0QX8t5kr+8vLsttukcTsQgfMnLksezDkx
bQo/6jxKkm1NCBkv9jkSuKawevuSloCleC03EzGwNGhdOHn0EtOyDRcd0S72xgBRT71DRXQ/yDJh
z67RzKY7141IwIS7u5638up1qItML/mcgYUngo9aVoFk9WrYkLZQMUlOQllBM6AJnS4q9jVZmluV
086T7fyjs/vk5Fk9UdyoQ6Sd2+5Pw+XSmRlNEAmdSn0qY10yWK7KTCAvaci/URcy+yuzWaalfJqU
RPbGP6gQNbsGciZVdrzurluHjvhnZ8zb4hGLjVd6Po4FPpcBZ23iw9Qv5+1RGpvkjqSzpA7fTBZn
sLoT3g7RbtvQEufnS1nSGo/W34gikmOMh2t3NcylQ+HstzbYrKPb2h/oshHK5KqvjImuwxRp6Bko
g+SvJaH7L/xqCU8WSgOPC+lRw6jMviP3KW5MJPr7el8Vr1xn4FlH7n9iNNFNiPU3kgU/PvGIyzvB
qJG9EFE/z2joxzwL7akdwAhmrDo+lR/v5saw6zeR35WT6MTbHcW0wF1O5/mQQAUjm6hzVoGJI4jg
lYZvUr6+/nWJ07B8mNtb5enSbPi2qRAx1U94qgzFihwxvzIR//4ldR9JqO08LS+TdYhWQwXtLbbI
7axXKLsrU4MwKWjo49zSJFg3TCWcrrSIKQyl3m4DAYnuL4iqFNt6znw7oz2l5miLbVc3rtpRjiqU
b/o0T0g7oDAuigdjjD/QtGqxWYho22Ix4ZziVAcX70OKw8RgOvQLw9X3uzUj8rsikuAt+7ZCnneP
QtaI8s9KtCKohu4mcrlv87w6m9KU1kU3LS4+co20gOCRMoWNozNikX0pi2JNlOf2JwC/UaVcJaSu
TQOHMz7c7lJcUDqvQRYuEOK7Cdjd3gbygrOu7c0aDw9naBp0zYmLMsGsBxl1LcPdcFE1+qtEAbaK
jeWCcohonEOVtJ73VDXNcbiPgGLqsSMp+3HID7CMvx/0XDMXf/rrm9eX6kIJfvbf1kdObCXIlPST
8kTss6MQiaTcxhbeEWjgTdUnxbGZLO1tfzq3QuuJW8bIu3yg4k0pAfFHh9zJnsWYnbTRTkraz6m7
+VsUuZS3P5u+ubXuTnijFjgb6v0m/uKmt3zjxEv+RXHCAD5EvlonKniJ1nwwDXydmJ5imIpwLH9O
WNG4b9EuEITY1wiVO0NdkRTs9OGVntw9fI4LuEvVK0jnKpBAYw68B+Du/hyaLeYuv8IayeMkjS0k
kvYDDVUoLX/xSQmVesCKBLyz1FFFvxCLZhHsCW+as1+EG2byxEobDm9k2fPdBQp4j9djHrIA0IIO
VA1PrtAoFplxvnsubwCOjRRwTN75hetWsO39zoGGkufzGfA4z1kgJX74Q7MmfdkViSNZiF2Ymzj/
VJLchka0HVlKusxJVYOYfBD7HCsj7xUYKx3FzHKfiY+nk7Tm640JsMv8HaUoca2qFQrIZXe7ye33
5CJLXwu/oWA0Y9tpiI83qu/FSjZG0jdIdvJRsnx1aCsSp+pPrsEYby7QIsUKV8RZ9x+W61ZMAZWI
WlX6oDcP+al3fV1NIpQZfedBMpL8sIt71jBNG8j5HvNPtuKpUUG4NT1Y4zusyubdP6XDRPFxEUJt
VXqWE+Z4EGmmOZ0Q6LaI7nKQBPoN5iaGE7HThbN1IveOC3lKuAFwV5qqXWcyOaLK30yP4wiiMwnM
gq2CH4vulGpw1SsmBOd5h8quEW7Te6xaQ7Avc4MRK5V+aSTWpyqbh4QNUKOp+YtvU3l4p9qQL/0d
wB9T+peQ2c+jYj6gUcrVv9JM7wrb+2HiodW9yDjyNBvhnfAr8xIyYxNWassSzOPv1xusz4ZcE3qu
38f9ZYrKBOSXp645M00RJTEaksVk4HULm5k1ttz4KuAIYmMO+B0DVuPVz5buc4CsHrkyTR6J1O7r
DAhyFMp1/UI4YMJaE3GF61VwQpbwZWizGkR9jDfEKbr0m9R7cOLZgPvICjf1jSIxGhP0LQEcFgZ7
j+fE9SJ8YDYcs718vFlFCKjoaB6LeabFexGRxcBL5Q+Ms3IaURTkvLHsTgMtz9xyRTClXOMn0tKk
3VsMzcl7G61WMVVlHh1/bMRIinKljmjaNAf7dhOjLyhG+9tR/l+ib/au2PHMaBQyvLhVIoh+sZPm
pp+ExcuZ+iOy5pI5SxIc0NSBS4EKqwo6+dAl/2PgP8Ql7qV8A4wDyRGhLk+R2rDPwXhqV83Ra3lt
XFq+z25DjSkDQFGZEw6hOZ0kV1/g3aomGU0QIxd+8s/boy89wTNYVsiTtUwOQiAelbs5lULj+A/I
XG1SVCwUjAeEPLDkAFXWkjLty2xmFaeRpP6PpgYatanyEBvzE3cGHCeYgptc9LDhbMHjYtrgbN4e
Mg9YtX4Fh73iixdZWgl3Z2UTGIOujc4R3pvZZrOAecs5v5pCxKjp2Qm+lUXUN6Rk23o9EX8MJcAn
y4T/ulNpw95t9slRIXSw/C1OLT8WFNLlWCsewmc/JKsbw864VDoACiAW5egpx5NbOeRX8hBFci31
GT9Lg5K9BmM+DqNAj6SvuUJH6pN0vtNQfkuh9qADGZ9aqDwTcwBsr8bQ3JX1AN49jYUaMvL2ed6z
lWJF/sAwP7N3LIpXnQvEN6p1m7TCADkoRRQn+75zHVVP+kZnV6I08KnW8xloSsi7yheBzrwuMZA2
ZZcMqszhYfWoCxo3smhnNduHz+aJ62YsjfBipxuG6UO/nDPCPS4IgCWd5rlu7/ElSc8lbDOcVaWg
fC3YiVgPASTrOu1bMXWJ9D08L2JqM3K+Mogm0/XcV3td8RUzG5xxpnSsgNeqqjemsbzfwxmSvYUJ
OplQ15HJ+/OzT1qhbE2ud3oVnLB3wcXC6gNVX8wYgtlgBrbHDbOxfmS8bgoguq6r5qiUbIO9Kg0G
cI8TYYe7H9WPMTtlzcma/9bHqzydc3B5nE/cEYQXIzuxnk7TOzomBDTMihMG4xAtqfrZx8kc8IXV
ZTtGqCWYAYIErMSkS2z/s8GfwaJmtOut6t1tkjp/y7sNz5fFy7yLH6Exc5viK3N0ocxdJw7AY/ky
2Z1X9qBunzfj3hrbLwUUTmH1H0i7G7sCbe5kNY3AtAaRZjtCcikUgKU+Hn+cKBXTxvBSLNGUka8k
C7tNsMxuvc5NhrclRI5wIhK7YLKwyeXSvIThk2ggkYXgwVDQA7JNkEXDEs7uNQoFHCp0hPsylE8A
9brtHD46dGP5uoLD+On3qX5kLDviG32LdpZK+F8+ymtq/eXmt7N6YuHTEeYWdBbL3UZSHi+M8ekm
p13eY1rbWqdkP6ZSKhb4VGLPuOzFhZB5qwen5v+D0FUV+OTtECOFbhIDx8saLV2/XY6a7iDaG7eh
Kns9O/PnIHFX4ushnfk/X1IfbqbeOU6MgOfC+A3S9XsyJoOEjl726n4AvB6f5yKIeo3YwRSaXBfq
MkkXfq1CO2nqfHW/FW3ShfpEfsilCHXlMqVdqgapE0ndu3ip/IQxsDqnPUym2vRQsP8H4ttDqz34
9HBZYKpaiMkhL40g/V1CDgsYZchTbYmBBd7rtaqrh4EqfiPe6kSK0ke/le3/ymsw9rnc5ud6xA3r
TfcsYOyS9k82lSvbOgiH+UYW+YqZpg+9LUH8G6OKngcokqcahvQsQzzJHORNvC00dswz2yKyGdUB
bU7YiNiJsIkr7QXv2NHO+lzMR8PmsUxfUl/YpSpxUM/HQDbsyiV2aAOVWv6cuMJy53gqTyln5MWD
2VCP3AVCmRktf6QkCVoqXjZqTZFrt1LeZ13FDYU17YC88WtSTtyfL4ab4H7Kw7T9KZ3Yh4jx9wIJ
51tEn6G40Ys1uSjhn1OLoyl0UoLhPcZsiwEcptIO2xUqKVe/2qSdnVT3Rq9ZW8iwOQTAvjxVBIGW
Nl77MQWKPabptCJMPzsbAr99rC0suL48u1bY9qddXL3FceyzIWXtrJE0N5JCV2mOQUBW+/o0DHhp
UCShsJjM0lFO+SWIGy1QsAIqtvaDPRp/pHQ/Za1C63wmJ04NhzJm65EfkQn8jZ9FSHvzX0lY7Cm0
ueC2asQpZr+rxMgPDb73emYmV/zySrMEfQGO/VOoRG6wVNfSa7yksQC8ccwR/+9SsXcfaa4rNU7N
/luuOKGqiJ30G/mkSR30NTOlOKK9hCI/x6vi3dHl7gfbTMrsPopiMfEStyamIrUrd2/JZv98YZBh
+k94e7BrrOLAz7NYLmnImwv7IPJDJsv7hBMRgssRNMf39JdMX3dv+gQd0nWEqbl3xkace/Lg7KNp
HZcxuMxEWx04ThNVU61UoXRweHsirn2qz75KZHkW9b0LUpmsFD1tfJukZGIFD8wqQ8/cKt75BvUb
bYlmvJ/czDs3Biy5EHhOrHemrkwqeD5KBQeWxaqUylpYbGD0l8xka4/xiDpZoD8Gg+QbLw6ZlUSM
NQmPJ/Cw8Q2bDjJQHl6rEyokxhhF6qSsuVLSX/Rky1Txhajay+UfbrEZUoyx56UK3HoYaVBk5P4x
IsN3k6SRAC5YOnd+O2jZ+7QJFxIXpZC0KJXeevgLcX/bYg3Fj7Ziws9e7c7kDUcBo4XZ65hLlHCq
jYQgdAQxu2BWOd8pVh40BtDfgNXYAfLNYx1cx1H/MFJ253Vwetb7/QeAx4BcgbjfuYly/L6K9RfP
8iwNVs+pxZfdC0jpVxuWb5NZrgNjBjUTJtcXACrZTrD/ZhakxaZdzq9tWkokFxeGgEkUmI8VRQHY
VdacSW0MwXpzCNEt/Zlzdi4yys3lo/kaqwIivqXijJTjzQLmEpTcsM/pbOSGgVZCq9YOfSudOirY
Ou2uyneLoYybXiPMJY5toIWeW9DxyIavVJlZXVuRCv/vdw9YhLBPK6uU4HlE8sYCg+TneaA8pz2H
hfEa7mMfzx+uoFguq0KG/PPRVcH55N9E3TAmoGjYFegzCeOj/Nh57F0QXTDTANYG43UYKDkp9OA2
+PoVw4R0eh1EVSv8uhlzeB9JTsBYTO74llMCPO+wBenzlQtYqkSM0T6DA1Yez2yK8YLRdLNpuJwK
oBDQpISW0iEJ7Ij18A+ZsObbs0D1vhmgZV85DTS/r1ngoSOTSCUJH3Npmx1AnJEXoDvqF5SnsnVf
MZfNPSXp+arjuNzYI+e3KsS8pnS+ReBVpotLJhqi6Em5HnXoBEepweeIBQ1u0x7YCv2N01V3/0Av
hC2C9RWGj0zNnSeW8QOFKitEvjH4eAg67GHCH1tPWeEqxe15Ud1IrWlPIdIEytd38rk/I+igvjzk
z2YblDXfDDcD4ulzoMBYwAv32JiKhHSv+FFltRrX2VTEXWR3kJttUX269+gh4fsspZLA67O97Ck4
++JCWPAPkI6BIFEK8gtxa6OBdifeiM1nupqLSWaOoaq8ZLCe191MPOWN2ZYBw1ewk8FiWa3uakAN
WSKjmv02kBcQEqFZmqfo9OE5XlzXRxO4akvMIyxHPYv4BL8tQeXMY3VBE1HXnDBQhLmV86h51+X9
O4f9H4KrXdlIm2HuQL3pz57Gn5QTl4Vw8qyVo6RuQVeGdsQi+h5bZRSEhVM2wjE9TKWCKJBJs0G7
XglJaC1IfvNETImeuru9LeS2xQJzV1s7XL3z7BaACy30VYv0cKngngcUzoIDR0vc/LvF7B1q6gSS
9QtP42snKNYgwNMxxBwmpWZK7LEhVtcGVl/85nnUvJZmrgw6Gpko2pMYNGRWCpLK+xFwkdk+7B2W
xkxee8QbIVjEP3qdlNmlxLudpEit0QKXDugCeuQW1F3YEapR7xrqwkHpOg+7d6RLjvnm+0Bcoc/B
WEqJJNilTpJ/Ywl3dNSuboymGaLn++CSlOYLSyIL3M2tIzAtGqo15Oq9NcBBOCT/kXFE6S93yJvs
MJjMVQh3LvyZMequ8QA38exFoUzwIgjr7+32cEOC3QOvTk43ASHOCn153KvpHLMQF30m9VMYbuLs
A7ETo9/Wnm1YUxFzpMO3KcbWWJYBcRP3ZDT5imPp0OG35j/op+unnpwOaI3WuAS5YtopYmMFJc0q
qu/3RCqBra38H2YXbi2RYEeLwMQ0UFxBzkzxTku0OYV98rXaBHJs14wcaUmzVdRqh6LgqVVRqYG2
363XUf5LjI7DXa/ari0wcPLb29sX0dcaB6kugvfXDdjZ0Sk4HhNUyLxs9eEtbATnkFuzJmpXsbge
SF/HRz6Nm3WgtFhTnNY17b04mfTe33yUUZFy26hsbLazcqh2nqCnllax7OjRb+jkn/159nD84m9I
AJkJFUGgC/4HW0Qjo1UHXXd/GEZmJ58NzgwSmPg86io9jYeHU1pkCyqzvSroz+cYinDM8brH9Qjf
kO7Kb+zIVT+0IW1h1oxfo1RNTsd2AzbZugW9W4q2+O7YMV156zYo06EoS1WOJifQR8VlC7y/auQ/
XKW1kT1jnsDfVFPplUYHYueU1CXx7sosCdHAN95cDFh/ro0vEjSjeQphgyKx85BS3dLqYCLf1zS+
tAHWOcRXdDqvZYJnaxjwgIstndL6w2q/vE/E3ZtGrq2AN3t/vrk27Y3V0ejGt4ArO+IJjjk8EHVL
cF7lG598P7oIKce9DgI9uTEQiLMyLX+wBFcz4eDG05XmuMxr5QlMSU23CsO8KmADRDnc2ethDsEb
DFKXdf98iqdb7cQ7QPCJs1QJMWcIN7aVeNSwq8DrOBn36jNtrD8tDnYUKMTi43urXVSGVWRZ4qDr
O6TU8JWV/6RUNbE/1eRSDh1/N0AoXAbMPi/58dXAv8UaCRiYsPO8IxkmLyW+e8p/Ubh86VR4WRnr
EPxvBSX0e7b1182sCqPz4yY2ny8/GgJqZbYmiHA8fkvdDP87nFiXTHsgmzSfbiM63EWHymMaQeJD
tiISfXUNYKdIjo7nV3+Zi8hLgrU7jQYNTtGZ9/GrKjXvHpLBQcwXiAgWziDnAG1ANu2PXBP90BmB
NHiZnG5pIL1iz2jtEY293otvVcq2/HjHpLufj1Ox6//4sVJEC1sc5OVjMkTJkrTQlOIBTCC+/4N3
MudeNjwQ2BwwZbSkZ9YtyzE4rf/DuDRFdUYP5P+/+boyJs/KOSWyFkEJww+4EAt1VHMt8jNaWKS/
wRjVdinhDUhR00mPShRmetXFo0qGulizwKCQsq76YK5MF75nq69cW+9nqsh6/KLSXf7Z7aN8O5zb
mOBSzdxGmJvgCltoocPXjoJcBmYXiq4EV1+/lZqYPuVQgznCyIth3upGcm2wtoH6vvRjyTDPsACT
8W92IO3Ev+gXr9kAf9vu09QoITLNsZW9OsYpGNmC+C1FsVCQDDBli0CNiFawvajKdvshZVEle81L
33ELUO0C1L6gxx3Ce0es1I9/byTXA7kLIZ238iRdRKDin9RGrZYgZpiyfPQa8m/6vOVnIk40m+SC
BcT/SWxr8nSwsTTIEtx5JXtRVCmZasYuztt9YRLBHyGXxuBq4gHDgqCbT5/jyrR3DL9NTWYbt15x
lWv/FXbQyz6FAmy6QoLr5577v94bzKGq9X9G1HU0EMZDjmT4B8RZBhXoxew87S48oCqU6j3q+cwn
4xzx7IZCZnDBAQir183h4LRW/Q065ZC4LDHgc2j646EhisSEWvr/MVU9CGgtc4wlZ8zFgbWTdr5n
1W5LQeJX2cA/MXx9+F/mpKdxOjgqJ8lAjbgPVPLgdL5Lv93odV5dBtn7l0hXJZN1Wt9dCqTrdYPb
Ay0E6EaI2pGXGeeezGOjwt3f+CUTlvJC9M6ecIqPQAAq1yUqMsvY1UvDvm1SekmYcjsnXmT2zUbh
HzBma+Ah1TQuAEATk3DA6OiQeIn5CLwC2HcNWiJewgzeh+0mXOPk8o/rfUm6uGKJ+j4Wh87op3vg
Kxmo0QnSV2t0DwpNK++86EonPfVxH185kPXHvmOs+A0KL26IHVvUJuF9/FIzQ0/PWvvQPvboRs2S
4VYTaeRyBXI5ML9dosRwCeiyF2VN7hYLu+l+W/i/jxNjb626lCMG5RF1KEUFSNijwGWq3/1llqWN
frMQ0Kw1ptmCJi59Bik7NBVhahPVJ20g2H1a1Rh4x6UmgdEHjOYFLrUILChsKuRP/aFKNvhGOGN8
H5b8MK4YXggbPVe4+SGdci4+2hCPCQkl9MhjazkVyQhrEikk9OTMWoksl9KO7eJAib37e90h+xYe
XxYjk9fuIwvoiqMrsvbw0TlG8wIrcBNvYAtJyM6jbgeQ/Y03hk5DnxxoNGNanQTpz24Y+YGT40B1
tQgx1H9EnoWXVzcCORdbFzhWp4nm43nPcY4QepP/Jv3TzEq/lq6qgouJ17I0shXfspzqQ89Xv+IX
9uslQZXFF1Q9+ZpjxULDr4rEIvcP2TdRXvwj1WDBJJE0JMPBdfLVZCQ4vt8n/r7iAR0/4M5JPTi3
4mI44vRA9P9fMROieTHalx0B4KThieGjtbiAKpVXF2jCy0Etxe8bSb2MoJG/5faq71ElUCc5WaFb
Km3Iuz7rutWzlvuwy66HiUvgVzXvkb9JmqHrI3qQCSTlo3jAJp+8aah5nILSoeE4kJqfqte99G8X
SFICyahD3Hx3BpLFxTzAGB2HbD7CqXfW14CtvFMrGEdRyPeKZHmQcFC4eUxEMsb4c9h3fELDouXa
VHLUfEYadO1dOnmD6d9Gb3zi+tRD5SiR90C33JsqPh1cUE63wmJE7jgmEp84Nbt+wYRygYqtJTZ2
L+L5OHWRzMpKbrz8cpXjUo7D6Imgi95a37t9pvFmWI2PZX06BK8e4pemTIZ1Jpa9A64aBHSDWnQ1
li1Skb7O3BuiJfUy0TIzhhGXe0sq7z+ZJazgeVdYWd/LWuu5HEaQj5UXpiCOAOzeFMX6htzOly/l
Fc8P85hp6+pzr/VeWsc5Y5CXHSXEqS8ZJ4gP66FqqKtBIDmIVoC/7wTxQVTizwOd8Morf/XxOIU+
KRfd0BkIG6Ihra288hCBkDAHNe6TS0ETmHrpdVQf5UVHYrSCJJLNNOAAwUqS/yryZfOTj7q0Jk7c
1sK8KI56+zUxFvlkbtUwFRvKI93l7n38ai0rGVCWimVEz4uNofS0J6UUMiuRE7yOBYYGAoXYn2VI
GnOd9+Vb9sN7i7vwHtOwuWwZ6SlIXdMCnD9M+1H8Rxmj96mA9lZNVbFGUck23Odlp7V/cu6zVKMp
DvNO+AcwFl0PrvvEoMgbv3jR5ZWhfFeMBnac+ED6LZPqtmXXoM+D4hIKjoRd6EU460Z6kf8MIHse
wDta9roDd2oO0oPadcfcJv/kQMtWsXYd0ivkk4royJtwB2jD04VAooe2bAD2XJhMoA1iUIvngppJ
nzM6cJO35OCcNZA494uFG4GiuaDh6Go6n3oHBsR3gHpq/SGH40+VgeshEWw0/M818kotGdTUH3IO
UNiozO3/VbaQ7mZb+HvTFZ8MFgh8Nr3uhZw8vrBISzx23Co5iU5u+C6Ezk6rYUcLlt81XvM8epVJ
OOrIB8EnMyWH8Zo5G/OlHpbUL2oW2pouNehTKBlQA356tvITnERkrfknBHvXLLJf0eRu0Kywc8VI
a4XzSbqyh1L3svxFYXxLN682JKEUwuHN3epWlO7WNrxnkHE4Gx5U1xb+D0R4zsMpsnkzc124XIEA
cqE3GpCzYWL6uQbn6VEcXEfsL1QrqEbqppE6RDi0HTzkfwZeIa2SPJne1K7bWUm+ZJNNGmu9GaEV
qcW/N0TJqYNwbjdVAbVR8zNEAfTfcXegKe/wpo69xBTsj51HrPOcOjiiNZC3f2FE1Mr2oN9ElNZg
iGA5PZ5wFReqCQL6uKxeC07wMjlZBbezacajqbxyc48Vykql/wTcat4jqkqH3hjU/0tl5BkKfz3Y
kVQUgEAW2B32L0H69baYlZAvUizjILMiJ86oCguLGwreDv++KPNdhiMZitKlmdDiehuTZyds0rHY
Fr7CHlmnOk10x1RQtcpsRIeZvCavxU/Yrb6fcs94cylljtb4L8oBaWdCzm/jOnCbEm+2oF7uMOTx
6fiJmOgz3Eq2E+8SssGR6gecEOlfzMtjlJesxj2jME7RfxC/27qk0mcWFKopu/JMOjjcRX9PGBTH
Dqr9kzd0nzlobS/bmofF+PvC9rXOh2Yod4zV+A5hhzxzZ8WlpF8t6vbmxemympFLT+sGLKEXRsBi
zt0RuWxZPkAMBcaApBVNf0jG8DkWMD33zH6MTjLCg1zObAXHxmDPhz+kWoABGKdJbVbrWN0L8kNJ
wm6DxH1yM5zr6p3Xu+Ggy7BradFz3yBeT/XPtwEbQHCibEOx+HwoyGYptH6hXHeYUjdlcXcUq/Dc
D3v+38P8iIh43/sfNNwl4sHbYuyeY+Dg/X2POlts95+kANqCcRg1r/JzWUcLIst6S3btHN49ByEW
Dwzhr2pttLkVw3isN+Frv775t2RxYgdmbnEVoVQmC7rSD4F73tEScHVoZasqZGKVEd+xBzTX/0is
TIKK1085nfxuQ6VS4sCd2kT0dGgZDNzVyo6c0393euEk/OZiJ+g4aVJJ+zOXXXukacqVeVFJs9YT
DkPZE9JgCozPYeEWj/t3t7UbndWMFgt77YmWZF8OtCq+l68t0bYJF5Jx45FIkxS7+ZTVKVjhlWjt
vWue+2tIX1u9MKbuqQSBgcGrcNmDqUXaQOsjey3SLv+HdY67YAaMtOn7C8clg3Qvb+QYNVdri9au
e1bmvD6BOdpv6+euZk3zpTqCdzPqbzz8DL/GgTZBg8GbFiw7ZIc1MzISzXd50ixRizgRMoLdpiU0
ydkESgfUxt76Gkrl54Kp5GVFwLhOst1unumiuhgAgRN7Sac0okezYTqgEb3hyBGQE8p1zRy1ge+t
pzfnj8NRgzzTUYTgBr1BN6YZChswJLWG9dodXoZp+WLXtp+7KxjdScHinQpY02ywLV+bzsCAaUqM
xIcVcTy//xAU+MMlU3wgVBzul8yGhyjo1Av9Oz8nUSPxEnGz+zPSh40pElJ7yZjT2RId+IuOcDRn
THGkbpPItpWGEz48ruIGLEMce8BIKXhz62wUB5TMDVgoSv9nxso0O70SkKIdTDKsgYPZsh+rxmc9
NpfZQSO9/mtHmzGrJRC4MxlByCa/oVraT1+Yr408W/+yJs6UwJKWouDqPXhLVlRj9491zmquDaxO
y6Wj4YC5MLqJ6k6x+uHxl3zqkBmhfXq/kswR+wGgp4XKqwbVH+NgnMUh3hfeYYPH+4ggpfnxzb5S
pwRjSqqbUVJobDRo0B7XT8hRVeGfSNmTqwL72r19xXqnMwx2CJe6rE8Rq3b1KS2MSSUlCKlM9QcJ
h8mRHVOTKfeKdutM6YISnK9YS8DZCrZegAZ7zuUirWiVriYl4VccbTEeePJCm2b/+oO3GCUdzzf2
ymglt/5v4Jtu0qg8vT4PSzpqko4jpav/46DyF2s+nMsw8w09WOKEJsTAUxA0PxpN6OKs9GKwmYNv
lI/ux4T/z0xR2Zkr2osy6zk+F4EGrebyjsH83oQP7+2tikDDw1uTPl7w5roFSqvATxIuoec1L21A
IDnQH8zvI7/7lFr2gxeoD3BN0vf7ceKwJVmEwy/fPXipPxdp9qnhG4COT3pYf3sc1MlbiRyBMwJQ
n7B76RIjaMPz4i4PwPeq+tRYUYHZxYTY9/BCAZxipttAkmhI4N081tVaovtRwwLYjy6vG6H58BHW
ffGIf5pRln7/ezbKuGCIlmePI/lLvYnAda5DzNffxVqvqFrsSJt1r47dW2JVFj0LZPLEAKbnHOxI
daSbdp4MMQeyRuL1RW5oUoy6aWmPJ/ZQO4T8ag4DGqc+cQifLklmM2fviSjFJuTvkyg1eOScExP8
rzLAvhQxFAXjUvl6RMHY9STPgLVmqUUedvmr7X/8saSeIFd4WYpXDA7Ju70sbUo191D5jwBy9ZB8
9vBmgA2vPjBVtPdcsKJ02fAI1Jx2aimAUrm2IQV8NuDR7rEPIUZEXmzuyB2I7Dj+4OX8yzKqPjZs
aKnLK0EpbXLa+pTOvK+CMxYBPbKqT+tMxdcNJ6JqcYtJjZMi7ldWE+QCGJFQyi6JTKsqrQ+L9uHC
R8Y0NxKZIkUfqBkHkh8qhNxTeq3OmOFVknKlAnjowngEUTFRRiCmnqkMgpmqVX7LNBT39988Dp3p
BDHmoiNTk1N+CO7fYxB83Aggew7vQC4VGINtsIr9sWw7XNfSl7VELcBiqySrltZthKCzQUWeXLAK
ri8zPR+oeUR3oEAS3URVIAvMJNxaNoGvKHXgC+uRlZaBb0f4JqMnvxH9+gWRchxOAmMuAtcIK7oW
Gd9pabyLWRHD5lyK7nTO8jlNsxbjVByhKBwOVVuTBwaoYcKMveeJ1AN/YWzLDr+mdQ89TR+rIzkO
43yC5N68KssXClvA8Qyng9D/H8T89bXF0dDdPUPMVKmiR1+vV1q9O1VsksIeEPrRcSvgKoODP6wE
Ia6T/dyucdW0PhXoDennYAiKDRdOlH6JKk09MPzdP9rGvOdVsIyQ+20KzDAZ9qZ59HKlEy+oYAQi
VaahxfY4uDtZt2eETolgLvXWzoSaAGC4qEVtnWXK8IT3UTRZPVipsmCiTquCBsPYCzX3qM9nQvSO
qMlxZAQrkl41LXTW+gDKhEeQdNsNfSmszoaVeQkRCxLRA7utA1ncFTYoFpFX2Mpf8tLZ6nggGgN0
ABq+X+uXkSC5gNdctSjalu411F5M/vsud3zKW4OeYo9M91zrsX3wR+On4gZy8AbPBHMBVAXAtvVH
2jULKbc0UFCwGbCCNWLzS92PPiM5r6ujMTCpio8AcgrB7nMzmg+QOxPkBTWa/gauJazjsWTYqAZl
Vz4riENlLRS6qQV1t/AZ/Q3oaIZiT/qRuMhqAP1Xwm/apUurw+ktRH5enx0yZ+yHf661vXEK1wVM
pUg5xjuYY79FMEyCusMjtbnOtb63ulYebH9a+vxL0bhzPRmbJ9+l0JUiSsyajhnFF1JJ5GJv0Rwy
TqB1pdi68214JAyC24n6dNWMvJA7sLkj9nYzF6MZ95XMGX52MBkWD7jyTKnSqXv+bpXjA3+gUmU+
vsp8QqbMX5i0oVgHMspR4NZEbwCn0XkCMJXsR1rwhYvlQoGoZjNmT4Y+uv7Ok0d/Q51I9rGteuTS
cDuMjuWWvUQKq1aP3Po1ifhI7k90RAdMuDDnLRwzro4PGph6/APrRXZSvwZAt8+gPQWn1Z5bCftD
BCsJs8OyHk60vGApNErWGTaUnK1RqkcAJlJYmfSNDBheVUEu44iCWnnb49YXtgu6+ovdmIPkt3aD
LNvaC3Vq7ChjaHRBorcVAcH8l1bdSeNuk5sI8Op6eEWEGh4eFAhe0XZQzE/2q3O7tnsfh2MyrSfk
qfvprsKVBJrhBPyTG16m+XnNZdx0zk9nB1//q+npcQGP/iQy3IETcDlPZ3TadMXybYFzz5a4rvXx
zq/QWbpvnSYJcuF6Jlgczzg9RlAwOsCATb9iHCYspinX/N4LgcZEXaZjz5DjJLOT+1HqE/vrvs1Z
jo6Fx7bEXVpH9vILDRkzmnChVfAEJLcVAVP8j18yX+gBvO5Y4VKVqpAfNOEL5qbZwLV4GoiXd+su
H+8eO/znsxZCJEpTkX55MCw2DjTMqQJtG8KdGxzo8Exm9ewAyVkETJdVB9j8GUeAnPdx5d0y3/CO
UI0HPH6EeQ40PrZQiFFP9Z6R2gCeyvo2ToHjjt5ahJ6NW6wtqRNibotkia4H1x5Tujdn5dSzQ+wJ
K3JgIhOkcfDKVT2CWU1uNrdUvEYtou63e5ogH+2B6ay9bc/rnr/RspSlYdWQDkA0PDCVHoAKzKCb
ypBn0k6xwQiU17TMHnrxdgdRXqRIj3QvqzWyO8E99h8dQudA5+rmiPP6hdjQuDh6scaLwZzg6hob
/0aAaTxJ6VR6TfbVctctip4wFIIqxU1vIlsHzR1KsvBAomUWyXycf9atIrvMXpqE/x/uLrx0vpwC
+KZYOekp8stgvMtUO6ShJM3z5Jd2cEM9UlS2Xd93+HLo3Z0BqNH898l+Gs4Y9IgXCUmjwaA05Fi/
RnOWTgcT9jC4a+91k/10VAAWdYCMbu3x/X4ToE/cZQeDpBfjwMeFfi2HqorXGcyelTDitFtv7DkE
NxQJnf5jWu7bjrv8JYpkcmI54xljg+c/mgzCbC/AdyJva/WKG7EaB7NOGm2ZnbTzQsUUvUjtMX/r
D5N6I8Ijx87jlkaHiS+4qZ/DOilM798g0lkXisTPnQcp4I8AkzOxzXljV89sA0dGh2e5BPdaaCNx
qBjBAqgKJs0+8o+6wL9CbIWW7spyxIbGYsizqXAxHFsvgsgSM730nD+lGgSybch0Rx1P/Dzv3XqI
kFVXybpXx0oUGB1uVNK0zDK9k1o1z14mY/Mn8B2LKkmY70U2OsDML2zqQG9FwH4XT5uCj+TEM61w
X0tzepKHl+T1ZbeKmcKCnFYl20SOGj9t2JWiqsPxtHkog8iBf0Z1hc3jHmqPDDhq2lHw9eyCi2gz
lETJWp7xD9h90jm60j39feeEwtp1PLx/PzlDrPty5m21tcFK8F8mDKqw9lBoDIuhT7Jz+nAnzqRN
0WWxBRYf6avwPw7TUzvxbDo4LzidoMOdNvZNh5LGLJxXOQdbWoNZyt8cq2H3VyIYHhBrs9iRbzUf
QTkCMniTxD1+sHB+IkeOnEBy0iG4JUKbUxeQLZX86YKScNjq1P6i1RHZ65PJmSXjrQUINnm2LC1x
EjqojGr2P1hfuHGmOuGi4FnEvFkXHLROYyaZOVeW/Qf/u21Dv2r4cc8jhCzppguovVi74005LNVB
uoT7K6AV8ZEvszmLpI7Xk1M3Li0P06PcyTsTs1CKKEcHLGP+Y7hO6YT+8HGcmGRP3l5kxD3EzroF
llHEOLh0syy8i5SzIM7ABLwiB5+EyXlB+xasPUfCFWdzw6SaRUKn755TVAQ2QOjda8w0DVmGXwlG
xTAkOONGoHx0mESN5XEUtlHo3gtg31uMiRz8MxLMUscS7+KV6J5MO7Mv8eF/9TWUMqMTU4Bi+DPk
OD+hMniabFSwfKqCdK3WTPntU5RZFLZaM1+v14fqWT9uUIe3BIlkX0p/GInMBUECVM4oImzXr3IW
FBNpxvUFBqi2Ket6fhzsTvQZGixDZifHPT14H2Woy/9DRtzd8HrJpd5GSh60sSXW2bubw78px32O
NdeKbkvMTLlRoNXz7zqT/mUTmo7bVghoZo0YAQvtDwbuTD4BmexDsIdPasMDDmJ/Ylr3k9YT8atx
By2Wo0ZNuVpoVoFU3lX7PLzWNUF84GV4Ik6irSAHXmOamsbZMrQt0r0cd1XTb7JLlIRX5uGYO50/
FNsBYAFLkq/gngo1Y3V0gAoYGlsusLoal3zS7NvCBbWakvHZLY+w78j6H4v16qHVxzZ1HNHU09BL
lUJusT7qrb+O84yIgXsKie0rRIPBlu1KeCR6kKwsfYZLL1a4pepFKmpJIUuXIwOPanXPXPHJDQiD
g8Ev14Onz/fQjVDDTscA7s+5RAn9H5sLOJQxxCr08yZjki/RnSkjU6q+CLEY/Pm6zyA0SORaGshN
eGosAbzUsm3OpSu0OF31wb6fPA9Nxbj8gdf7rm9qlfHeS5ZPCCIq7hpUwo3OXjqZCH90gdsGMYiB
eVmlokZyyNZCPYrJSq0OTB8F+5ufyyD+wr4mVRPnbFS9nkUPBrEvhsCCG95oUBLVGOkUPmKpxsFE
dngKeBHszYjH2+ZwRA+LO0Q/Hb06cuE97SmGWR2enTTzDYngaNTHxS1ObO9NIrs8/8Ssp6eK8Pgl
xl9Sgkl6QUr2muL+3jd96kMOwuvUMCGmsucJx8fpKHIKEhqG6O5i9k2h+Pd/Dh6qODWSuI5bi5LF
II0vV+EBMgOv/ceRQJYbdv7cuiiEQjIsFQhZYJIe/ZUON40jPSMpRbiKIZ6y/cAom5oqe/GcWuIh
Zod0/8g8OeANaJaNQrym0LQMpBdyUi08VCHbOkrqeYRLba0avKkeuiDOsP4VqH3QEnrL8hLFdIAJ
1alIMxTngmlsXZrk0jEaYsLN2Re6J9JKh5Au66pOHsEdxc9wdaLfLCwfBVRQYUmUxI4yW8vTAjkI
RM3RGKu2U6MEUMn7JqV7m90MwgfQkzx5t0JZgnrzYqQpqLcW2s8AGBkcuvEizXBe7A1qVJQ+1qpk
7QuLhzX+0sXzQYMl5rLymrkmDsFpCugxuAyCi60Wtp+gN85rJGRyGDy6YKkODN0TUbi2+60NZ6Gc
yq6sp5fsGPz/k8aU+K9+223Wpha0xGBD6+xWvwi6TLtpDU9IBc3R1kd2ymXnK1QWRfaf03g4kKco
sS2hreaKIb9zdsRBiwOfRieK76JUR6IXpRE7QCJ71luqxXeUzn4LjMBSWfzarjuEJHrIa1AOgPnM
qoH6idReuqAbZGpR3hYs7DamThIIfoaOKIYx5+NbA/4shjzy/DA9ANs+7ZGvnnpmNpgPPIY72wMj
6uxolS6NZSDSwNbYPiocYNGN7wiu+4rJvZ0mcTFltRxTrqypoPNYN6th5MTxSxcNOuXepxhNVBWL
SgojcsAeT7y3Ej/lqPiHRDkRc0dQwg8C8QT2FHOHTBAgUS+LoRr+R6MW9Y0F5WD2nP9Aw2tMFQTZ
DVufGbm8G32WUwE1gbVnkiGuLj0mLU2YpqzHI/ENOl6/K8Q0DNl+8vmsoWKsmobjraEIHubV9EtC
nCODfIRQN62B3W/GJPmSPtGBqLjLWoXWWi6ZKuEACwbdT6yoLUxBohdtS/ZShkSWMu4TG8aF8D7P
/w2dJueZvFdok++JVTuYIy1he6nABIyTl9+je8rt8Yjn/pytbapUTgidjGwcoTZxIeOLXV0pktnW
O4ZN6T076Mxbv3fnV4CpGhZNIm1dKCsPESRy5rFzwG+LJZLshuR/a+0y+Cia8IL2NY7rt05vcWiR
rSTYVZANnC50lrpIMSTN6RT4N3GqPCTz1LH5XtdXdGCDcE172sln8aKJQPCAaYgsvDXwhdsdj7fO
TohvVkAys6A/c9VCxX8QrrlT0OhF3Qw+cEBnSOsC24vv1tClarYZ0ILStZMqOHowVQ9Du1BLWQz4
H06zwjqGuwuQrEAwOUhZOuhaaqBp/m0QIOXZ1Z3/sxn3+ZzWnY0LhN/KigqJZenrYuJrnY5BE+1h
VwuKW4xejq9Tm/s2eH0/De9mrBIEoCQC8FVxPa2uhbNCNWqK2OUY6aZqj7Gg9F1ptxLkMC0NQq6E
JFWRtj4R94d21hHVKcz0PpUj2q5vHWJW8C2iVNR5Q8+7qGyh6WKSFy4C1eRAbQ/hOt1kOORpTZVP
CuMC46ETgBjRn5sZMdPuOwH8KDqgwkgnXHmJnv3ff+vvzHulVm+qAdZ4B7uLe7PYIPDH+EawmleD
IuNeHKyxxtcWIZ2xVSprVlaXiXEuQu6nJtaJsqlgFhJ8iMR/xANgL2mIARlIcg0pXpYEBulRaCNB
5EWNBjkJkeCXXKZ9n8S9TPLFfVFRZey568S3R/737gOzXeCoTS681s0/Ji/zbjfpeKtP4rloDOoU
qifW/lbVRX21nLusmwaQYyvJxavdPC8dii0vgqrVpRc03FsS8TV6qtGK4RcmMVaOkRoYyJDcjzb6
FnDvbAZ3/RZqg6dwfR/O+3R3E/ZbJOVrGkFAx14btRdOoSBSNkgBxygDsDUez+KaqMD4hC/MLIpz
r/yAf8Ay6jDRkuNRaOiEfyp1r2xFvgBBNgV3gSG9QDelO2gGSJz6pNCc7f3hvHxBZza+7V1qnm76
6U/GWbD8BTK5KsZ10ZG+mtZI0H1/rMAMapUIpa6GsEdepQbWxqUkCYULtiyyTrgpjct4onOIo9yM
5VWl/ScIvw4xVYKJc+HH+pGOAjhtaKrhCVbVRG4KkiXzUpeAo8kd3ZAkCdbtoAxx6eyFiEPyWrxe
PoFi9CFgNewTR/ug4hTfU5vXD+GMjT+ulBvmQDK67px/WdEFhtcYPyHjNKPKckEmxMYjEDR80RPb
/+FuSkS1dZJHGIJsHJ7T7IX1vjez2qohbZvTIvHYtH9s9ax5nu5WMQS88NJV9zoZOzeN85q2FfFV
DzmOf/CoPSshdc5iObvKebng0HuRi7WSkwF5YXvwYwGJXc9jLKMwDkC25tmn94YA9GQca23PjmEb
2PbprBts585B339vX98evbOiOkgeXetFjPEkkNJ6A5CgdWGMvV3R1yaaN1evqI9nldBfhPplijwD
T8OnbwJvehQQhKOeWqgw+j9Vu0vmJ2RDU08yU3/rCORQSqmWOYEzSyk/FLINif9rJg2BqfQNQce4
J5aZiv5tPNjF3YzBAvFr0P+j3CGMTp0hQXTwtL47v1P1kVxgTEQcYg4JoxUreUG2XIzYAk1RFRRF
sI36TKB/e1qrd5fdfGTWV8W21X/lMD0N8LixetPYiwV2ZQM+Egj5mhCX7cXBUNpwFoa4A8SpDq53
mCLt+S0z0SXzx7M1rwzx1b24l9HP/jIWbrh8zXq3f95kiNl52oFpZ11nqB1LF7/pfRYR8czEA9yT
XqtuQwUec6LdXBp0NPbcs7/R99yfo/jS+GQsM4sHdu+ukT5PZH6S+rFTn6L/gaGInpxjKUPsWP9g
K3M/4//S45bbv/5ZuXg1QOiwhruurNtA0c4yVy5ymWjYnaEOKYxEERCA0FAQPnpA816ZmyKxMF1M
akRMpf+TQ6p9618BczK9gxjYMlATHErwhVIrciJrYu4ibMGyO/k1fCNQ/bJZeWIdrDM3X3YnYQMa
P0H7CjDhNc+dQdVkaaxdRYKQ5nh1tIqrgdBrERfzQUNVoGCRipGJtZ/n44vlrmwSgzm7Q1zM3iC3
VvcCLB/1bXLuQwH/5Nv2emIylKz16pAq3NBrsU8QXxfAENK5bXjgCphkivqzDAmAjiR2phxB9OpA
znEcFH4YxOwAG2XlUOP24YbG9r7qPJMrlM6CwDEJYCikARHqLI4Vhvquu6xH0A3HLYaVR+IAYslp
Gp9wbgzI+ggDuPSHaKoeKieeY2IeNxZgdjWezaVO0PwJD2Cum5oR0+6iGhpIrZmjTTzGaQtRvXek
EZHhXppLcfrK8IdAy4HCUTC8C8BaFNGoVXm0WytJVmudfSSPl7ZEeabDxC8SUKJvFY8jyFj8WSqT
NV6YfLVWbV7KguqhG5FktQfkLr3lCN28r4ER21GBBZi70iTNTuVplI21C84LJDWlXUmVT6vXoqL5
/7fmuoCjpLQ+KCBIVbakXEUcPoAehbdQflhpw9uTb5k43AMZnnpUKOZnx4YoLZhyoW7iusbQv5Xx
x2EbUP+DU2rLOtHW1Gx2WlS/y6zj4AXwn7O4uWAUShz4uW1k+XaOhT9b3LyXLVLIoIBqP5Xe6Qdh
PfYfKO3LrS7fhqR6Lg6/YN15o39jX1kis7o7CqvZGrn/SSjCCE4g6wIg6bajwZ6RqcgLVmwnVFxo
3MxlEBd8aFEg2coaSy8UquD5+G7N736oNVsxvhzvCADKL3Ci+1ylHWe2WJdUVk6FvJd9sEicmrOF
LaEUjn/ys0j0/WuO2+PKOcRaEF0EXUtp1WznYIq41nxJdFagROG1NJ0Vb9xnWm2X/8HIj5h9OedZ
5CnOv6aSsG5AIY53V2so2ShumcFmzo6h5Ulw2H0H2PYYaKwZPC00EMopBYBKns5kykJXB7RKOb9Y
AFwYXGDisBKbGPYXwG0jo0alqEeWPgQdpPlKLELkIUw2CXDWWGxicX5Tdui2DUrNgKevn0/ypGhP
txmOAtUXY9srvM0ITx0pkk0ATqwYHNjOkTsHPEf1dIHfHaL6hmV7K1X2ypujqB7StTVMR7Gkj9oK
4EcXqy+9qOBh+e9TaLMoN+RxDCFEZ0/H+pErp22QjhZl9HqtEhOx8hJpoEMm0NzZkLzzXy8c4U8H
2iTh3dxAzEPAhg8imHZ/zlanccYJZijCDOHac6fB1LJMH9s7hawo0XePQoL4p4kTtUJBprmlotU1
8MkuCyc8wwwQec1u4EuMRL54M9Pp8jye8QSz2nxETpJr3C+d8Xwjt8Be+/gz4fFQbb7E71jY1d6A
QFEp5nnh7mawtdUfFewJtSrXbU1inq79xuTn/ucPsxdWhj2g+UtG0wXgLQ9S7JBAsOaL8PtMt0TF
W8MGoxGTBeCzHU7IAZPTCcWU6n3vHv/S/RtkFSlPl9a9+u8rrlaS9iNiWXBRdQY8JU1tQDrCSw1j
9UuXQcmDP+ASOwLXJWr5gnuzHUO8bGZaiNSEfw5Zn2ITQE9H9Vw3iaDYz9LVzwnrfcQ1dQNe+YQv
xXHD4afUGACCTM2hJroxCX2BFgE+h6Cw5YalMtYIULq3xHNoJyDusSAZeqhBE/kJZ4VOheyc9KBy
16rK3my2/QrjbEdPg3t0cIfwm3W6cIhwLO+jVHhl2YGmP4awq41SLc3dLl2Gi2EehwneyvB8LmDQ
tn3MQGB8Tfp1vr0AfxmpJ0OMbNJ6wVO9Hb/1I/Sgef8mSvQwiYVmt7zCGaGvvUzQ4iYZm74cbuSg
26izgzODWlPqn3kuM8sHqELtXpnYwQvsv5Yoi5bn3zpuFlkIY5I/f2na+WIic/igk87oerKZLNXx
Cm+VqNbLn+EPqCa84V+bbRXoOMtQh8MW5iAl3XF4c0ps1s60158opRy46E/d+Eo7rfrCQmAz83FN
ERXgjcP+yR+WnjgDhy/CdRi9eZVcFWSS2baiB4WWS/3koulAxYSc4XYgvEaOpEGNmebhDJ/JfR7W
F4Vq7y/JjpMm2yXjn4NxgjL7mWLmgXUMH6eWCxUrqq33pn1qCC9EoFykzuHA8TqAYMt5s8JTlDes
vMgn2tOb3vIrG+63hPQOBkm5vyHM3zG1lpv5TaQnk/0tYcToO3CbaykNVt47u3Nx14g3UciPoZA8
v3m/MdvlLfz8XlXgt49nEtYRxs2ClK0QLFGij/df5RDMRvH2ZQOun6siNPr6BnqMrWDQ8UcGIbRa
1CzAX4ShZ2Nq7StxZrlfC2Ez2vPnM+t6bJvWCc9ILb8lFj5znu+KlObh+3iEJY4g5YMfehW8xNXg
rexv4JzsRjZNhcv2FeF+aecfO2Vy4ieWcy4V9ONyt8Pw3yJjvFi7eraukJnn7Ynvod6IFEUdyD8a
hXl4au69vZM6+agpNws8NvTcNrKBiTaxLDt3Ehj4V2SK7A1mRdCU5lfE2NyOxmTZy2rXHtH1OtlH
rn3iFjSpAUBqAjnBOCSNKrTe+A+de+XwYbA2AkJHpAYRDjpWfdKdqsDwJTibu0HFFmiEtxcVOlQG
IRe9bhJtVHxE4Bt8hMwiBLSthfO3f8nx9xFGojrazSLX/Z2ewnk30faiAVzRBnMcBse4NcMJe+zk
mAlCtnVhPTKjuZbnKuX8Eu3LO3sIyQg7ynW10r6akEPpvAI+VEU0yeIDoO97GkFIgO+6bt+pJ22t
in64M6vgt491ZLXOGmQAgDuKlbQ82EW+ZXmWMHN51rGxjjLJOA0bqc7ELAWoz6n8O0nQyqEv8Zsx
UirP7elW7rN+eaDY0IFk0ITRtJcdPyGn1IEx9v6BViVxk0lF/1ls3wS36NiZSGtaazM8/9+uj4kX
/BD9jyklm99qzbWC/B9MHXZSpW+lzEOYeIhtz3wWgm+jw0+isG1za242hS6YZOhxpBfuKWElZrGM
Z9ShMDm0ZHiMagvbC42MVyQGHtHIaxdwxFv4DSkGJrKzfzHUkBQsPbVAGRh2H5WzmHErC1NkUxUp
pMeDZGTerrd91sdU79mZxfGJ6fO6d3Y/ur82OKRxThs1IC/xYpCjDY98ZEvkMQRE5XwUqhnGESi+
mOwB8qlcEi64KcYnuZ6yFLN1kQSu4MTrveT1nNkpH7FqmPu3vHL88zLSO1zGYxaHf+winh1I+KvR
NA+FbOumwHzYhds26GeWDFbrzMJ+8D3s4L6kOsTDBY/LNs5dQmIQ/O6/kxilLZk4tkkWyVrwsPBI
5Vzsdtx04z55nvZuPoJHmY+NcPtpne2bvLFGf/BBlii1qsLqGcbR40pDDUiAv1ikfhrG1q8jDInE
leePHXRYTQnYO5qfyBL+XiVxsvDq94r4wnbz4J0cUlFSnT0FOB3BbldYngjGjr/3avGNx2azWCUi
GDb6AtdpPsZh/7hcd02LzMU9DOSdseoUtH36QOwGy8T4DgE/LA0BaZzq2FNK/VjW8Wtibv5hkVjn
1nF0UiBXz6hJVjCs2tFLcv2X2uKxd1eA59uUqcEMy/+QhFguyruyGS8MR30wLuwUCdp2OeBK9VB4
y0PfoUfcWOXwlM5gCAui0l0OuW5F/NZnK62eKPdv9WGxezf263qYbTCnAtdmIad4G31Xakopy+/A
TcPTgyNpRlzRvZAXfUzvFfRZSSqEuj9o8LwXgvt4Cc1N/Z2Jsnfgsec+IBm3Xp+jDTN04WjTKWkt
ixetNCNOYsELCqdcvGbOymiBHEsIRDuPMsXzJO6b3Qjqt+N3xQ3NqL62SzNNiVk9n3u6dOiTexvp
Bkd2mXnMnRKXPS2yLR4bNazY8CvndzSTXlmBI9RERlhp0dza9VX8WwTKygFaEfLYuQZRLN89OtlY
PI9bPK8uML7sCyKqzg2cdvMYqTx4oXtcLhr5ZCxPVfF8UKB6lIuuy59jypxpkrh9ZTSwM37UpWHM
lODLwP5g3hgAc+UKgCPqhpOvsJpNVPmIYtB0eFi9Lwmh2jdLHxCM8X6MDKhsMhiIFdvxZvMy8CP5
o7ZvvAwHcFKnP0cny1GKhw8/YrTLYvOilPqA4BWHqGkveIpvSQgGk937eCWIlhIq7loJvzrs82VO
3j4+bUsSe2JSKoQeqNjGmrvkkyKiciJmiQMuRN8SjoLUkc2RyQK9JUNg+ZlVN2krJItJ1u8ZSr+i
SQDbVxxuqY4vZ0BDczzkaS5SVJQojPyP6z1ySJLYRGnaWX13+aRPe4+uUsRwwHsrimOOPeA6lqtQ
9J6+/uu3d5CgpL/ai/1jDzZO9cHswqulPxm43owS15IOPkIXGIiXusDB/UKhAeVdqFvl0mzC+Qd9
GwBIWvENq6H/A9HXd0AZRCxfijGo7Y7zIVBbfMaMM3B4DTSqTsM2gKudLyisa5G1UXSJg8CrpVxY
o0IREvy31ss1NRgRSiiB/nKejrACG/zTBNixCy0GOhgPaJTGHBJeZfc6OCkJjNQg/YNaznv3Oxjg
sGrRbZM8pgy2Z0Fn6PTvZoxKLMhTioK1rjV7/UGcMItGTM24m6As5OxR47SFCvz1QRFsCs4X4PdT
FJQTc8nGjmnQCd8uqnijOPF7tSMzCKZl+6zJbKRIJ6BUtxD6ShVF0ylEoa35l9L+RH8V/mXcXp12
eeMNk2JF+j3TqruIJDoosZVRK/Vr7bJxhNb/zFQBNEkKfg1rrxexOlPjDQ5btC/dkNFPBvGr7oIr
hGns9RnB87HAQfcnNnNGZMicMfe0tK+Tz2SOOBvhSlnmQa6rFimwOwpktuVis4L+eF/Xw5D+Lgwf
BvaPCxoFVZ+g+I4hy0qd5780KucJADSRSB1HbSUo0cTJxJI+5d7SIsVYPMSrNPbtDoz+LRT2398u
E0zWk1AWi9r2XLuyTFd7328NhT+v2GViao76+XTaZNXrxtEctNmaMzVMXPzDsQWm+dpPRnsNxogm
6OdN1Xt5iLtVM2vB9KlJVNkcMbkLdkLm0xPMbIPTSfsWP6XmhuQTz4iZIliI3HVhvO4eOiWfqhvy
yVbKli+pvrpqdR62Z/HG1Qbmt+DSQNRUTfRakteSc0p0BFIhVihUI5BTw9UY/09agt9nI3EluFUv
a9F2hPvOsUBlu4jYYBVYI49iQUsLfZFTJfv9DMyaCsFv4GSpIM/b0S81VeLV9FULACMD+Zi0/vn0
AmAN9+36KCkb/iwHmrzNr/RIvJ3630OjbIRPKL6JfYvJzmtWfw/+vYpOtKX1Xak3dS8btQzFllkq
T+DvHMfC5+0e41zBp7pAf7R+ohk0hHW2fcCI1iRkOk/PnSq86sAAOBXd7YAmKXD0oDkL0DzURWVF
PazlFaNnhSFyooqoobkMjyI5ztD3t77YcL+EL+qAEb8m4UMtlMvs01Zcgiay55RniHfFK2VOoijZ
lkR1yo40CFEJ78eBu2XJHqHgU0raOfMn0ZxPB+N7wrI68wLW8KrrPtbLZYLmIdPBlQvslqi29hvy
b8HNMoHhc0iCQxiC4GXEstDS27ptGfPwg9cnLrWTiL6RyBm/bwCZ69mcQJTS3TNo77Nz84BsI8cL
/xajf4kucVG+wtdqQxWS4KVKcVFcq27zq9itW0D5Z7zxtRIBOheABAsGsw9Vg1sSmc4DX0ClRHKL
5QExO2qn73OLtLxO7vVcAleZVhfRExgV0Jvwl5itgB4fEg4zfn2vF8/bkWN67WljybrFe2/pKIAO
sjhTjRcDTdy0Vs0phZr4ORtBrKt27PtGtwgWHITgu8OJQOB/UBVlc0UkMz0aVN9dGbjjZLPCEAyn
3CIZs8KJK+Hs8B/aqXO+QInNRXrPjCUaJdkJkw0197qc7oRwm0wn63VHwlMogCIDi97EaMTPwOYZ
MTugKMrAi66QL5ENq5vTDSdzBtl9+QsRFcKNrXoB5Mc+lVAbQ+z+py9Cxeg+OZCcGClDJFpk8K++
Y+N2p+IBHALagZetmL2l0TgfhP5XNPu3FhDlmXp5sIY5AAu3mevPC8syKsqILZ0D8Nt6jyayn4gB
bcGOznYuLkbq6LyPSqn+erBLMu26dEaqJk4wdunV64Ll+20jzAXOh7kYEjxAkmiA7DyP9VmbtYDy
stmr8wcMo9aeLVhDIQiBO0nKSOWjuw7wBCyr+HimkMRrCNH+UXKzjkd8ygV4lW2OR55v2ylB2iZ3
BfQ++Ynr/Y+8Pv/Jz7CRirDdGpjJCLXMGXk64VdiVpa211hgRY4tg0XZYq0awf2q/P5ItREHAr/U
Qyz/LDamVP7oc1czs5/LEnmYFATaxiaFqF7PK9W4lH9DXyGxVNymGab74IFqFPXE0GUy9ZdVIhXf
aDTRxYYe15dTPULMaKg4pJltG+qGFq6FgCC4xtapyVAMLkrAQHsJLyjOyxlX4Vn8uTFMz0EbpQB/
aupOFv5yNc3lYwxqiq4k48feS8ZBgUpJZeFerWJpkZ49BygfLpORUSiRWovA/uvptSzQ8OgH6j1t
oacepbe22DjbtPGN5/fViXA6xh2UXxzMrs3QT+3g29JGX5TUDrFGo9ei0XDSp76MwlKZRFkxbEzh
L0NNmEuKQETNBa+OalLYta2Nu2/ohdx9ltwQawr0dYrG8kFHMjJORebFej7+uS63vjJoYENjfvM5
eQ15JCFY3qmPVnBHh1QFqV+mLD3r24xYeg1kmS5Pd/R62FC8Akq0f3IcjKEoTV9SiKvdToVsstud
Gi1M608gyjyrxMVJO2sNCSrnBs1+l6exYJC/pHrEQmOxxN1IWJAFK+wO+VakKF5B56eq2KL3cF/J
9YeoucK8MExQEtt3cgWGUfegt/zdAAt5OQTVz6eW5r52bdfdpPuPBhfg7RmJ0C+Y0GEf1zYZAR/d
i3tpgMJBei4fD/nC14pEXkDFHI3yRmdBx+WRPplPbJx0MbxCXsim3AUvBAmP+QulVWQC8oEcgFHl
Zup0KkTTNP5X5TZzB7raTkkdMQrhYRY1kNu5lgZxcV6nF+k8TmMp2W9lKP5Y/CNCgLU1IVzrk1os
VTFaNJS9tAr5vHwcsLTaNyBz7h3IzW9tju3UnqcocFmEtYpImh6z5uehEZv8braztX/6i2VfbNVC
nMG+PZ7G+nLjT2QJGXuLoyMsjWiC/xnP4g0N6lqpgz+MPguxVTPpYXaziIklqCG7020dstnVcmlM
MssOKVGk+emHonYqB5dU88mTAfrqHkEum95Vhkb0bHjLuUAzuHwyquSnXb6Ca5/fe6LdQhv0/tdD
p6y16zCmkvI/mM+uqfkcb/KWCvfIqQx7JTSFT0qiG/YFs/Ho1PVHrVD35+zgGc3zSNzacQHX7mn3
MJgjEWdSdn/QZ4zz6HhEdcBWmPrItDmcyUj/7Xs2ukAwKYGp8LgBHJ3w2Tv8bpFyLVude19169km
+fO/LVmdT+WgZb4flmkXdBFRap6+4bAvZqth9knLJYsmCwq9GHc33NeD9RMQrQybemBPQ6jlR6s2
yVnE2+AseK6/LMSo3vggJoPY+A1C2Mzi3Fwix+w7v9UCqcMkuMJPmhMLeI0U/+Y6ghIOPsChJfhq
VhI93F5j7s/DOlDjr9lDS3uEuMk7/+4JFdD7zdnlLf2yOuU537HVC4m7wieeLugZsRePnWc6o1m5
WgrsTmq3dITDUeyJfiAcfwI9/h4wqQx3Xz/TfQgfNkZVByYt51z7CwRRqaiicF16M+qItCjO5VN1
jQkPBqVYTJdnkYowFxSuHQGhDy3ggi4xfXqJEpr1cdDFw1JmbeKlxby2stTsI51JbRv8Ia7GjNsy
zt7WkXL+6FiKBsHbgitiK64kF7Uy6QKinhnkpspIxI2nxcqWaqGJ/A9YmiuyG993xpUWMtnQbo6X
8i7j6xDJOWuxQgEsk66FWkEeKCm2JlXYjQBuQWCMCQ5A1YgzQlNcgCv91SQZqZr3oDwdsNyrG9Jz
Ja+yhHst4+Ua90cyDc5sky+6Txb0AepcJu3Ekf4Q5B9yNFSqwc8cxHy++VL92T0+xakPPW50KQr/
PnsVpPcB4TdruPuO4jruFAhCqqLXVXttwT519qf1aI7MaFkzTH0drLSTTC1ihLiWDB2RBRLnLr9d
FmoOVf7rg/QoW9MpnNPcUHS3NLJKZgnGYFmqjksALc9hDOv3XoQVu4GEk3cW6FkOf5TiWYmmYDqR
O7ex2SxA1MtHDnkZu3z4t39+SOEfcXSRMQA7IpJCNrKB5gVg69VoWUxal7U2A/Dye+snSbBPl/FP
lFfM7OQSB1/lh9anuOxgt8RlMWKGSlrSO4mw/RYV+SxTHcA/FAGQBjO7M6oCYxoBzAfHgDrwOgPb
rFYfw+GTffKGuDmIe6D0CDaAu8bCbE8cMF3DAJtb9dGEeh/xdDmfk4trNJu11fhvxhc1T/YkxzMt
3PIS6ed3ue2fkrBSnEjmzkBWFncGIr8Vfig1q/ZroPJUgLNMyVWKr1VRDQKbSYRM2me6OuERdujH
yK9Zj+z6NHptkQlQWatFxHNAeb+zXeYGF45uhWRIgluJc78qNNOLCS479qqTi1nqZrJW/GlIFDa7
Y8pzwaFifDMRNtMQtC1GnHI0/HoKSGg8LwCgcQCbcxvSb8f7xsgDkPjza1+lDcEfYJNVCLC04WPo
/5N83zpv3qh+KCEuiVvvGTvZyEk362nvm2Ed2yRLL+cLTDAsrUuC3pZWx3XqxvjKXP8uLxCrTg1E
6TlfEVzXMKlISLvKMlIRjPK3EdKoWIxA3DQID2ppddyKzIwCQFUZcCCuvBasS6k51D+DpL9aZS78
ZKzgOLql41i4LJCzX0W7I/ftTcyUm9fW3U10cAn2cKmR1+sx7yLqev25O3d8tHF1Sn2hAB9CEobi
ZECTR0qaVxlCpYJBBpvUOyiGzwrmq/KLIXb+fetZbmLiF0lFRd17XrcmCbnJgh3Z3PECyDo80nnr
dP6rvx+3UtYaH38d3vxNktLq3ItAvc7OivkQsGRyG0VKw/9fUZwyn+og2/RoKU5v59uaQJa/W28E
aXTSYJIsbg4y8V37k8zOytuh58W00FcYqcyotitr1EMa57nN0mWxdmNUDHXPO63R/YHgrR3khxTw
V0Glbk+A69NZZ9xpgbQKlzgS+r7Ph2qQF/YwHaGd1DwF/HPcLtI8e3Bpl8t/Ox8RULjWFMiNFoJl
42AdNJyN+oL51hXfIq8e+xqGIu/1i46dHl9UQCl6pVF0MUCu1jfml4RhQPfpXIk30JSaHG55filg
suJKgyyeaMl9Je/Y7Mfp9ducbiVAi3I6KeWG+YDyQjWKNfvyS0LlZ8ptQqMl38WlOlKJFKokUH4u
loCAaZ/HTh2/Um+Zd0B65XZdqJJXyrtllMifDV38Nxz/dWHaBJLWGT3zTKJrPMvczOPCMaLFsWWo
mrjGPVZykD+f3RsckkblwDWb3UlXczPwZB4v6ZfPyxawjQAMooI2/aE6yrxUe9ynp20UMAu0+4Fm
ey6lFaNzvSjrYyogymtTfxWk+goshXhq3NZ99PWWgRHvBRw0f2ufXcvv+mLZoAVSE3LsQQjY5HQi
cssuXi5iVfTiUctKVZZo/QijuRVBH8HziBNh4adYI5NztK7G00HGFvrCXMaghTAneRCMi1pPeppJ
DTLzqMDcSxJy9lJsvopgkXtPFQWEoESvduFvMNw6x7klEA1iDkWYMlJuC7rOBJqZ2+CEEPgiG1ZY
Wjt5gwTpCXHrYxuI5MrhDm9ktpEZ2/sHW7r00tIgfW+VhPEfiprQR7+bCXg80bJQvirS7hatAYmS
zZeiFQoNg2ffKir0wJoRAw/oupMGqOTs+8i0LzC3+0PlnWvmU+scY1AyRD0aOflYOHj4xmOaZGui
2mVuyIZvsKPZ/UT39XdkLS5NaMrmwhBtdVXJG9q3pRMLekku76Ep3CN/gcJZNhUP2iDQQ1YTrWTJ
r6HYfZHR1kB+iP8lmj1fL8aQKVz4KLXDevVBlhfiH4HDhmm5xvKOPH/QIafGVETI5IRndbb0AY5w
QocENj1uGAtHHFyvpeyT3MAxqB8hrsCOTMMJXcklHmlNjHD7OsitAzHEaKOXuf6NxD1ywCdn4rNf
ABIO6qifMNcAj58OPWgLiDnY3dyY2KU4SUOxOWOdQgrMM5RjO0oSamJXZeVW1mM4swHJM5Tpy3Wq
yOTPFEujHOK9S+i34/jV4kag8P9ts9Ii4oRYcNaT63ZMkctV0Q98Vri9E3YNXUIMG+eqCQHpAtfd
8jgP6YXk0ogohVPAESp5RoenmvHFJLezeCCiaxf2dpLnuj4xVzUCAsJpcio0kUutx/5Sw9aGFLGa
UDEVtqxBSFGiw9x4i8xYhf68Ok1nwisfwyhhKvAvvxg6o1XN485nikeMwUEOBthlc7XpJ7kiVz43
K4k+65OdAvYnJv4hgLYMFI0PykFrrJj5AeH34+7b/OAuf/zSI1hmqTaTm0cJuWj6AzuE1qaBNdbt
sLZOC9gISomxuOcauLrAksVt+smIGmUPqPKBo3BNFKCRS8OVrRq5sdVUcuLc5+0QItNn/LwG7ZhA
QJrniQDdbFYpJp/y/WG2PxkRmW9Sxpgf61Eiz3vjjVNDaJFAOiZKOPLqVzs41Kbyuc0tNakTOQdq
CMkkm6gkNq3LGKD0nffirvwpDt5FioAuJtQHJd4NaOtXdRA8K7r8vILpK+RdJXQ5EVslLJuCn+OU
4+ruk+uSZ7c9I434Y3U52uMbxa126yz7XttNE8KPGqoVwUq/afQPbDngfY5CH+8BBfWsyK88Hau5
wZPCgPffdZ4TWpQDAy2UbH4HsYo4+hjPU1orQBkgzGuS7Bc0Q4cE5uh6zpQRa4vv5vep7EETkOvq
bGQOC15pkv1tphOPfEbmz+yUfjDYJ9mVLaWQf9cFrJNk0N4NzVXt99a+LAlpjkjHfQhsEU6xgFuW
KsNiYei4SoBf3S1tvA3l4fp0y1jQEQLsUCUbvDHKtUcTVHSlKJ92oSQW2ohvBRNOySn6nRjOlgzs
hzCDEQ98msTKDzPRQjKJr2bCJBSTVmGd5BqEIS63RbJ+WPz/XfiZsLIR5hXeuaoDhyNXwLcCnWP8
6QguId3um8BPPdgdA6r48STe+DqJ0YMx+pXtL5yaq7CR2Ig/c1/hqoO2tuGfSwRzub4H0b3VhfgG
TctoEOkCOoHCUkGzorUuO+uYOt3Jw//2EZbOva+Cyx/NmpU/b//mhbVRMeRw2+lAy1rOtRjrtYwQ
7hi3r/CkP1xeqkyky4U78eKnohYiohY/CvTZiGkJ7kvy8nugUKK6cTeFFrY+5L4YttIugTSNNHAe
pn216YvGCY+sdRiaTRZayzQhGi7CALGm23yyoBVm1DZZXMEFzTdiJ4iBYR2df7WrAPu7rcDbxRQT
cG+GqZkiyevuRY6gDF15SjWvU0z2MO9F9nQ+fmccui1Pg8CcMXJ/frTAScTG6bzvQGR+J9l8Rps0
ofeAhbAWXs9gcxLxy0FQzWWcXJ79uQRfEB/KmNBIklSs1Hmww5GcEQGRAaXKhK/wEf4D/TZxvRXr
V8ulD/7PhYigpSkNRbPDbYBD/BXLWKnyUF3OW7jsyZzq0D3wNIzzjzaAZ5sSaEDKbm5MCFOJLSl5
ATAxXR9opZk0GlWFooGQ2DY2uDG3HUXoZJeXBtL47q6kgHnKibnhIYgeysToAuPUP9PbUZzYjpxv
CSp04aHV7ccrY1VaWZWrZL3nytGDXR0/FYTXj8rkfz6CJ5MW8OYRTcMAiN8hu29WX7gm3DFbawFS
Um6QksnJp99PoFRportdMc4oHHebD8oWTn2I9ypxN+uOCU4YsBhVh3RJh4bNhbZHtPk8Pjc5X62l
xRDeBrOkTNNvrSkK/R+yOIm6ozR/lDmUbjeFRr5ybgdntCcw5oNpV4tJ6i8FlLl+ZGoAykkmcneL
D2GCLvYIN1UI7TdOyLR371TECJh7N8q0Qi8iUX8XVeUIcJJrEDnL5KacmmWwWME57pkwU3fk5XEX
sHjny/jpsOeeurTvZL7iohvxUpbkXF3P1A0MhA4rCY5sf9pPxJMar699lYfVKHZpaQq8lxzgqCUs
yOIc6LnkqF5VIXfAHdOXKNay1E6u2duWO3cmxpvPXdjuPxZFfYShVAX2axRD0nhxZpskIEEe37aM
KG8bMhxZH9Q1tLg5nPZQjKnTdauApsJvR7Khb4zu81ufJnGVnAh+4VSsSiCT6AMya7ezNhUEFUIT
Sx9jYhJZAi8IFwH5hD6iPNpgUT7V/b6St9IwCaJPHfbS6CDhuXVk2hgCQvSmuDRI/SApvP0niNio
qzojM4+G13H7OZyQqOvPnsDS+bsgYClI4qMdmMtipwAqXZr8ulJPVHoEB8pCVj2No/6vanOyhg2C
dlXYkv9MvCuZpOZQf/+6vSvOz3IFLf5dWF2zcciTcGAAPuGcSBZMAJpsHqEVyihVvAtHXqvY84UU
5CSyqF8rr1Y/HM8RQE9t6PEMc77WYbQBzL7EM6lZ4gE6m9z9thJ4UVinYkI8b6oshH/NIkBINL99
B7W+GV8gSQUHOnpfhLri+m48EOFGyAuhxir9earE+Um+AaChDKLxaAWgonPEChYjvj7gqtbVNFTO
AIgco9eAOsRVI0pa95V0fnD8yRj3a2I5P0swe0XsstP3zepOiIRHhT/gpcNBGYR9kAPR2IH0Fei8
FVN4tKWGlKxR0h7A2/h1zqLKCQEEt6rXaczg714YiWtUDG7wQ42JQbRT+bN6n+6BaluyNPgNyOfW
Owyc1MWijy3+rRE65qD5NpbMQ9+TiR6xbn3Ybql8dvaPKejdjcUfmVvMpd9RoxV7HFLWj+WSWbfs
/+CSDvuvB8LoIFJC5ZGtcsXpBz3fT5fzm8BgO7Wo4x513J484V+xRMWmMRW6EmXgjB3v+3vmfz+k
X9InKQ2trVLZipJu3tPla7fvA+6bE0j5+FWvMFj8YUNzSXeB91gEGTFE7LzctKrZ5Pzm67OizlQK
eZzxo92xP0YoXlrRI0XGZaw/JzmHdPuw4YMTCvuXNJPSULO78uoEVY/ffw+Kh37zii0U9BKyDzLl
wtH2NxyJn53rx5GPhV4guVvzdYN9ri3HCFaTWvbt/qP9YInk3Xg7dyHHZhllUf1sil14eq/QjE82
Tf7UBihxP/vKjLPBAr0qjJtP5Bp9WElGeSZ9R/IKHGEo5zCNKaHWO+E5F4w1+QCQ6MjkXyG3OqE4
YBh2RCEmXQBHdvjwTu1nHf4ln08zXoYu9vaIbpBOanBgZqJZzF3Dg5LeScv9srn9zxV5jbm5dmra
MY9UDhL/QnlC3gv11XojShi3WjrCe6VHu8vNe78zoQ/IYMfibERBiiiNQpoQKDcZ6FY6LkvbwDtp
0KARbHCdfwqMCQuXXVbJPcQIIrrQGOVv49BCZECyJR/Tstofe46D5OMa7lK49Wx9Q/0vh2kF6lMb
zQ1tHdod5AgCMaq+LNoR2I8o/NrIT/qPQ+YXy59imC78x+TjbHNprHaxuuQqiHgZEPcY5RHHi/Us
bGtw0Tb3IgE5Xfb7YOfdWQwWOvJindPhLj5RHz691kHiWg0FpOWWdzPvDuf808l8oCyJ8hq26+hX
pRIIiH5+nAk8eZnjY35agQpuzTAujzTBg2I71LLyOmEpsk2tj9TiMAS+7Tt21eAGKf/ZOlBrkH8z
/hrs+RzHPQQ4o+bWEeO5tbAVhtBNFd6DwCfG8l9cZ2+pSUv5g4cf+Piy4MI5KYR99Jr7BxYqMTGg
cp+i14Ns4cCIZ6aIHJVhxl7/58kQQoFL2dqDBkq2F61BxWNdBkfBkKfeA4XNpEVMKS/4sI3ofjk6
MnvzV43heSNCJbSlgvGuT2wtID6vkGx1dZFBNOyRUNOVKRFOrMxzN4DePqd3Ijqim5vVLsZsqr4p
j+vz98uK5hxZ8tc8wFc/I2yEdMT2fs4U9PZC3LlQpD7U5SfI3ShlJFIkQknxV6qq7kU8hk6ZipYk
U9PXapjfk/eLdxywPRGhL/oVpcmwl1VSfRGRVmOH3YjfF6/de16xd6tf9s593ad9urVD2gyNTzNt
xhb8DsFsVQFIXC8/Cj/PAZa/wRI9csIg9+ZsuhGlB620N8MBmRbkzy/q49XrQ4OBrwtS7JFKJgAF
f0Gpipjbg0rDUVJD29vkzXNiXOg33211AujnGbgCsF/ynAlclgx7KzUMevvmjt2Vr7KqQzltsMDl
D3XEpdHOrR4tXikF4bxw7Mmi24hfpaavxZd8W3YYc5YfxyXzg5JNlBYBazz3SFcGhx0wNMv/nlXU
1/Nyhn5Z4Dx+QtsRzbyT17s04ylXJj5T1xIkHzienNx0R4/R833nPwl1DlfuTa7biS6VIkiBk2J7
qfM7FttfAxQBgU4Fq91goyM5Ds7wAcCl3w0t+wHA3RnL8VUhD+ePZ1w15th3uDnczK9WfSM+Hudt
bL1/V/xKVLjw95s+vzj2veFpLvqBp1TdXYFtlCQ5ApN9mKnc8snbzYdasN6TG0UtzQLm2Ra4YKxg
bui56K6NsCXghd8IW/RLDWvGi2mG+XT8jYbOLqpoteUEr0iNrUPFtcW/19pnGj/qqiMCXfUihPLL
gSRL64efwDkN6CB7VxSQjdUkblxDWZaKXvsh5enCGY/DgoBavZv36uzSqD/RhRYJA6b7yPpqa+bc
hy6Y2HvqVwsON1eeq1zvpyD5NEKNso9dz1RGb1P6orss7oUhLhwP60KpZQbS9cFndC/6BpTLxNWz
h60Ihw/vuLW5+V4KYXhEb80xeSCH47f172oFz0EJy3iC7D7kPe1Pxz1E8/K6MUgH0Ead8IyrdDrm
lPPlydd7PyZmz/0h5yQ+oBTqnU1SLQKPtkL10QVc9Lk/eqSzy9eLSe62iw1FMk2er+MgpI7e7dRh
KlWfham1C4Q6cfK4Q/raeT37RL5iF6Ze3fxZp1Zmrw+d+sk7rqhwkEYKoBioFNaGBnpI9OLzJGq3
mOgEhuHC2kTI9lQasSge+oWW1hYdsOpPhXOOuPntjQbty2OKlfaO7qBC2xYu7PTTCsJ4BdM7xehb
2ffuuHJLCBQdlpI303pZALzU+tI1ayqEaxMaa15OliMFDhTYDVnl58uioKFeqYmro3rwZtIfoUA/
pB56ImPwHgvowsKls8CYkK3W6G9qKmm+1KdIFi0PAt8dOo7SiJd7woePYaGdRG4CxhHw2A09uIZx
tr+W65ZsF1BJiABHslq5qQSeB4cBM/lcT4NwHPNyj4nOQr0sX32j0wgP2LH2bol4fp5WXl/55xaY
uPwm6hWkIlAOm2PTu1L+uTGQ+anJ7sKHZnecXAwG6+oJNphayhEyYTAfkEbo0VzSWhUSJYukcBN6
sWdwKwDe924l1B0nHhwxAA0131ZYj6Kv2CsABRHUUS7mTuNOYWkyovrAC7JSgJR0MrrVsWH2obHe
DrvO80OyOS97mshvzQANEf9O61mCoNulMq0fAJ3PUuc7QpCjkBzi65TSq2w4OPUEy3eOowwlYoXu
6e0tcwHKu50xdR4OyqSlXbFTNdvlzUzZuk82FrvqdM5RPsRQtRpyX7b3RaokpnYGergUrMUJTnJd
Nz0zpebtP98jpG/JJlhSSPKb8vc1WyZjvuJLAN+EnsSYM5uxcaJ895cN2B/KEie6Da7qb/ZjLC1f
cS3wTxwzDrA3dmWtk4FArmk0jKnH+0hKWjZQznEjxadWGpEjFMoKYSFDhm6M8jgPIYteu6N5wGq4
dfSR08dWk0Hi1NOyIZFoXKIFv9mabXxXmPGywCWSGolXXB9TtbqCyDDelMtj4BvsvxxaMAdO0+M/
cwcpYDxaOM5TXL0CRFNvICHmkuGWzUK78jI6Ch5e/6G4+oJzNkE0r/tlUzp4nqFaYYE/Str0I7Um
V6uXsRQFSFPTC3c59RQB6bpggPoxq9Z/kfvewPUMV6ACvy2dp7G61JMUQ3aP96y2Yi8kTVajTqFc
QKqLKuPCvm9qZNTekmHczVsX6nbROhIpVHFzAyyhew4JWrBYANxzpN9K+/goi0ZVvBPpM1gRQ/JH
JT/iBAzgDiM23aV6+A3Rs2X7BuS/xfXPqqQIfAsyOW7PtqXCws5CPfiAQgHFvTpKH2Ma05MSuYRu
6GTLY+V5E6Wnwem6esWp9nUjaqMavQAJm7PImmexxUQBIxEZViLJ3ARNELztGLvzspI6dXPKl7h4
WwRxVbnGzAPB2RtSzPxM8PLij/ygs31QlGAiREo4IWH/y2/N8x7+YvD/dW7hKM9D6oPWUVGjLcNq
2i60Lp6JklfwfbXvQvScjhcthWlsbnP6n3f4KnydgVuMfwdA67ERcy8/OatuoQvwu3vBBGBRuQnz
ldW6wVF/GTlX4GkUKdSwQgBIFsjH1j3jyayduK2jRVzQMGdrTamQ1CxNUIbb3LV8y2wjYT05CNep
alQEtRK0H25JKb54L4DfxE9mCtigkcj9hi+lc0GeRCsmvMPM121fFDAs4gj4d97M6jsDuzk05pww
5GGmK9Y9PAlzL5anfPpGJ5T2Tk2DmZM3ZzDh7tba/xty1PjmUOBiGdFZJVsahA5s7LnTFk/b7UAO
NcsSMYVNyC0LAn5eMGL4wMhssuwG7q8piIu5EY/rk2IWjXVavR3RCdo9i+vVJHOKOXsjMCpwG+jO
IR/pI/L6En5D+DUNPfZAO5tcWmKYi3SAb20AAmYtKhv9zL2gDWLOzMQ2PpcT2aXuurav096Qs7rQ
RSqwHrHbI6HGRfU+fXPkkBozP1C5iLwybM9TrHOM81JdEEri3CuPrjTo+ARe/as0bp8ozuaHJCW7
qDHrzWS9YG4MsXZSJ6df1Z4bV20HzyAMfUcnmWdh85X7r0uW0v13GPg/ey11KheLXXGv1AkwQNPO
VhHim5v7EBeLMNzAp8lJmw8/ioF20v6Uvcn3xggJuLNHUlziM7o/0o7kJHLJNTQa53KEV7nMrVyq
9FfgPlOr+55BMNyLcMwhuKjp3EoI8zHANQGGJsdNwk5nRPBUZCkaUK7Hj1PRlwmj1vlVxneU4uhT
al1JqUJMMjCWHDpo59yVyErX6yWUa1PwA7uqOD5qsqOnciovGxhLI56UgXwQV7GdHhzLdElynR32
+kjCqDjQplPeAtEo6S2qsV1ixieIqqpjvrBz80eNmr2p99A92amCzRJF4lZZ5nyhKLRDx0F/0y07
5d5LSG025HMm3FVkJXvX8EAD6UJ7Z2Yl9LcuUHo87OSRYA/C7e4TKA1faW85tGeJyCa0IeWC1ax/
mMsPRvxoHxhgHdJxLbCI7wLR0QUxm5xus4hneKg8xh++w/q/JF7SHlLTCWhKyBwYCbpzoU3yUqIz
DYY+eVFIplDqVdF6OWdT658H/90WKYZUHtr9BASFHZEhtmO/CmUdL78FK5epcR8sdMNhR4D8+WOJ
VduEyZYspiV33IpzlmybzChoSwkt0vS5iN+eh5yh5Szm62jl90b/SCBIVnUg7RiRUu7jkP1TZm4J
WsZdzs/epM23oFhiIf+w5Xzi2L/hNesxl6laaKRoAlf52Bi+c2m41o1kaqzS50AsGjjfyafr0k3I
2ggKVlLs+SYQ/QUO4iNr54+BOsNWZYyYwD+q3iA+j0V042ZbZUk6quSYdVJEkKPRe8XYAcjn0q3u
npysMHcZ7GcUajVxqKyJIGDPsjgJBvZ+S+dJY5qZD674kDDzJh6mFcDgGagl9CWl9o5ubd7k8nlo
zNrDTZpY2bigRsms2aI256d7Ip9TGjoSs2HPn80TVGrdpitfpPX2aQ94N+vn6fPTHGCL7xShtAb6
y2SEepwDLTIkmfo9avjhEU0J5rOfVVG0GuXxZ+XPDBKXVQ8EFaA79HCoafcUgzQsoAprZ0eMkhzm
0iqJzq0pXl1htilxX+ZJLnaOmb2N0RbTpiZubXS1S/kNg8hwyIktVpwPXIdefaSQRZpVNlPQ3t4y
46alrla908Oauj8H03nAGZ8kFYw4qnQoEr/aCwPigqBVCTFBiu+uCDxPbwjjZNVnVW6vhzsxLP5N
vXvKa68RgVopg0lrifL48mlMhYfJuQPP3HUqZlZvQIrT79fEifkD0grDFfmXkmkT3W9hV9ACBeUp
zlD4/xKh6mk4kbSjRO9b1NTe20PkvTdaZochoN7yWf6FoKvL0Y+nozvSntsBKjYrFqWeXtJh3CrD
T1iWo5IogpoNwMDxhJ6bFrnzbUKYScJRbKO/82TzoDw5Ik6KLtB6+pFdIpx8RMTVe+brrST9YRqK
yg7mKB0K1wMVSwhhRjYlHkORcn51L0RQeuu26TwgxmljKl+3eCtg6cbS/I5jliyXfBqcCY+pGi+R
BsD3WGxgZwH83z0UPGNC5T3vZhJP0KWEkBqMvd75qI68dhRTHAF7guJP+KLQy87wZBT+XoMa/IiL
3DqIYxGwfCH2RHYAYw41ecXoqqey4BJiijNYfIUp4qkSiFGV7lwHWFZX8NsDv4qnYY9+Own8yxdb
36xAW6NpHZEPsNU+fO3LxN+xFN5zcJaKOuxTzX/Bpun8PVOUbeE0Djew6lK1utJLa5hWnyx8TbTV
RMrcV+ZUm0ooknRJKJvv801AvyBdP41PwZMsRy9cM+lBD2c0U+D5Sgy/zxTZA7r1EnEIsSAGPjcr
/e4EY1zgg0JxlyEAsDmvDiUQtw8SGFzdEr/6Mn3g/Xh6bWg1CSeP82r0vJ9Xxi3q7Dmv7CfNkirp
uRxnKuegzweWt78tcwOz+sbj++mRC5ygQdU/n44SE3g02GqeyuTNDU/wn1RbNpONzSJ5d1mwyrfC
MKmKu6Vg/O2eoUXMZXGYTkDmk2310po7eNCwfPOXZX1nMu81j6bi51iutEb/VHegkodq3+r2L77y
dNS3v04Ru2Y8eaBtWpBpuw8NIsYd7zcXOr6ROJUTVgo/i9AzIjpBZ09e6JPewohFb34Lqrsvc+yX
HQluWRDUEVY5u3lEbWW6pqrWsPEWsf0TxLXYietWg/aZ3VQ6zCWPmxwpZhBNFcRnyb0fDSbcTupd
buW3Cnmhh1hcYW9tnRMQ+UK0kwJuRvzrX9QaoXIo6qMmHMq/fjUS2D1LqnJZUs+XnJs1wv1IaR6H
5o+wcvi9s22g64m0hHFApMvFaol1dJbbYAcoJ3+vEOxwqKw/GyCi8CKERA5o8b7TJN+nAFp39L/q
AzeIEVt8fHarjj0K4M8e54snNgfpAXKdntGmxpJk8kkiQLtd+pScaDQnjMNRxno4o7Wozb4cmcQD
sXTfqQmCIlIfRxeOalgNQATwiEX6xIcKAUovHo6YlF6/2pbZkAph+JbUG0cMi8pZhJfKrUhlOSwk
cYbDFhLkaX+s0Vg6zPhaUdBkikCw2CaefqjV/Ek1/NxGMiXfu2CtwqoIqTGekY71LbdnATirZE8C
64iJfW0vCRKig+aJ+Yt4grpQljjeuQCODeCqPe7tQfZzgHaUe5f7VIMDFBwoZUxuz6GPE+WQ+8Vr
eV+MYCNybBXz/nHLzG3GwEQIO3n38mT+qc5oC5SEeMYZSe1PLtOLej4kxWlvywjHp3OpJZjoaAST
g4/nzAwExmp7Z2UaWNwKZu7qK6nB+n4E4CQE6cFfOXD4hOsMOj79zzzu9vS53wA/pBDvnuaFQOo1
sdH6+j6Q9GFYUphz0/ren4sSazQOhRVN3ZJQqnZ90lgBJc+qsOosBKJtt737lOXxUeklcNZP9F4v
AOr5dYIYLN3uzCa/Q3cZNCKanVUuJUS7PJTP0FeYUsdeCv2JhH/CihPNNprsGbUK79hVraVo2Yzg
79pWW82Hea6lbvYc8NNvWkrKsJz13IDV3fIYFKwHZn9TELOn40NGGVbJDyJlSvVpOiu3xit3wWPU
dkwcCn/k1G+MNULCAsIH07miv7Go3bDdpFCB+mszh8WXSPD8LjUxpZObalcz6Jok6Q5OBZEi2tPX
1VacrxeKYWOvgUaZSBwvlNGOYiQup1xo+e+sR22ZljV6W481nVg4KXX88WmvWHCzLCpGigMUxKaT
hEjfFEGVKOTFd94Ss9ChH9knqkipkYSFnC2E/x3QkbEcGsPmspe43cfY5G0T8aG2r9bvZOS8b25h
eMtlHfcDb7f0giSSp+X97LmYD3KD5sqftOXAxsudtdhTbnCYfleO9fznibSWwTF7RLu8Zlxk0ZbH
jtLiMDx6CajGSU9cny5uZV7lzc/dF4Ge+n999vceuSGuuW/Pp/j98N/ma/rGJjkpMkIEvu+1GiPE
iAvFHQTraaJW7J7swjNZ6uho72YhffU1dP0ZU+82NoQf2FEroaGLTLt1AlNwRGnNVwVr7JjsTUSo
eRZHGwJNm7JIL7NDM/c7UXow1xv363sLjI6DY0nqVCULWrkKlhva7D12yFXJRq8TPxMJdWVQewgp
wnIWqwv5BwR0EvuufAJ4yVwWyxkMimd/WzcqRmd13SaBQGwLj4NrYUJYHcR9Fqa5qy+oiB/LQEVU
fDcaGfmXVEw32rcONBc8blPT6993CIhdNi/7IwKsBV3uZhLFTKyNRANEwKxGyfYdF0Hqn2KUaB3w
brmX+MVfvl4H6/CFrRFRp1zfIgefUm16J2pmdE9+zEnGG/2AyhW1kL6f6K7CTxP5AhTwDfw30nsD
1jPdNS6lnBHhvSg6FUvfN54quzf6P7fb13sLVnZx7G6/dK/ysSDtzodEfIjha5xXYTGCWDkXdd6I
Lr/xB85BGb2TF+aGN6IutIgv00vlnYGyi+xubII0e3bWM3FyFO5GgT5DLHXwQhqCOEJ5PZnrmU+M
JLP7S1znkx2yboxKkwAdTXXuR+yxIuQ0/yNS65qp3K+lSFr36oOS7U1V+qJ3njUZgYq2alfJjwdN
VaCBKf4ud7oWH0GHjulwEa9zgHY/31ETYEOiBscZDXTn9R60zAO2pyqIOmTq8j+RmIV3UDLkks3/
1vm3+My8NzdpGVYthrqiXAjFftzXY7XA0TbCnC9GsmON5i+4qny2YOpYrDNrd77PP3YvDKTnVzCZ
OXm8TyF+817YeFr08drTy+DwF9PEJIWKtrTJVkLp67cm9DXrv0LGV7n4eR7AdSJJ1K1pw7Pr0dFC
hUszjsz02Ej2yoF9FsG9S1vekC9uD+Y29NeEbC2N6jQyuDpwzvn0DJ4PMKOCWZr5EpbNPZy8fkUY
zEPKLlzoRPg8FDiRchRuYJvl2po98Ep5/g1z1caJMQzEsg1RTl7EW4t3zEhcIOt2c3Mvd3576dxL
8iI2aqDe8Ia8lEV5pWuxm5bmYYArfXvY7ewCLJ542gy5AFqFd94eTI55zAbWEzX0rrxy+T0U16Uf
28YX4zYJBj/afy39Sy2Ml7Gz3WaGUhvHmlVoxlu3zbJnJhFog0US+4rsNivzKnWRhG8gmtWBJcrc
M6V7IMyCX+/ESFO/ses6aVBXXHvRUj+QKh2CabUMmoiZzqIwGup5tNrVWhIntPtXN0R/b6B7i4UO
4CQ84GI9KkBxFw2+Q+FGXIClB2n37SIv47VdlHXiY61y2zU4u5LyXzJYUcnq70CqDZeJv16vL+Sb
HIk5M00N3XNbxjsbtrneQuc1cvfsxAGAJM8ecDNzizv3N4nAUlRNKTKyeYcaQ/C6h9RmLCfnMWjB
pVpNefWg01LEfYGWrkc+1FYwwtshLaNWpESMTmUKFUkPY96UG7r55Az7x5NBSMulYc2/cqWsi8iz
FjwCTmwGDzAhYJ8e36Y+5w/wQlqS++oBT0dMs+BMp3MrlihQ3X7o/PMzj4ZwGPBu/gWHDPjRetI5
fYwHaggmZZrWEHDAEjvC7xgAq03vKotMuWk81aFgg7jcMGHBFAnZcipHjilbcGPVJ+3HNYajslRH
Ush3uegRSFx8YD6Mrz+MEnB152JS0C5JqdEqXn10BQ44mb/3K0DVh0gGBUzUq7XssB7LcvH6lA8t
7D4d3YXCEzT4/GhoWiT5Ji05aphpBz0QfftmTMim+MlUad8HPWUWcj0xyh2iBhy32uMfhZc22G2P
X7mvWORh7mNe7Wc5wTVTdNZwG9G1q4I05XcLsijHQAa4ZJonjU5Wa0Fs3FpvAokXBJcKIyOhj/GS
hsKzQbTV/O1IhGNTIG0foqEftF2Qdzd3j9aY9j2NM6pVuJz4LRMAyNj7Cx0GoympjajxHeIiwLFQ
c7eStrmeRRc8IGbtJSFJnSWJqSRUTdSBWMaJVX/LAmPkTThKQQjWay8w2Uv+nHZv/Iv3jpIwOfdC
Q5rJDqNRHFeBsYZ88Lub4+1scS+l2KzqTbUyQe4+KlLcNC9TW7QzQ9TAdU2z9K9/j/GvigLMkQra
75h/BKi1gA8RqSisE0JJxTrX03gVQsaj0qU/gDymtlAY2lR2MM/RpRIocm/Mnwb/w+MU8MonXRLc
zEnBS7sWOs+WE0jxiJ7EWskx+Rv2Ufoh/8zCCpR1gIIp4BPYKDoXKDjmv67J7BD6BL7e4VwUwKv/
8NpBrJSexVeZgOgbZiXCXomhLeZBiUIV2Jyq5idJlGR0G3x2MBSbzPszaKc1oKxYHNKtyJOOoXtm
nGiJ0d8wElOMq62HTt1V/IyCMFFRq1Y9GX4vWpQ4TibcpQQ8Gn0fkKc8HDzqF+a+nUFdeIEpvK7v
f9O7JlJKUGhs1abtszn+TCosg71OsI7V+0KeZAVvcTxSWQxdg4Vs7JL+TjsqhIHjM4/6SzeqLkHL
LXcGN81A5TIS8o3RYmdvZBWX0B6KvvESTTipDoBZTTwcr3qh8hTMH1ZQ/nGB09HLjxxj3sttHN3v
4JWlFWwQbenAjRcucBUfL9r8POnhdylaacKbkxca2GkDDdG+rnFRvNWaxHKVHK7TrNQ/UhV9W/Lz
XE8jJjCVpAs9E4/m41zSUB5FzqcaOI/oipSb5VLJFnEdgPUm5LBZTfKzQjaykGsgEPfAw71/lHMU
Go/s4PgVOz2PT9dEVCsGXv1QBU969n0WDBQ7Rob8mAryonPbyd91LoJvr5Z31uvwtR2N2dePCj9C
A+RMQDQGT5CGK0SOP1FIVAQ5rsLkeNa/KrlAGCNedtBWEoH+svDEFP49QPhfxs2eCL0+Gvh12wUX
5nMV+8TsMSq9CtS1k8PKW52kUV/gwnIb5Czd/a3hnvXgiM2dgD9Cv7ucwSuFv5bITq4nwGrSR7Fo
ZWcF6iXrLN9EAu77y9hmesjKmWeJtxE2RIfz+8AHY3rErtrTRodntvBxBSn34NCTEOHAb10j3G3G
xwGbukyBReQ8wPZKtY0rOwM2j+NygiXRcUi4oRLskgKppYnYItF3zinRbd0blTDKQhA/CzROgq2j
LDRCFifPvi6dkZ1VUozF6acgEe+gIxqFhEj7W4f1CXVoafdrSzuptjBBIFe3ZzpnoMIZXZ1Q1Uux
EMA/EQFPlxAPYhisfGEa2clIuEQuOUPPRYZ0ew1xfxngqmEMSmifWNvYKUCNfOxUWUSWU8iiCQ+F
QaySp6aYgLquxUfjnf8pSsjnd7OPcuNgtDpuSger7GPaV5LDbt3Ikh1a/aRh0tomG8Bcu+0sfm4o
BIDOfYH3kVN9jDt7NbogUrMC5IqFE5gtKo2sMr+zG1YBFhHpj8rqw0BhOm3OvmzC2O251QJZJtEq
V1P3bf/1GiVyrQUn+a5XwtWCuTskBPhZtgnAmPp48LuExUCw0Wlc8brHDo8XuwjXBvbdb2o03tuf
O1rZz8ZMVuxiTQo8y0e3iYvFfZvsN9xX7HohehIwCY/pSEQ1FmFfA97+aVHWkeVuV8fFSaYBbu75
6olLWQ+G7AjzYkoGbPcB6rdY9Mmp2FjilSJozE+Cbu4V4eV5jaANLble5YNF0Jr5CWB6fSp50tj7
ZaeazKxk2MMrBLP3gRfIxUo/xtULPoQP9ZoB6FXRUuxyCom1t8TgrETrvkKU4AFVeeLl7TJBV/dc
iGwxpdIzuetPCmZVRJJnCPB0PkByURyzRQLykDIylM9+K9i5id9Ht/VKzzAAyDlbAsOhLKfiJ2Nl
vc5+YK4lnfEJQHjn7EACZoWGysFQN6GTjncuqMA3FPUQ8KEfM6RvMxLqtPh8l6RKnm3VOrtsKufL
Gb4dZiaEXrPQF5CyhUHNSCrK7VT7jbsEg0sjBQKPFOR8ug2qHpUHXDcrH4K4l/zXqNaEpMaGVWZq
EYE30Y/3MH6pAbhQSnu4EBh9OeVAP//JVqSMRi/tZ9K+6yWce5gbzlBQLbKkujuD1JEJyXXghtdH
VqrEcTyBrhWZJcV6b1I1YgtHVug6dPhkEiLxles1y8u0yg4ADWwYjKH4z2LpK5ZmSGLfsHCnF0B6
aRS4dUlmFHrNstnQ8Gjxy6C4l4hVSkJsMlAVObgdTeygfjhZ9q/K47WMLl8gMolTJQH/URGKgQ2S
1y8A/tafWgqV+PB0hU2eJpZs11TtlwDv2vzoxcr0AxCdhoIz6YRRZQTwRlUe7nUaVVQxpFObN7SF
Q3RJrBnpL0uanL2EIMT64DaJiK9/fHphRvK2dKwtN+1HpE292RWBO2RCUgaEelnhthxRW59IqeQ0
l6x+qbePn8IHx+TrdwtWUkx1pYLVKNzr1kIg7TuIN+4DTLGjv8dCE2K7A3b4g6146g6iXRoarHvE
nJs09GSKffxQGBhJ+J6hYzlfEwjFwFyjvkDdMM7I+z/TIIZIU5O0dr3L1WFMd662aHl8QMv45zp3
aIBbtxkUb96PK0e7F/zSURseV9RUoc9nSEKJI3v5aKxXlH+m69YMkoDPczsqm4LVFErsByyaOF9U
LI68bJnoCk4y9IjWrVUcTHkOKCU9LEStxPooJqNkEKhhyikFLjQvbGFpMtkEKqYeBuNkZi6nbXFN
87kG0agtq3hXTllgPExzl9yJfZkUf87oBwbzBMuokSrsmjyOAr1+iciVDxUYvCO4tJ/2ybH1DodL
lnkbRW8iNOjo0m28tPMEiX31o4Cjj5jLe/m1yilgQfCJvrOpTLVVkBZ0KRxk3GEvWgApk9ZwPdOY
80KcX+L82fDvFLnecc1kZxdAZ63v3SMsz/t5dd/IByPmTazht9PdolE0dyr2L/ke+3GfLOK1X0V/
AlD4t7V47vhVE8ty6PB2QcUWM9d34JuwHUbyPo2pLc3RwXIul3tGEf9rCG/t8R4bjSl/xCcPrBlm
jAyqoNXf+jq2NBq4bnn4dl7jVO0yu1yVsPLShyGs3Gd/PbL3KoBTXfLJZ0cm1cowdx5IphMaVYSY
xkLzSTeIVIwCD/c0a3/u+x5PYDkXJW5YRB3ClZRAUSyzpNdoAeKYFpaeZV0uNJy1TVeWtge3G10J
idrt8EMRHHxpN+zydrZDWKhDpe8f848Nl6sC1ys0lAKWSSsLOcMYQTvK9HgyxOHtHnM15yVw8DJ7
64oSoi90RckbbTGKD+wct1uGKC1hJDycjCsyFEAXWFaNoXapEAtxGLsYlcTtKBlwi3PaUjCblLG4
mr/ySACQlIMXZC13r+twb9TiIgM0h6YCJQ0O1Viy0/kgJrmGQPzIiYHQrVpXk4yaG8bUGV6Jf18k
0oXAyDPsUXVdF9sLK/dxSLcUpCzHTzlcrw05eGTOeF1YOBOB/TByQsWeuVexf+0K2opRaLmPTgtE
/+JQ19bBf3YxLFccVel7SZk1ffID/mebHuiGz2yvvLrMzgTh6L3D/F4+ZPk0Ffv7zIex5pwOAo8p
G6fxJUA8MW20B4sUTmndxxl+qM7ricxVjDM6MsVAGIDERGSmNWUEe2IjDIHcAKAZPSVo8lalwBUB
+8fqjUR9+uVi8aXdNh5NXVM+L7zr5IGbMawa9OVQCCBG8d+iDJUnqioDVYly3jCCYsyF4GDuNpay
r+5qtHDDrTOuywTkZ95Rj+7brJyjp3R59HPqrkp3acVHNCW7IHQaKXNUS/7uwCRfCgZZ0lo/gOTV
73rXzeBtjH2yeHpSFBBitCwBaAwSCS0Kd/k9U1dE2UOGuU0xb3afda+wElqx3og5BhuxdDag7CFD
Wk/0AeXHJlZpB8lR3BNkqhk6J6H93bZ/HutRapBWXNJoRIEvFA25F1ZR4HAdVsI10iSQMj2mo2x0
yxAjcJ/NYq5agOREHMNbYVV8Cbstm+B1h1ZySW3cI2KxlPhYaHcBdWgAobz+pECH6ncWZX+GcbbS
v2woT6tzju17TTKdwp4fsUvAGjJOICDdc3zzbZ6UGnPJI8g/p27RRae+pjVs4oxs+9v/w0i8OycY
NIqosljrTovxRSQwm+p8LqMlZpQMccK3mc0PBI0EqLE79YoJNvDDrB1kzQOQVOufyBPO2Hn31L/I
mJ6jmrH1piWooZwAp59WNSIi7NJ2aFuk0MJhVBWQfmHhaPWSyZ5mXi2Tp28f/TCllMBcoIv+24Vd
gggFRJMpOSzwwUsn/2cncYYBivXXtJJdv7SNL56ytVSqIIVtAnny/Lgn/o/vd6TFG+89gleewup1
++VUqngto3bwUVQtSgzUD9ywF1QKh7dzkTYdcAwZj/LWflt2iCf3xs0oq+dkmShQm8z4p1PKiWaP
bRb0MR6WtkU/VKEYTQYJgRk5Ub1rbbt6T5ESGBbrkaROL+pIbtCVnTtcRDvPRtvA180cu1YbXliR
sI6pnn0HvbtCjcHSBhoTrYHM6DNFQdDOjsq+s1DS8Q6pBfIQci8vLc6Lw/kJel0VAY+d9sUSt1Pd
nGyfqZWwCTqWsSaPaOvEZmZ4tGKa+QQphmfL4Iwed4/RyfuTrkU7QmmCpIHDHy46w2bKlpeFzPo7
SbU7fna9l+m1y4y98pT4IbXk8lvLmjM2N2Pu9WxHh8FwyhpJXiufXMYC/epzy6d3jEtGUY2efSAF
JyuuImgy7xJOd43js9a19oMKdIJEDtt4ns9zOVKs5B3rmTgvgP12FKvmHyigXB67+rIlv6RbQMFL
9e1klFwr7HDPvhtEH7mGKPcPXyk27o13Fe1cYAiJ8DWMZPY7VRcAw5f2krVxkd7tV2c1ZcAzDWJ5
dPZaBGAkIpfgyfKLHvhHxz+dgI8GSlQ+aADlgXTFm7KZyZLhrsLZharHoGsSYRwH9p0aCD/dAae9
dcDUBOtrdT0XY/QsFb8dV5S9XHUuUeyhNPMLHECrizCG4/7Skn7r2OiTFDUCky3t2FAqgeOqpIxK
dj7nIv7z/F2fOyabqJe69EQxv/TqEOhZLAlhmjK7SZ/7eMIIfxDxTWpFYs+8l0FWgIt9+k4gZtV5
VK7Dn/cavgU66abUAcZ76KAkFwCDd0b+fKACrtd7HFcETzDKH/g7THHNU6udBu2LYvQP9ROHSSUP
9+Nxgh7vsbUVjbsjzfTtyE9udL41ACs3mL4jCoOwiw19tjfvSRhNU5JTb/wSs8XDvEF1lTzSXYPO
rQUL2IY7x/Xixv1Eu82tVF708Tt4u+kVMuLKC9ecck6jeKKSM5br1R+okFdqgU//rJgtkGm+3aik
XZMp/qI0OyWeotTTlDz8u4t8EpRxJEfzZF7uqUOOh1zvPDHo2doY6P8PIdkNOxkjn0njqbsw0ELO
TDhyD3YkHaoVjUrmfJc1Ey33TLGGUkOFjYB8g7EkH3NrzTE/92VrmcB1NARReJYjuWsDfTqk8Dyr
P+U30XqsugescVjLfA/XO0ik7wckr5/M9LXAtt0bKfgMz9+0k9G7UovHaulXSPQ5E6Wvw6yGk54/
F4bUUVdG95oWHfn5M5JfyiVajsZnAtCcZ4hMZx0tCLn2h+VdWRlxki/ytxgqsKfcQJLn3DjTOyvR
SkJ3FeB/6lQzQ5bhb8YGzB0+gBPTH2sjs3+8xU3tIYlzMJ5o3zoBtgG+eywyCGbaS3y8omS0hEHI
TqqqRgHk/0UKwZBKxOQ08VBOuMj48n9JXJBYvuXwZcJ0u7ZdpN0D0sXUYgFMTkumTKqJj6MrKZ95
bucezo8C0UeiAgrYJOhrTfbYMWV+dcAGJkxo8jw5yv0CcpPWL5U8YLwhhNjQl7S31cquDjNAKDY3
eYdl5IdD7wcDhZrDa7u9/4I7vQZFg+0C9Ft4VgdcbP3YDw2LOQ4qgj8904rwKLFhuHkAEKUQiNqW
wkWtFNAo2n9vJWSizpH+btVB+7F9Em1MX14uRRw3djlqjwdbRw408uPaaxtiB+yHu/XLFeSE86Uo
EN6caNEDEPv+lw3vKgjwQkMa8NV89SCjCzhe0nh0Ybst8D4z4JKefXlyTxmutQZq6tkNspU+53uR
w+AgAYTjkog0P69Hv7ArxEMUC4yeHHeM1Yh9qPF7SUVUYNtIKdkRZOmB17HyQd+2W6GOblioJCqd
vfwiW+MD4iDTN2KXU7qZkTlf46WmEj+6Gw4UyXENoTUpMEkZxHH7IZOkhM3YkHCCjS81qWcTFPyY
fLU6/nstL7ZgQmUvyqn32hUOEaGG09VZ3Yr+tOYdzIJ4APwrh3AyKXRJ2rt6Vq6lOO7HBFIG4y3M
2F47AFsOG/UTGMQh/MfKmmPnNtmG2PaKQzKfYro8MTRxopyCM0NldpifAqa+xzlte9K4U2Mw+FM4
i0HuQz9EzOUeA/NtMu4JxCoUFZHOw5+J9QDKDJc2at1WRcXisfHSyZfxyBzeXccaFOkci05Av085
Uph8gDP6kYQ0TaX5B3g6Xdda9iHJDMfSJ4Z1iut3Mm/o02zLx271DDdSCpSFIwDJi8hs0iIm0jYX
6PRTP0tGI3XW2xxGZ8OYUc5YMpKTjOpZZxaSg1biIaFMPTM/QSbMK11jzxx5RDeGZ8TYNLTEey0J
/Kceh1xYi8lD5c5QqdC/l9cdezqWaRyrolbwRcvKuUPcGSlx34+98znEKUhxcIh+fAJCV5hXPK5F
dkODwvj4jzLhJU5nsIajh6BMCvq+g2oTUcvQd9vvLGv+PVujBVCFbL2pPoWY2WAEgmIw/+VyoYXa
TgyaRPQTc3L6RCA2htelcia6jkuGWE4dKg3Ju2f/bH5G+AI7yAbQ5Fy2Qxxu3h7Hx6SlrSBYlzgH
5kIh4qRzY3wXemPIDhEykxPRI08xqGdNp8uv4uPrJ4bmiLncpT5vUd2gRHFpuHhcxakjReNA/EmK
MY9VgYUy/NaI6IZGYvdEEUGHy5Mq+vW7V122/hWwRrTeDM6yZq1oi5I0PIWrnHT7l5BZGeVR4d67
hWxGq5LSw/Xj8ypzpAkRAeTgdCL0yUZs33g2cObZHmKUd1a3jKRlIZLgwqByhiRZWDLZJiOnlvke
06zBMkcTMox59qlKbKHN7HluRNkT0dOiZY6w2spchvlqmNjhuGs8YOecjNq2MGHEBgbSVz7IfSOn
VuFYOvcetwQ+9mjuIsG/ibl370U+TpoiXW3TyimMsSxPTpW87RSdfQHHGADL630FddBavKyMr7hu
tgT+gFBkMnHQnsL9yypoSDnRK1uP+heLyEhqWALkPcDD9VYRfTFGE9ChZ1AmkjYTTJahL0BpX+Ob
Id9stEYeBZP6kemfdo2VL652uJzsSpGG3Q0nYpvhvH/QD/FRBCc4P/BUpV2ujQ5wQSlW4ZBYrwlg
SROUAAxS9Al77olztI9fjZszO1SAfEwfjg2uIG/aElTlL6qrwiDyWPJejuziQ+5PH/cHZKuc/3Fa
d0zylRUL4T1UNwaOqLFaY2Giiw4qe9/cAIM8E8Ovigd2rOORxc17ry0gVZRmsgxecp2ZTfm10qCQ
L+I8P1HpTQE46IlZHTiVLqDsBhH7yrvSc7+BN8+y4cJlvGsMmzv//8cAwNLo5quQOKskyFXUvK4O
AUr3i+9wuGLPmZSAG4X6qy99JiQiDIqKyHzIOtcB5j0EILpPM1cJ+UDHSmtZByU3mcxBIOB5XtTc
j4UjkT9UARa5l4hNIobmkiF175qeuT8lQIYyolsRX0NeoVRwu/ZbKBAieMHvD7gfG3l2Zk+awoO5
jWiZ54MUKFW1OPKZxaFv0aoEbRwEiEXlzmOiBpBO7946dkFyYygxA13yJ3H69g9lmxEBl5vc2hnU
uYfpCjIWr0YgSTPgw9oVs9HJOSrSCUjW0qfI9w+nUroufmWKaK3OS0iirO3SGjlZw4vtxoNGMhZt
0QE4mxKgfQAqknKaznRBVya1O/2liQBC08DUrpmhrgPDAFlJRY7o/ROsZ8Yjly0gAh7NUN7lEDnb
3vY5aURFGP+yGQtP6eelJH+qv744ikMnaD2a1lWfb5ZNRkoO5kzOSNVfyWqYp0qoeMSBT6dfclvt
kbT2Jv3cmwnSQB/yfCLVOcAcoyaSL8CJQEBzrEHSRjv30aF6UpbTNwUjBvV6SPJNt1JTq+KFtMR/
NqrvilVDHrbKAZW8+J/X6+Hl8cNFhOMXhR/7+TmH47glt2ulMbvPYER5iUw0VHL2AkXZ0s18rp3Q
D34u7v4LOiMz3f5zD1YrBkLqIKiVgGWCi9yAuIbx8w45CrYtsBUuMYddnBN04scsp8qkKst75sGu
sXXlF1mqaJBwsEYmrTGPSgBjASuAZx4rRnfZnvuK9/uQNRJYm1r3xR780/4SgPgwfpkwastyI/+T
iiVupaS8z7CbaiZ5/Jcj98utQJRAbx8rCQDNQurparVwc+xAVNK6G8zQ3wdG+peOXz+klRFfExYf
Y9AXJVR1fZePgI9As2lCHc9DWU9F9VdzjuM6BqLi/AClf3gbVDUfPIKlAlT3balKBGLz5tOWv7re
jztDxFHfVTIwgkYK/DUb43qtz25nMWyJBlbmLG1jkvRzPpFV3AT/A/dOk3eOMg1nUe7D2BeqAFnj
6dXEKFAoJGo6dtSlCsoRZW9d1Sx2BD+xYLROHXa134ha5avxyuaVK6F6myA7LlUhVpDSEZiinfSt
P6eSFesUJ8l8lyb/B+xkZePb3j6WG+9/h+oAiw2WoxQgN0KOjIeMPRkqf/M5qrvwklvvjHIHp7p0
InEe9+J86jai53HqOAx3jLhyOR5jHh9djNHfufOvWtq6WreBd0+8OXzkat0Ct1vLKRMVSWBgYyMk
aejRru7AB9jv83Dm7Au6NIi2Z8JbWa5naenJ5ntwAEh3M+HQbqDXgXuM9h0/9ZQNGMPd2zGVaaJ1
d1yuPAoGE4zAPv898PdLnHzLiEiB8pIZ/hjAIXlHHS0DIfDXYheNvMM+LQ3pFfHyKqR0KvTBXYWt
JDLjRRUC54qOFzYoar7Wdg51bGo4K/jaXX1eRrdg9ogEleqSDL64qy/+aah3gMD1POE0L2Akpnyj
oPcr7dCGWDm3nsag9sulNlVRDx2/T1axFSWpUZN/v+3ZFWpwgiwMHeRzugksnkJ8IjCGWDitBig9
tCN2pArfaBdCc2HFRvtNOk3dOFp13hl39+2l/R69wXjtvXz0hQNz0QMDchQo2J83IPWTSp/E2JRY
M8/ZbgzlGBycbrag+qbGO2Qv2XnrkQ9gtll2xpCPGxoB1W7Ths0cySMToYKUAxjkhQObJmsgK9j0
CjItDhdSiXuJ/Z1cdREOqeKvjtMh/3Sh2tDuarunXB4FptctS2g7XvLplTo9E58oNpUJCccBMDQe
v2O8ZkAglKYsjTVmgaV6lQtAesLWRxkJBB+shPctNQpGt4+RWTNWuSOwqg2Iz4/dbTuCNVogJJ9i
Tugi+Zb9tlVDRUvwzqh/7vSCyG3kFDKKJ+g3et/bS5sAUv/a3jvWQm9KcBf9twanljl+K6jWlVd2
Eg1sM25e7iNAr0mlWbIZCO5DGPiwH1bJ6Rb2+LH+EDuxg+61qSxMYPc9owSX7EqhISLZmF1o5cvm
rO/xjkcYLsTcSky8fmgwaVZhW2dCtaR6locq3DGt9vVKxfiA78j+/XD7uDEXCOCBj6E+YJk1IWjY
jn6aueqFMVh28vtEfuNBeceQKN4PcUKGhzH85l4X9UalSO19IgJk1r4ZjqFQs+H7Itsfe7XF4znp
DepM5rnuRryxdrK2I5RRGx9dbkYOmAWnHYtLehDA8lq35z1pED0nAImhzCaYQByTbEW7D5V6c4Pw
3XK4Ed/450/MP3oNxrMj9Zy7Wjen8UkkQVTAWwlsaiMDUHyG1H0Sw/cR5yVYHIq27hFgAhMS+/Hg
O2YUUYWHg/q7GoZBQeMOYt2psEYX8Zoolq5wj9CNzon0N6wg461YEE/ZQRJugfIE3e0/34if9D7u
VRZ8izB+cJpArfZW/pa4dc73g9Wz6+NPSjMSo9bA/CJHsxDDTivTJPHSZpujhCc3Ri4jy5rDqv/3
tKtwEezridezyQm1/Tl60wlQw9rd2R+ttmVdpeyLF76RrEJGtYiuknj/ks7lmnFa0X0Qv3V04uZq
k6FOpahUWpamifKv+Zh8rHiLgoQyDC09wT9E9fe6mfQ/HF19F+ZKE35aBPzto8EzNJuqKmtQEPHU
3hfaYqrrvlJHWYnZ/lDOPNN84gbEu1MzfHVu8Jk7eCTffbdfgOSTxt4Zb65CIQo+rdcHpr4qc82D
dW0fSOI/QMzYrK49MOZq2dqj8/ScEhLyhfA2gp0dIOhdhn+8t0C87g7nDlfp3YhwYu+zUjGAR3tZ
Bp3PZxDPhNIig8S1lb8KrXt0zsNwZUxB2+UzxIV13r1K57fUy9xKXYJaotR9X4MWiFAFF9VzSG9v
u/sPOmyGZJHVXKogB9ZoaXuCCYQ9T2GFInyms1HDeuC3+xzFPc/RNH3DhNyNxO/Lxfk+PyNYBZnG
CG9QHuJ4WX4hRpf9sc3DmuBAKrpvlijFuGWpNdnk13aETq9d+EnPbVS66N5sAUtNL/GnmKxsKOLK
2oi4OIwSKDEd3muToQ8iPol5JbG8D2Rjkce7dG2w/yhMQYY5He+JsB9DF8vYXDiLslnOMD/rA97L
CRGyE5cwt8Y7Narhelwlir9doFp9BLLLn6OjMUVSyTsWWCrR8QMpFK79J34OyQMAbMSiawKB15iO
GYtiFLVcYUm3HAIZ43ptIBGct4Hm0wU/WMJss5/FGpJxzEUVIGBfGQWrr8QEOybWKhbhp9lpsMJs
DDlzxA99HH4Vw9nbY6MrG37y2ss0JE/rwWNlBqlWdJOWIrXPyw23dRRsIDGYOcFHMt16GQzveYSH
sCd+cKHS+wzrHdGID1XaU5OaqlAiP9+NVoMH+WhbPmROWe2H+h8fhWIZ2o8npKPOIv2pk547kWi6
IUnE0qTX9OhP4ZsGlS7D7jeqXiSrCWCW/RIPJrgDX6moA6IZwurtwEjbJNYyqPWCU7GyOA97/xPZ
g5/SUvAlHOZZuzuXakO5BvaGe1B67qh2QSCIpX5ieQzhzlIVuflz7Uu4ionyGxRT+C0ao6TAab13
oAxRIjkign/WBbKC06gy8nquNZh+tuxjLsV+V2Su5r5IAFLhnpm+UJ1V0RG6cmc1mSrmioJOU20A
1Ij/EGvCD+2Ev1lGaWbvHj3d/7TRdjM2GzthIG0g9+I2YjwD2CQIpRNHhJylaqMJdgP/MdIgDXNS
ZD6itKhGVBFGco1qp3qAilZ9/11dMKx2xCRrNDKVmVBkyynUxXEOUbgponGkT2P//hnlgVGEoCM7
7sXebIxnZnsGzW+l2POitSz30GfAf1Q5hd3hDmi6/ZjBXmFk1p7v2wduMN8ZdS4pniWWD/0BqECY
e1AaO4+Sf91JTzNo+ikuPm1BFpCTMySgQ2unMAqqhUTbVkyRxsKY5Z4xNc9g8vOa4fWnct5xPfdN
R1YLAsRPgSFT4BINnpT+vvgJSrr0YXPvTOhKljo8sD39yHkgTZKuCg4rkN7GRF8e643RPjB9328h
iFsoMzeKv6/znt0TE6+tUjdlzxyClHDXOaco58vW3LZnWg3PCmpc7Jurbvk1rQFmNgrDOCK3+cW/
8xtf8Ct68ZmFrEYqA+rM9s2hy4xfJFYUTUXLhGidk7/8d/Wi/oU9vQPO5dHhwr2l2Epf/9WIwf/y
UV50SRoKGfcVSA7uaw9o2fruE5sr/cRjxt01x+QmxG4lbiBZa3N+CrziWunOAnfArCXzYQOuZWzF
opTFMwEhvdQezBc6rOoKRu+O6QH5KvMjspKc0KxifZt1I1pS/oeysRsCoCQFWscoDZB/6wcOEZw6
bPpPiKqjs1wHPC2K1KFC749QjqdJaSqwmWNXkU3TmOB5roacsf5R8Jl9+ZDaNhBvZDDJSKpQSU9S
TwA8/rcOmigo42iaI/DJMcIZn4fJYOeo0sLE9Pj/bV5eNggxIJbtx6b1+wAGPbexs3bfkGBUomAU
dh/fz8NkfTUr7Ix1UA2g+stq2kK4yj/MioEo1vgm7buVBxWKNr6/HtCvf8+aOVyr/JacLTVANyrB
Tt3AVim8ZKeG6mH3j4IdDNlgXKXt6/b4btLfa5Ifz0Cw5QuEB1ZgAIdmYu3PQAnH5NXkSA1FU9uS
F4G+ZOczWs8XA2wZ0C/RUokaozb7riYG+mUDcrovmr1cC6OpmjDFn1krLDo4tZX4EQvhOI2bIoZd
lGMcH8FEaK8cxFFl0EUgiMl/DGqqoi9ndp0zIgs8L08X6/T5LXResJ0YKp7MB+Ax9KEr9cTzyLVH
wjWkK74Joq7uCHk//SNDJdJb9fNlvMhkneEy6XpJ5dTs44brUfom66TUT7dVADckWkU97OkMVxl+
f23ldgEyIXsY5FpWpBdiFCLm9K567ERjOkRWyXpJ8rbJOr6ruTMkYGsdQyh3zg4yd0VdOvfajYQ0
I37eWHL6by/LiJ5Jw5SZA60bSVx6G2E9ea6sL3K//4Pr6iLY15w1gCLN0P/CD7cL0mQJvucSzYiD
52KIZL3w5wihfID55a+akDoOs8Uu05nTd/uoesZdOBMy2TGPt02vO7XhJnMVLCeNry3F/l42ymF5
O8ZuAa4EE1bc4QqPnW05UKnHcQ2mxS8SVSP2p9UM897d9akMkARH4zo2MGQM2utuHRtAqk0RGrrw
MmoqHF7GSVHa9ARdeqJWIAW5fXD4kfXfD4Av3ARtoYFSRzQQqUSfwpAn2mRwm1DbyEbITKmhjB3K
850MxIVYSeiyKAvKkdI6TIuakX3sE9oKNlHLXYKUcr76faIJh+4NTP2XdIGu0fCc603XOIacW2v5
AY0nUd2tz2SovD+UeCkHXa+H0YNZj2Y4QfWo0z7BLpoJ4yVOBQpX112lOl4klF7LF6eomgQeI9gM
2ivDqMDmgxpZCHJyvJsjzKbPWxddjfgtlptwskYgWVEMXMDUn5EZaq3HOpLvcr43hvY0BOxjiLIM
MG7aP0cwvlyq+tba/QHVWk62DkS7peXM+HQp+PzOi0YgrKFrb/p335pLQuY6Mfx4K8WZXuvntVnD
rJQ97MLx0ZHtXrq9ra19JWB8o9wsb/ZLLO5xmi3LAXYNxPVthZ60Prq/TS/PH4LlkxJxzJgsqKHp
gYR2Aq4lbxeVumaczCDTkr6DpsQ4HvZMclIt9vDR2YjSA7ivOnUUJakrsSc9FTqZjZCjt8Kh6ZQ6
sNau5g8RcfXmtvmpB9U9VTYfbBupXsrTOVrBwKH3leaJGU2V+NCqIIz64kzGM9kBT6FoABHMyyOe
YrrbtDEUI/kEStZ3cm9cFKp0JzLF4DnYT8ioEEvKh/dO/LgpvOE/Wodch5DyeeQnAgeoeeKrtNhY
MM/auFW+MwO6s10xpqMjecTOwJvHx5Wa9jwxvruHQylQq6Z7teuTGDxXM8xbzFluuhcazK5HM8TZ
Iii8a9DFDbpgUkj8lg8Fa/R12S1DegoeTKsbCiO7YBADDOlwR0Xt9m+JtTKof3P+phZ5Y49yEqeY
YJxjQSFtcAzJQbewbbC6BqER6kE12YDuW8NEAE7EM/47wpxRnFBFIsVBwcuOmGmjA3WqiE6pV/lU
7Od07DsRMbIGrZvnF8iHTbf/7eejJ+zcDeuLfDQVR/akcdet7zIclZd/W4AcEvi0W3EwxjXCdIeu
SyPGq1bU+ZoXrBfwq6JSLaNMqMkV8xcbT5xiDEr15rPr3qCMTJPfxVeuVHvCqHyvW6WTI4n/66XD
2QtB5lrl41w8VcqOmsoMFCRarrYPtlnUemwnIgwRdDDcgTv07z4PfloM5UKqGVc4WY9ExB6phW07
Xow0I3cTqZKBQKbFQ39geL1YVOD9AomZIMM/nyiLEX4Aoq5aZRkroM2PyJSixSFZ9oNbKi9A83SL
OzSPD4I8O8To5+DeTLoVfsxFzTNjIvdc4CcJF0/NvUC+MaRXqJ7ZiXzCK4I62p81oc+QpmuHGCjV
ylRXFUrC2vl9gieMaJ7mIXz6MrBWqAJZqT3ENOf+T1qdCpL5W7jqPLa4Szim8zVVaLBhEjc0+OXV
qW7lfXtv7uuFzuBdlfMo+ZCdww4zlRqaVKa6mUdknC7FPYxZ/K9/s6b8ES5euEF3VuklOUiU5o1M
jLOL8UWUHqXF1jYkWYtEhMS5l70scvmCkCNGHS1p7RmyY4FsLb0kR/C/8lu2XCQsxMQBlIemXq/D
418fB9dJtxRCPgq5QPCOwhNfV/NIGxmKKkHHxTyD920Avx9rmlHNEDuYRCguEOyhnwau0r2qCcP7
ESeoayAX/pShGm3+vsvo3HihPxnt0EbbmpshGhSKOiEtJ9v+LrklqW4VswRhqlrCKMWPW1H756wI
R5yXpzrO/7Uenp/lE8WpP/zQyD7/O8gpB08Spv6NgCSgMc6t3aKMVvsoiSh7ftTLyJrWYutUARoo
5W7tVZW+kC2HyQ0Spkrk3SjXkVeWhoKPpT/jZNeaiAD0euZ5QhJoptxLApJvQExVmqGIgowp5AMt
gmiAgedVEk3fTYeMHvqKMgokeMfHqhXuyR+i8MST15ARGVUgSy5iFZlyhLqSVXF18k6lS1KFS0WA
g3n0G5zejSPYlM1z0JEx0izcbhgrYWfC/tUrIfO4pXGp51Jo6V86cXfTtzA1rgt7jqwGDOtnQkf3
wloHmrsmvRr106KgwmODUc5gjrn1ymSUhgStUg5xc7peli9fhEjnHVKaWu/IVeEcqJySj/E/X349
ZXNxi5k7T1R38w98ohXiNkwAm+g5O5vqYuoZE8saQVbSCwG5FxDEebKHzp1BHNlcxBAtx61LGLRQ
HcEG1P6GoLsIH9MANowFo3rcL3NrQ3UWfbaGe3TDBWa6HvU4Xul9qd0DOdEbPFrLYPsC/XDyML+2
qMFaUw5BpGCAjJ7wsPeRjZ1H+8MCZuIVL3ZkDc7lsAMY57nsaEaAFGWwQBbHSNnPKZTUIBldqFsr
teA4OrTqEqMuAKZ3iOm6lUFCVZCg86kzGlBmnR7pzqWHh0VYI5Wao+HyXVfvV6qdj/hMkARxUycL
KVE8C/yXCSvnH7/7oUTSmnp7SRslV9xkA4SRBXf9XcBSovbLMUimRbYQawsblhDc/2bMHpY1qyJ5
UtdL91xSYToAkDBv8B0Iyo+9IPVxtYB6O9Hh7b+nSav1Y5nqAgtzD/I2733v2RDW7ItLdzq96kT+
1gtoOn9wRP+xSqq3LhIYJmK5g+KipNc2BVVHKeiahe+i5gkwAyC2QwDBsYxRjO8n0+Cp1Z2yTMHt
el/6cCQU46kdvzFYCox3xlesHsWjtRQCOT+FWTUah3R25fCSeu1yKv0Duys8odrN2iCCO7JrFFJL
S83t/QAak0yyRlfiJR7rO6oHekKrEiVXL+XcgMPMDbD8Bl7vA+M95QchXh2vkFJllzn3f+Ac++ST
aO3um48wtaijDvp+nNSEFO54NbYMiOBh3xKciJkb2oIsu4jX9S19/abQY3VJTsJajpspb1Mv7vgN
rkSNiXcsmmkBZL7nBVk067fis438K7Qr2+TyL2DdNUKMx7FYgeb26aiQzB1sGdK1mwvAzBzblW5d
syoD7vrKVfAcpxP7zgAYwRG8U8xal8EFm486ywKAkaHI2t5pKUPnT/Qtd0HVHO2+nvNQYlJZhVJF
dtnwxLOJi2LACWNE2AdpKF9X+aLpuMeTTQQyeatZSR7oDT7sN7VtHMPUTaDRsgtj+1K7G1P9Emyx
pZyu0/4zevC2XuD/63nIi02cRLqxWFd8pvVir5TpvcAsn35LTpn4yH2IdY9DC20zsqGt9tMy24MP
W2lGVAPNwGPK8i6uFNNqaduy4SOxNu6XThTfy6P7rVqkHmfDY3e/fLmVUxbtJZ5scBKiP3jSh5Xg
XtbXL+c+RyLvWcSjgA0Ke7uGSs/fyuuwUHkfbIATq/WLNVPP/Psb3QEZ1Jq+NLDByu9ydbNKtxeD
RUy3v5ThALlfPYsEFiCa6QTycmU6cRHJGrq105FzyIkOmQSMsYobdDx/cYTgCKayaMlDjG1CLBaQ
oOaoq9+ybD5DMMO/OcftNDLqkxtixLpHwWZm78KRLLf7QkHwLBWgx0/B4u9udnk/rkLGm28oN75d
RocU/CkXAm6xEt5N8rfVJ/p5xmX+EO1w9Yb0YgWApXVFnldJNplV/qDJz3HISwJy0KCp8K8vB7QM
wGUjWi2prGt9gEwV5kqfc3Y67GV4NR8Nfw8jLS+ul6Nbgevvfd6lOra9HHgOT7gRSdvKRoVNq5a8
ZonbDxffaxie/mKZ2lWghR8b801ycxiLGtfxAQOj6HzA0Kl4vaAkqbllT1XykHcuHfG7aV3nLaHu
xxkuaYYBsPIVhagwI0zAbUVZ0vbNvfXGQnaEp9D7wDlea3ncpV5tv+7mSrN5Xj/FrMei46Cpyzdp
MPDZsBKlCfNauscyVLb7fOtywlPjh8pl/RJDb4WnApspz7RhuwZEOZjrVsGex3VVFeZWYEH8LQEX
4Z8giXY8kD3GxJ35DI4mlVInZ4HYBzSDCGBvORLo11Q3LNk3uSHfiJ8n77tbAzkbfD+Ujn00HBb7
tcSFh4BlU+FfqysNJUejNA2My+4c4WQAXVCGP3SQgqLt+IRiYdnnFkbbnVy70W5em32eAZoDF+u5
eNQBUypBb5ucEsWUw7T6znwnmkB7ykoBQM6g+nkzRmrppRnbLSrBFeil4rVkpr4y56f4Yl3ycJ92
igpnmanqEnDThO84OKeMcN2aKyzXb0s/qo/RbCyePoh8in0/ZU8kfOS66zP1NzyKmP1kuNOfvT6n
uyadwy0QVyeRV1bg2BTmCAIo8mSn6w+pb/52Gxk5lr6sz53dnypjYTJjC/ZvdE/knNcTS3N+w/iV
0cD3EBUBbmPtrnRxmHxv0qhFxacqjN1h+6kTXGrJwTHwRIpUMeajwn0wByZsaIbEHb3oXKfiisgB
MBzYqTakXUc5zKfRLAv3Y/sVJb2ffeCmEBtj/4dsY8uF6amPAYQ2fqSwkHhEftcpsMusO8AO6nEW
HY/g5z5NN4JOsSL6ZfivK6qqBhqahalJGiDqkNQX7bDHOU+IaW8W4T9tZwlZlIF1f15y44XMNtdI
1y/T5l2e432h2X1AMtaLw5yLdVmxCDVheOVyrsdtVVUprIERjMyhS99ggFrc/Mklx7DsUvesT57/
/+1h0a6CfK9VwWu/vmXLtPOoAy6d8gugDiaXiA59jl8WCPfgjHJu+FNQyi2LFN0sbw2qmFs+DOfy
5wJBWzQJj7VQZKM7wqFYa3IGpeqMI58D/pbtTchM6n8xYamG/NCU4ceZE+Zi1Uqnmi0rtv44ueIj
Ho0rOJJ09eUL/eXiXRkHzc1Pd1/o4qJIdp84qzDQo+oMGBcuWpjR0g3yr/LTPtKgnGa6ET1sdmeZ
h84vvVdnufa2q+fKOLjfG6fwRWruAWS2ttUqnhcezSt/jgWIpAho9XhzC5fBAlsJ8/V1UfXJDLab
lRp9kKRNNAqPZbKKz20/G45Z5zdxJnNXQ7GK4zOvXJ3EpbWkJft/9g2xgK46j3m1EamY3vIdHwvC
VLw7lQDEbZDFSo3+YEkr4uKvtUQzvRUMdSnoA9rsbcT6wFhZyuU6Gg0Gb/Hvl4Xf9efd5pBUmmnX
VjHteaEHmXSvl26ySFC1nyexhARi3zvkef6riE33PRbx+1p9QiGTGsQ5dLEdeQJhpfORDLeStsWs
Km+J5wOBZtavFzmpRfrkumWIE+wSzECRMzsQ5Y4xfu5eh4BgiXdTQHihwnXXYa1WtgYJKrYsUe8z
1tc505CiO3YovRoYO3KQU/bv2VJY078Ctytuteys7bTsOlr3U5OpVWFX4tWKftdubM8gbVi6lWKp
mIPiqDN5LwVmnjVrM9q91h5PrvwO3ywXgc2pjN9gXK21zhkeld+aiAVCIqrQ6XfYYqq3D6Tegb+e
6ZGqT+S569eb5FAGnYzb9O7ocHQQm/lyNKfhSSNCACsaTYyBP7ymF2w7aH8a+0HTfr4fiGEhft3O
tavyEc3w8tgh92TSFm/9KGve8/YzVF/il1mcKkDwGSUPT2IIywzAP85O/3/hV7THNs5fdSfcPpWq
RJRFi1pB+raqWtOgBM9Ccm/OEWTR2wp8X8VHzG/QES7tH2XoSVgA0A+LcUbAb42mZ7qT0Ap9WLuz
ExBReHSSJ59lDonIvZqZ2bmi1k3oWT1IrwTTY5x9L42AjLA7D+DEwUDKxij06WkSfZulVKfwXGa/
O6CPwzYBbTP+jABPLzXBUadURLYbLmh3N5y/qadA8LW/hv4nojIHkWYeTPH5A9ZBGSOeRqHqwdsy
7hkKcbo2xu4f1YA+jBOrhm7I+2TnRWLptc8I0+f3Q1PpHhxdFdv+5uYweEBMSctJN4D/ZT6XAybE
1qIN0npqZ2yzeP40A8rdduuOs2fqchJCUCWX9L6n7UiUsq+TZ/GlcmjbztQkOvOfLtjyXaaTiFdy
CVqnEYWMTlZBCjbE3PxeQ1zfzIsQR9zuOdBqQIGe+fFTKXsc7jgTkiTPVyt0fpPSpAHtsnojEIaq
iOpe9Jq/tSzkpQbP90U55BCPnXNU5xQq3ubZtj8Tb4njcubUy5Au9qs/74YMhOTeoySIYX+ZCT4y
3xkQ7sWtTXVC6V6a/UVtHzk+yg689Ipb9jd1kiRXPqJnXg9f6WFp3bZwNBdotngDwgvGfFMhzJCf
Ii1Zm1ZwODIkNgNFS+q9ECK4lA0o7MHpVFBxRpd2UaiNYkiG77FUDAp6fMGATgfyFVTVjT/4fCty
ruvivv+vmKoGwOPbzoykDE5onzWaIk7J+XerAFIr/Teq9TxLjHCZe62Gopx6akoZaRqS+6ctHVuA
WjNXluFa9q9T84AWSzcJVKUpcd/X4eeJhmHedOrE9M/sxxzLlCdm7rwbuQ+Xpvqrk47ZtNYJO3ZO
5HhEqLo34KwhmCcV2qpYZ1zq0+ATugOIvS1Mg1uHv0O1vsJ2zFRNyHxgiFBrWgQNnuY1uo15Bs0I
GzTnewRMQryf+3LEpeYJEC89Rm8TxCKrS/mV1fCGZT0unQtOWoMe8s49BuFXZYu/QuHmN5+vdcK4
UGTB6h2Ec1zntcenZjyPK4BkTw2GLgBLzTAuVwve2XEhR8uhKlrOF8bsQjJXO8CkihJ4frO7KSdQ
cNUzsiqtfKtCHxVnVf8k2X+o9XOWAjhe0bY8uxWGaHg8f9ER1pGXoKzjIuQDU6C8r45/ekvbpS8T
z0qyJSxfCJh1lqnLV8Mly72egU9kgOKv3dewXHnqfnFoaP9BzoAfQ5xgAV968Jo9Jf+2YmKp9m+7
KvF0buPxAUWDwc4sxid54fgP7DijVxNxvmqIVJrNx2YePJS+pIe8mQANZup5AIqx2On3Nejea1Rt
24OZA4NR7pP6ZPbXNkhXIlzDlO+K2sBXg3c081Wk60Fyo6lbsvelIA/UZ5ZGjocqEbxBbr9YUVFm
F6faYahrmnmWfqQ2lYH3mPL+NoCjicOzCp6Qh/f13xEeX1kIEzyfKwQS3DJJ7uyqgt/ZYCTR3keo
3GtwBv3IiKFIA5VKlNt2+5plaj+PveLc0qa9vvZyWf5mKkhtEUP1DBwpTCXmGYzlSP0PCbEXSQB4
X3mD2hqqDrnouIOluVvc7WgnFG0EBfBNjBB4j/dD2ztB+fMhg91H6SamD2jtwL/QkKoqNrIh1jyo
V0ioUd6lbvibtJuGOEhatvjYs0C6NwqnZkFSjLhv6vRdy3nV2aC385HXfXI7bzYIZ6S9Bnz6KbLS
QHrHKiCGczz8thjlVM0u6+T0DELStgYgymMmm6x6yNf1FJnD150D7uVleowC06znA0Hr55/6ipeb
a8Cy0IZOna8peIgd1DQUmwrXVM/YHaYJTapY0zeUZG9EIL69G7VsDsmReohaWrREPa6v7pmffHZ/
/CnLCbDTG/p+01kSCHiiO7UMRceFf2uY5kA+AKqo5Fifn6zLA3KWSGOUTL0hQ5wCoaB4yDN+Sk4C
+ICUGecgNUlVKadLHbJr2L37xyXmWoc5H3qc3G2Czw18A5aqXA1bo6SS+hccjRXk31CGFNkkYwp/
qvz+AA4je42rYqa0C8445tJ2n0kyruif0O7dHGIqdT7CHS0ORGxu7lnBCX8vjstpaHJxY3J7I4tB
nnS63WBFy4NxqjMqRzJV1Zk/ZG/IBUc1GhJjVZVmdWnPyatD3u2+RSRv4/eXTprQUa16FwQNGQbm
tdD9gFIp9DA1Xheo7tHXPtrvbZXOf/L/LJqCsqAeLfQhmYouq1k0EY/wm09EKVliu04N78CHfuPl
VDmWs1/W7CWpAG1aZMleVngAu2GWKj76EkcbBjisAXPtc++3y4MB2uSCvTBM/up6PEeqNPc90MBZ
3tfFU+dO2i4llCNYT6a7ADKtr5pcfsywRXhNP2v5jR4sasHlZ/vcFUf/eUNyh+F/iQUZUVt7xoGe
h+t+2+2s/Js5K7/LiUYJPWG9fn/IU0WLlTe0jH83YAbpKda47rWQofI6x56cl20NFGMTq23HIece
Bwq/x3HuW6paE4WKrmPIuVmLWTs7cT1hwbifS+okDuMenb4JZq2gulAGawYKb2ojS3XEJ8RMlSwz
5u2DZfT0RDEMKjWLAVEot71OlHm6F+xloTGD2mdFh8jsIC88mHljTJ/YXl1kCBfqz7t3sEe7Pu+B
79azoyBlc2EA2I//nwq2XsnxpsZ1CTX+CYVsLc47r+VqXpQp1WNPVd9TN/7FTEn4h99eGR2u33/Y
vMtQ96HHqDXL/NkioILIG81nvFBaSXieWAPK74j0CKKP8hR+gYVNt5XNHpPQJ//oxjiWREWydHSz
0gWtthKGXg0YOmdCDJ+phO+uLHUCrINa+YK2NOi/f4h3L6Y7x6smJ8VL1dI6dgYIGMhZgDIPSASy
pV/FiiS53EdGDVL2nF3F0A9juyLTacQ7sreyd7FG2M5E5iYe9J+gGTOIkHb0bih6VoKp3+BskAOd
H3tvbFSKNJPCdkCfUhxLW9QETe39Vvt+cuiquaAQZSnCMaSLo3V3EnAHWcj4ApJLkl7UwzQbA9u+
BaxB4Wt6nIJPD8YEFYMXPYfOFPOAyehqX7yyxIQmoWxdzTQexmOih76zZFVh73RzrwM/qHhjgAVA
nl4KjOKVKH+efP1Xs1Hvf8cKtAd92uMdDo9Kr6D9A/ZYoFw/mErz0w+G5pWM0nkVvNi/0LEx6cSf
UG9kgcd66Q8ijhhfhaWBhofcNHSbmv8wz2a2wFyc6L09AC7vVecLYwnQqGj+gJWuB6IRtWschdYa
fkhpR5xbCf49+CyKv4MxGYK6XLQbGn89Qln/rwamBGiDvwsc87KrofcuAP65mruBeYWDSwO0ErT/
QXLw15CSnfHQEVjrn0vE5O4yBUUmbiByxVysoW/gRhSzeEfvIMl24TXRxX6N5jLdQnv31szLUeoN
4QZz4ZepSBI/HiIFdTFkdmgnUJpIr6f2ZEhUpR40CekvL9s8BVcU9OdJxva09ZfxP80PTAnCUS4j
rSxiNFjItzS3/RBxd9MYXTDzHsmzgVIoVOJoRGPp/gKMs0YOCKY2Ocgee7Xb5Lc4v+mXC2WjTk3E
KqsnEHB6AD1LzjsdYEVqQMb/UriYfyFJ7lNXB0C0BgNzvByAlXUWm21+0q37KQzCRe11JK9/HmaV
spBaH1fDEFATWHnsKW7w2qZMoIEm42768rRXjqkEJcxnCu4GOtM8uL5ddp8Xio/j1rE3j98HKQoF
iTbGfIDNNheSp5CYwUCBjMDzND+EDPdBTXcOORUnFynU1scCUmiqJahydltPbo4+KevLv2PTRsAV
ZnDoEwjhQRYHiNEUsV+L5O33EPz6Utx6rrdJEMbesB6ycyt9Lq6cWN98o6cPVtDkI7QhWKhqjPF0
E7BAzWVaqiZ0yIFHsBEhAtCoFDv4aIi1/lgHXPQn0Rp7q340IQsZs7tjsTW8qQcqyz2TiBnLBPdI
j+mhjjMnT+kThlVCH0c+9bSzxMImt0xoEY2Md4jP2GQmuSpQ70vauBETFCyznF1XWqgLEb9WlQL2
gUdkBHf4c4rofLqA0oSfQHZSrUjQvj2DnJWiXGMPr5ZncigYvr4kojWyQbx81T7JKQMFKIHkhXxh
5B4hUcc5SB78Ts6CVh6IYi+NUx25Lq5pU+hYfE2RVhgeSX7SEdCJVEf/CQdZC7AjevNlUSMmNJrD
xecMrAC96y6N2UWXr573Aeo0ThAvplsyicoah06HuLqYSywK7q9h+zZj5qQk06xpLurcXrcic8aq
6KaDoecd4pyJvI30R5luP9nlOjWDRoV00288h85LVXV91YrhfcVXBBaFQpRFElEk4Hwrkwa0U4Lj
SqpneZ0dSu+uGWgwXEpW/wsYq4loZHlpQ7KyR82BHlRMbfN/bwfEwIEfWK/rMPgWjKrJp4RBNpxO
W67wxvloPI3u1Qc5U11nf4+X+2Z1ZKaZefhJx3SPw4MxY/xLPBrvEA7EVp8y+DuVYe47mOAvS1Tb
NzcW0VVptEzkp9JofDVUoeByT4pmxQVX0g7/144eSPI6gfU47xIT/SnWgPiHIY7zYNAf8KxWmwfp
6TPftxTn5F71y5Vibufp/KrHBaWo6EnOywHIxR1IQWuDVjiZJbZ7LyiB9s5aNRAcCgrwKAp+GfIN
fZnuztcgxNdLwm0OXxh3wM14xT6oJYo/5wsR3PNVSr+094RG5r08xa+276wIoL1ZG9izybETDn75
VOExZFJC/qJKLZMM5IImhHcjZJSqwouQfBiABZ+eTUk2tgrRWs9KCb2vY/rK0DccbQY0hYG7I/+/
gLwXVumV2I89drPMS6aE2b4sZTLdH4oYDYsA02IMbKKzKn8Vn09O4fuHuExI4euY5AKnhtFiEhvv
XM/DGzYbVq5rVkPOdLhySgmozdJe1wcthDz4d6soUmRyTno3BCTh2uQqCdwSmIjN2QGuyYFQCWkO
fefxwbehqLxZdwlgA3WH5Tn6pCFm4gClyFdbWxIyrYL/yoipsOrVmGom4oDQ3Lprzjp8sjtsjnBs
ePyRfK/iRbkfJuVmK41uLfovlo6MFvH7ZZgGbOlmL2FmhJKbiEkjY1WzfLT6qzOISMfcpPK01zSa
Q0Hf3tV6uBqZJUXzh1iWxw4qNFdFQNbxyXRD1DonVAyZJyhCtcBxiOlSOoHYDW06l4UECHNrxM63
hhntvIN6i/+d/tQkSXCRprnGOEd26bu2YCb1CAj1r9m7Gf7u24CkJryOTgWVOydYTQ32a0IV8+Bj
Ik/TFDyZ4IXrUUXKlhXMB2lXvMLXpmxntKTbxcoW96ZSEBJedr0ykVH9sBLYPM1cxwWAqZ2FoHtT
PTVGPi1xfvqj//1hrY8HoWgiNakg1yV7tiBAMmlOzaUK4wWMBIlnO1cMAMTr2WNujjdSnTrzqGtU
HBCoaXqpOjxGnaBty0jC+CwnsOGbWGl6ZW39gQ5/1r508+F9rPcqXzO/aoYUniyBHWl6jv9ssMPf
l9/fUdrhV9Z7/PG3omzxS4VTBJfHDJCBfs4Pig81yJpwHiDsQrG7mfwqde0tzHNNNLg2ObggKsRb
JcCBrDuX0WweyPCoXeuI2Q7Qr5e8EgcP2/bdbbcf09YzGh63e8lIDKDyWOyNfsrhgj8MuSBsOhoA
XPiRSAoUY3KYf7yyRdVaixnwWWzBT1sG2QGhn1gQUdhKmyVP2UffMjusmxT+Y3iVhNFYVBtJAWVr
tHOj6bDpzNizKo358kro5UhMmy3YyTcMrrOetdfmQnPAMRWGbcoHeFI8WYyZoTKYr6CW2J2buUob
MYqlhu6/MncaykTzd5s8JGid5A4XYLJJTxE5FO2gKGD0bf0/QzFZFI2c51DBgrH0jqADGemCqbvC
ppQbau869qyJFLDEvYXBOBqhkQIL77urAFh7C9wa25LMy/nMttHbo34X3/olPxKLhacO8ncvd9Oa
qsPx5AK+3+DUxyjziq2m1j3akmoMapy0DOv+ufKFUXzp5ukVtX6rLmRdBewdVImwMmyCj9AKhird
b76J1R7w5tNZvfQ+EC/0duYJBmB8dyc0zcxmv8KPi8x8QAO1wvGM/CQSmSjR7KoDXPZgGjyKZhzi
QVy7EPd76sVnkjt0Sdxz+HxHuvMt9dcJCHeZ1IdX81fV44nGV+uN1VXzVPhgCJdjw8yhqCDZrZ8k
Xf/hp0/KYLmN9DbwmSSsXlXjCo9/v3dr4MTQujwNilYWVwNDwv/E59kEXaalDxRvc82o60WZ//w6
9NY6MInqhgc7IQ8MwAIc3+0OEXjeKf5wIEDbj5CneyUmYWcRc0+LpLbKHtPXyew839TTmUcqx6uD
JYfkpQayBhbISjIUeOhSw8/DtcJ771mj698IzOTF+Q3gUzTCy4//CJXd73G/Jd4gJIDChKpS1KNt
lHprrcwdmifA1iyi4vC3kCjqcGU96KixtYsTK0pkWosegEhiJLbOMU7KW6an0pA/Gfjpw0umQT5T
MLcWkT1ilK7QPPuuRdBbSvMk27aZNDjkJjiUN/N1HgRV0jLv0aAWFD0/KFCUorypJb5VXTFH4sQn
ObX3Tfkv+sZmzZHdLbgarHJC1ZgyWQKCUAOf8lITNN0MCe+7yt4tNwSyGyO1Bu9AtMsbi+svFHvQ
ScETU3UTntL4tf6pGaByHhzN+VJh+mOf2HOjn+q0TYxLIYsuDb0QQ5iYt7kcWXVar9PeLBz5o54E
Hir/dCiilkEKTAPZJI0ZIW1G1vyQ1E7WrXoawJ67pAIY05ohK5xov6bfFVpgS9TyX2PgSZRtGKgY
lJYD3nxdGR+uF/v2CHJJaKzzW1e/HhHIi9HGWvSYywom3/kO9/eV/Ilv+PiikDRr7lFqFeyOtlG1
1P7BEuu06dAIQ3qgKGIoBzG0CAn8Tphd1e/aJ2EVMBKP33cxn63Alzap34a+EQQ5xw9JKl0BJWdx
QNrTEBi7/sk5wP2lLGbqvRpofbicIc8HdPAyLddaw2B4NkSV9Wq6KnJsNLLCUlFK56pTF9ZhjNHA
YZJ2/dfN+ORNmaTm44aqOYDiJJXwV+hKL08Tjm6Y+qxWmpKe/Knm1AC6I+9CEvafWEIrl1aKEaRw
P8BJDoIq4m9IuJGKCQdF9biWqxs37190a/CDahDyz/r86CAzxjqJpuZNn6570rI1659jPtvelhWR
B9zekWh+hqPq4Wq6tXg4NC+r3v/07dnuNdETkU8nf5DjX3BR/7TfjMMvitFoLEi/EN5LN6b5UW4G
783f6EDogSpriq5egF0TPvtOLKg6JoE61bT5M2vl0FEvl4TtFBhhnhJfnPPqR/Fj4cG8ylGmHlqq
Sd8ZimTSEGNeszDyxh21NO+aSprpltodQdr59Oxr96QtdQdA35cbFKkHz/unqkuWquRkROFeZ4kE
cRp0qGap1r54Z1zVX1W9QQmj1RMfi6zp4Z7amCRVkqgMUdV2XCdehAvR6oVZyYDBS5nVD1RSBTp8
9GUEK9EJmbR6m4MgBVoJJVT+lIlfbpGG2/ovVh21/0d2SznbyEeHENyhQC+Z4gzJ1EHcby/woai5
Y30ZPpwVvjbeUC+BtGJIIqcf4UEM+/cSlqU7jBF5I5s6T0KnBgAp/l4Ke+LOtymEmrgmtY40P1xD
Y7U82+GR185+XVkfIEe0ToLuWaikDdOT8pucp/scOxnTUrZV+8pOtxHgkTbQJMfFIVcKvb4RfUjo
lwT+rnieB8gdYqhHAbZZ5J6lP8AzA3jAD5QS10Lxs7k3W04KS6BA22FBXtHJdngBWA4We0yyHFo5
oy7inmvtXnyYhBNDY3KVhF1mM9xfMk4Hv4Cx+22ukzbdUPL+dyNWNjL4r7ScCnrf0RU1qq1P7KCl
v3Tv8o+HrS7ZMy2hmUvnC22iYIlgQnLjS8V9uD1pbj7U+UEm2EcZ+r7pMqQ0UYAZhvJ/VdgY/S98
064ujIjghaOHlfkkl/0DpkTEUVpZsAZjaGp17P8h3FjyO7Aw3eVVqbUvGtNPlUUFYf6SQHh3mA0W
kfDQ7krMsjW96gesqGbysT7pqv1wBechucC5onmHRJV5q85s5a0c6oEb4y5q6WSCh7htc+aaSNWX
NPfZ9zSeJmwwhi7mK97jNYaThBXhEjsaO5byfgiYtbMx8rDREGhIlKkvlOESI4uFCrhLnnz6HWYy
QMHy4RmzL/UmigAEyLEa/ofOa5dfwQZjifhRvU041LLR0uvhiSEc9rAoTu4uTr/5ce1avsgmeNQU
K5GWepwHoCCHBlTqrEIvHWyw+5g+359Lc2s/7XWa1k7snVfpL00gaLukfbPZJFOkdZPkXqMcmnb3
Odhv0rYFEkUlUfHt6vKjpPtxDyd+OwBAekThvNBurfVMh5SOLjdg83EjIlrijKTL0csxccXna/Ue
CYSsatXKHh6Fd72+6QCZxDmRGXRGsrhPF/d1ye6jBqyP34p20k9C+4JGvxZS2bZf8/T9R5YHys+D
gzV6P1kvV7vrO/Zm13DKgFpeT/5mMFsv/t5BvxyfJMaxjJkQflpUWh61PQjMz62AR9AD7aUiTnkR
4cFtsfogCUa1siro/BxxnoZpxcBKcVL3e/6O+T0oP0OWLrTuKYOUFFUzQ56iqrgXX/K5B3TE3XU1
AS7iU/z7qZT6yWSshpH8s74APQiUKfoSnQAPscfDBcPlQT5CfFKXIQzTdsMSLYATVDOGL0uqtuJO
WnZxBFLLyfJa78huUS3mslbAmsxAUwtrJvnJAq3EqOXY6p60s8vBOQLs7sm+dQKd4LjqqMRDUZkL
MsywANqTcioo/dX9OynOHU6Mqj/oMaSlPMf3OlQJ/HURa48IpJ63y8fTbgIydA726fknZ/EshaXj
CvYDTJvJoQ8EiYjUIekuBLjYDQLvimnlNRAruOYK23b8G+OQAfAAjQ6RWw23M6a5b6qvAg9BeHiW
Ei2a+ZSwfmYEfJi0Tg8M0vcy1C2JCCE+D9ku+tEjHhgJG6RRcK1CBgFVazKHKcvxsnagMu5QhC9F
Dyg8quwAtXFC2zVsAh20rcUSCmEmORqAVBhwKHRWXr9kw8TLLw8/kLJH4XLwUZBSjgQnEbRvgYgl
+37QaoFmHB6ts66SB00KdYhMHuh8jLecVmr0mvUNF9FtdrzqvF0gWISLNbkhXdlybO7uLhs8xKxN
1g2fd6+SwwB2pH6y+cB9SnRo6H0n0XAdRQujK/Ea3wNmX//jEhOJQgb1Uig+XChVR6VHz9o2jE0E
f80DId+ceXDXhZ+4xyOhujP3IG9evGbijdV7UlNZMc6n2cIgUP5WZdGj2DkpypT+lMAKb6je9vYM
wT63d/j056XKDaDlJ6K7atW7MLcM6j66YjuHRjmsQK6H1o19cFdesAZSE0KfYMpackgywpAIbw3L
jFYpBq0EiV3iLOoj9dhKKp87inY1wOs0B7aTfQK/H7AKC35YZg09/c/9HVU8FdnrLQlZzdvjkomv
NofCLuiIbZFQkcWkt1xDVX7j3IYT3qeiZ/+bQZoDZaJk7BODi6kUMD8yPm/rs/KpmcA6OJcj6L0C
71Eyua3KMycsOAClWkf2hmb9/XN/WwtPOoF856TD0ZoI5QPcc22NzQGpanA6wzTKbUk67g+5pqNN
8H6/zG+Zsfn6ca576oKlso8fLHwFz9IIcb6YGRaU2Y5BJGAD9XOjf0F8dst8Yje83Ph+5Fr6P5mw
iHtFJENpjRj4xzNXj/SB59Qn9cV+E+ZljLI+24r2UkWokFvaPxlhuyWxu0zEPF/g5oNUwnEsKiXF
KXXCbyKTG5EJDyGByEtpMqUzz3JaRM/Liqkbpr3wIxAKdkpZToJDzzWhX4wIvFcHbtI1R7LECOJI
pMW2QPIrkrD1Mda0vbqBj4vQ/LZ9QbBBqJrOHcfkFo1lehpeskDJInxqtmqnFHP7+tWNmjT36t8I
eG63avfd9oAkYm22FgQG2vZ1kAGCHRDt6Nlw33YmskDT8zakvnpycFimysi951avgFKHZGSiJS1S
Nt3ELO5a+Q/b6bHaga1Dc9jvr6DFfo3fw5jO9I8RHPVBrQ3bNU9fD4E2LtusHDu+avHIjP1L92Sb
P4zGXxuGFaZXjWCAna4BcuMQ5AF6MYqKSfTLesnibM03OL6eHuhKKTQ3CqezEjIX2QxyaqqFjrt/
i6lQJF8jxKIkvDh95PbtQErWUw+6nOYcrBcdjS1aVCaCQvyqdaITGrUJxyO1ns8FrF/lHlDuX8M0
U1ZNsC+ToBznJLFkOOnpUsfFXgNJjnTMlNiytMllAghBAykK7rJ3SEBIkYfFeeEYyeErm/Uzh6Ij
wVjHDGb0eI7NWGLI559Zj7+VDtrVQcuXivtiJrOf84bfFTkZ9i01xO5v+WKJD2H7fU8eyZcxTdcT
WkVxcZeQ+yi1RYRCgNe6ZpYgiiqieI9wRNSCWd/kLWSlxyF7ojgsGt/OxfqWXYNEYYuUxdreTlY+
4JxTpEUmmWhRn6SuQ28kUHW09koel10SYjrOZH5/Of9MCwzkvtcT2GidWvcc6gHucBZKDEHSHmko
SJ8r5+5+gyMUpqAp+j9V7yfB3Zl7E0232vgWKJFylx+9q5WrU1+IZwshEjdSfD2dsQf/skpYHkgG
rRR7GnSEgia7ZwOSYB534LhEC4tQXJOX9ceFrBmeP0Q6AbbfcWBf42V0fwEbg7oS26cDHaSk9lM5
265tWu1KCk55Zde22mMKHJ2S8wIKjWokLnpe0udz2FNAuaGMnD9IQOirnDa0usowAstkABaCnw6X
6rYMDdiL/kQKl3YRXj/Cb6mIEaf/Vgghafi3mgrQcs3cx5kPGGzfCFcfWzt3TUyobB61ZHD+WVgG
Za3QwTLo9L6dyH7dWr+lReoTh1WDH9LxbGlBTap62grCPgWdcZirBk9L24ClwoT54q7KZg/Z0Rpp
qKjiDZ9bJsbuIudtWJ72XyDu2t+BkXJp095VNwjkbiBs4KbMOYmxvCl1iPDD+vhDTd+l2cCCXhdR
ArOIqhP141TbTpzf5XjHd3zVlMzM0159Nrm+gpf3vg0u+1051YKtU2O2btz2euejFuQwtdFTRsOY
osuH7YhaWq/KY250ezncVS9I7mnn8IqW7RDMPrQeE4aRmdwONrzBxiQ2BVFCu2n9qJKTcVNMGvj4
dtlWhWsESt6wDFfdbwOs6XOgsRtXntsrRBa8+Qqf6c8gKI2kLoS7JrqZbhWMZxnYbQkH5nNe00QR
cWVmc8hVWKS3Rm/OhgJJU4qzu+Wmp+duXOea9uR6b+0geqcyK7uz2fg58mbLqPZ4uljEgRLBuIzY
x9kuD3JKrzX2F+zTYjxYMpgD1dMbfCz6HNmjxCYXCZ5Q2l19CZhieOOmacHWwcNYCBhLv/VYnjKx
y8u1QgA+6/W93NrpZ4xxa+jHsybM6OcDLpGfwGAw7c9iGnlSNmETrb/a15YeY597R6fyto1ueCMp
5MgOjrIHbZ6HmZ+91ebSaw4Kcfuu2ZxDm34aTkn31DLYo9eptyjgrlodYqH2nQlBhM8xldXOU0Ip
ClWgO0bskvVoqqbpqwyCi5NegswClz3sw5z6KjT90UJ9RtIKXzpU2XZ8xq8RE1BaygsNVFpKueM1
IKzu5zb/ZxYjslBSPuJA0FPtn22aKyRS4ZZnc9YvgUZTOC/mhWKgDRvURpuax45mam9VKzkhaApX
qGjJYXF94drQSXcbAnZOTjKnsZzhBnnjqxkP0AcaH33Sw+dHffqbrxaEuqo7Dz8bYi72bRPJ7mrX
jOYCVjmYKrp/t54q9QUtithbb+WgjuoI3qMn6ytR2kr1ix7OnjqGC+NRdv9lKqbrJzo/eIIfkTIe
1cLR/9WGLkGT1dWd5ra84v6kz3XeTHW7YYZDFvcfo/sotHajmydTwzsyP3Oh2e5SnXhZr4QO51y7
iykDvbLDIgkyfHbibMVrUlLOiGBdJMIYeoE9brnouXNwR50CZIw513UGQzS4ix0lAJsWIb/628dV
WdzKJAG0euutTap0b2FQz+FXt6g6OVW4OjZbGt9TosPtCcxASfvcXOwV+K5Wc0zSC02+oN6x5VrY
FddPeuK76Gvi/rNHhbpYgcSLZdKKBSv2xsRMjwKADUwu/ue4c/vfidVhuCxWUZLDyVBfrBjiTjqO
O/tJE9mDJgvYdxspf4oiPL1Qz2Jh+BSNJ0WC4xI5zOA/HRZjUxln3iXh3S/0LuzmWVCKZnbexFCg
L/ZcKnFCwCN5Co2ArqtVIIbb0OiVyUUTfUeSgF4lazrAgtTkztYCQT+9yLAH6JO1oXLYAd8ORB2b
Zq+ELTOapu2FUZizOoCbXzn9mYAt8j52nHMvR/p4+EHlpZfptesRHJ8JQ9QKzHqtqLriUlnEx/3f
mZeHeiZbbeLTy/Ndn3BgkjEJ7Lxb3t72gPZ4017/26UWTtIiLgmcDahH9KznnQMGOoZy/9uP2Nfe
3gUFgnPFaflj2HrWDZkgklp04QOSVolkklj7FRWW1Ij+OYU1YynDkjbknkPEQ+R+174gnHQ1fzFY
2BLG3sUexpfdv7xX8Qfau6DKaRmYJqzb8/GTdBaLPObFlQlnM5JUDe9SDaGlmw0fcL9KfFxUjjBL
Uolq35EKw+ewO2BQZbiBuvLi+ipqRlRJBkQ/6Rx2bOpGrOOQRVdhSIw41BpO6TBBjP6d3YRsHdwM
wvBPh++zSSMdvRLN6DDLHUlB+9OeP8tf7aarJUD9tBXuFhAGEsA0r0j5kZ2nvbOHJ9I1wseuVXSW
FVrDsUG7UFA814NI21UrDUkQEylAYxTyJ+e/Tuf9cnlO/nzZ+R7hOVcfx+LdDnynmi0iwHlSqy69
mYolgZZO2XXWPKwiNTLDgUhNlelu0bMPaP5yq8YBSIly3BoQ8GokyOuPm6xUFpA83BC0N38fQ8nC
383dybRpsXPtdxODdXjfXI8E84XkV4B6VY9TYxSocRqH4fFjZx7RIUxEVvd2a64TM7GM85yeBqHi
A/UYmlWCqlkAnH8Q7lm/rtwi/mD792bF6OwF8FwunSTBE9FtKf/kdngo2uIwqhmriQJAPZb3/kPB
2Jov74cA7WW/uXAZ4k4NMmuqCQWMxBI+u6BrAAJC8IhvcTYGX+mnMDpFXcEyxCTODFb6zJUHWzyP
xlog22aB58gzqzVxMqO8HlSZMUOiIoiAiWOTMTTgU2zvMfRmzD5a7EC08cpL7x1MSRKxEcPXy7r0
KWtmpc25GNtVM9nUhQt6zlHQTUQE587C/YxTfuFSno165q9Qz94a1axxW1ja5t5NNV+/SCPXnhx3
D9ge8WFwVBMhb+9KAbuYltxyOrpQoCMjbmiPJiJpVG9YLwpZGY4P+ghIX+fGd7W5I+sphnKyIfhT
uBsVbi9OF7HJuvYC+p5JuZ8hhWNNW2aRF9zShbsvNLykuG42K8jzQcGixBY8N1kiC3kes039DRjO
eD233CWQkBxjJA67vZUPNkXULFrEoADLltaZhMl1EF7wrr3hCbPzxwK5hVBIXF07YTrsLMT+n3ak
vGWd4Hi/QRuJv4PHxmjaoyyXleiwuX6lC0Bd05yRW7wJ3i5yqVpdQ1HlMigm9RuA083hdTLmdL1M
MqybjFCJ/bz74wSi0YdmV3MOPGvb7mDqSgZSJefsNK6JXvL26qNGkqeCvGybSDHdb3CGx0RkRmtd
Tf5CpWneiDt7PELMC/KLUPF09eGvyL4+o3O4Rma/hZ5gMJTGjLil9uNCx+eaZa45Kv4JIrlCeZ0n
4TMSXUgtmVLRucK7V9XA9oHID5xOb7I5UglMpzexXuD0JyXEqWHpBgc2LkUP9sX226QT22Ojytcq
Kp4t9LL2Y15TTiytoX1eiO+J6oLSLNer9mIE/TYWoGvcHSHcIi9veyLjyFJ/O1RCCTpd2XeHAm/o
y6Iq3qGeQJYal8WXkAzJc+z2AEo/Ly5Lxbxhj1SOP/+SIH1qcRqVOsY0nnaHJr/69LtApi9Udpvu
yb66Jr6fSZaaFG2jIlVnclwKEDKcNmSnD/smpXIj1Paq4HFs/TRh+Ue3Alqe+w+hTKsXjuojUuwc
u32F7eHqfrJT3FAWMrnJXDslWsiY6Kp/r15HPMSiCOuEwPgy07Pvu0gg7I6l4+BpbC+yM9E7h5Yf
MvLyDyOUU7mZ+zc7lwKJcrI/B+eNheVu04fA/ML+NLytHY/ZcHH3ECub55OaOqOZSWiUCkwnuWU+
B0cRs6QWo+n/oQujjB8h/DRuDan666/L/ywoJci+02qIHuPUd3VP4nhWSaI2Xk6eYEDchymrdaS1
cTH/wTrJPOQ8waQjD3ezTWuqL4D8BE2KeNLk5dMp9J0O1Elrlla2mWJ9r1Xvjpkk5SpB3DZdBOxO
NCWJhEZ+JTiKTbmUBS3T8gTL02YOg6QdjyeMjewBn0KLtm4jW/1wwoypquGxXKJtew6/nDfj/be1
NSRCaN/Gi4xFmEwBA6lEPT+X+VEhQ1XjAoiosS67FVxI7WyW5Lpl+rbfPDuUGFNcuwvBTdOyKYRI
fhccU3ktPXXJZSrqjP40IoNNF6+e7S6e2dvLgCj00+xZADdi0XV2usI+B/vM4E/ljIShkpSbqZSW
z+HY6gUJSUPHg9D4nc6WlQzKQv44lVaHsXIQGHrNyOKZFexfy0GT48GLEYT+Ic5aM4337KhTyfDZ
tqQRXeLQuyf+j0Cmp73hUdQ6Ht5H4bP+c3aKp2LWwzyM5foz2SktBxgOcGp2j/Z3fFYp/8Z6pJKg
aRmGqv80vZcTdCmFOdZ1BYUfSNm/wckE56ZnBFSXJ7iKtrc5ENBDdM2e0+yFOvG+o2dtFEjfqM+W
G2Ktgn/toO2/ltsr7mQZulLx1i/WpKK9wo5QUCYxpRLZJp+R4tuRtbOsOGhyAVPI2qC0DhzGeBNH
2E0jod99tlyGc2gCJ0OpBsYFUAIrMJTw4TB3mr+IGnhKz62h/0x1CTBLl04JHqzeNjhcL69qX/C2
ZVgI3g1DEvSjhHZTUWZb7sZVAGtojMXPWI9guvFutdC9hC5w0sFdrYBzl43IVL84BqDpQtZjZSqi
FTVGn9Ti+eVGmG34uxJ9w2TUZ69Fd5aW6y0x3pLGaoivQONiylyXP4Slxs5LrFqSuHuZqKbOSabc
03er39ICTTPdss4P3gkom6wXeOI7iFcZj80qYVhkK1SQQ3boSO1mwQZ9sz66kE8MEow96fVUunv+
8FlGawJY/8eutlgjXSSWR2sSay1FOpQT7dQ7kl6Yc/q0j9MT2n2K22OrgN0MON2Hh771nIRpnJAg
DXMfH71lps9YSf0XcjvSsGGfUXUCgkilzpvp86hSYATL4PRPryifoi3MpzZfpQSLKZxR2dRA2nrW
3gZhVXs3bLRfygZpwggeZZBBDSngJfxuMXuaT2d5TQLqQBh3A9mP8YZNA1LeyCy1xQ+XnGahEZNw
vbi7VM4BDq+0nMtr8iXfxYbAKad6f4fhSnPwKPj5a1Ef4Of7H+cgjuluD3tdDpb2nY5Mn76kIh4v
B/2G+o0o05I2HavuyPio9qtR9isFbw2PRhwe4m/OVI/E/89GhKZFV68GjUhCN/3Kz9XpydaAeL+4
Ts6X/j8fdBnKrTkLdXgcm0CLTg4xX885wRCIYNaB7YsCyZMGgD4X+SOqgVAH5gs7KW0Z70UmT9tj
sKmmP/TQbQVTJwdOFQ4zfFa/Xp1/R+BQ0OIokBcy95jYPrYdj/fNbTLTMlzzVDAuefPlOuUPiSXY
8gSlPeuQi05ASxnqrS92FBw6/W3xEDpeey6zXJ1cN9i5HNWMlHyZfNjlpdnGJR9xkcBn620Z88xo
X7sK/hWjhbk/P2EK+52+E4bIvAollUAHsPWmdr5eybHMVaUTqPGuZk38iqhPsM9QWLLnKS0mEi2A
/PM/Es8CmBVmVfHBUb8lAzZkuQfOZbeWJlK23YFHXOPWkjiWKzudgVRTJiHlQYJcKXSVtdxjgXFj
TfHDjTuQETynIExBSGebx0H/dn2n50/Bn+FqDF2TU84DhlXzwc+rScg1lQvpm4Wm1IZ+GltLhf2k
ZzqS+zz1NRCDNuvoBbQq/yH0wjnK/U76DM/90VvQowqx7VppJ50OwqSuLLoIAqVfp+g3gdlELJQK
ZbEgACp8zG91tGKQVL6EkIoYGAq2tTSPQ9T47Pvx0blyiEFGv3FVmpi7iq/oe55TPUkLmVGmSM2I
VAB5vi6h55bLZPcFdGRW8xrF0SERaH4dqW9Tl9CakFq+dqFtjpdtfn8xzxSwlid2bJxRNaLGE4AL
f9GPUXgPGAtAZmwohI79WcfqbievHLnewMNOD4V1j7TeFnMI64YCRY//+qtPPaiVkxbQWJTo56NF
3CwTWiAQZEy4YQT3ie9NMQy5aAig/38KefeJuaCgVc2uReHxS79XYbV1nHNp8Pk3+4MVORf90nmG
brpWUMDxg/eWbGYlyhKc+Nw7UDVW6f1eReuX1T4m2s3bIb7cfjTrDcNQaoFMMNeUqTgPuSFQeUzL
bYlq5+iIYNfv01fWWGQmi5LFaG7YwRrfJ9CmhQnBH7Gw1u2E+5pRyUIRJFYVFHkyQMHe+Wr51dYc
rHMGtzqBoG5xKPnVL66q9NDEfJSa9V3vqxheQNUullHtwCePhGlcDzYIZDFRcBb9mAyeB2VpZZE3
+H/Xf0KLkV49Ub7tloxeMLJDAO0HtPgRmib+AqT8AtAUEu+ILuOol4gahMXMA+kHOKPK1nfwkawt
RronefpKchTYB/W5Z8M8e8s6Oh8fojfNlemuLD/BHGJ3KcCb8NvRjpTv85O1th0LzYX64heHxA2K
CODluz0k3vnDXcLpIHnSzzI+w5yXchSMshSW3vMJcgBPZKQVxdvMSdZjOv00PLwgoI2R2V6GRlXC
arNhYoiviD57Fq8xgxvDwcMlRfhEleSga1Sv6x0TfPNwIjXzbljCg9O+UVrJvIwfiAVGG6kN3+xN
P5omiC2PfmGRRmVR2IlciUoQkIiq//Do2ZdQQuAahZmdFKxtHbYwrb0GipVnyBkBB2xVM7ZtYmJ4
86GmQVpMOqFtkpPCv1yGYUA5Sod3OZJoOQ2HHHLejsRDswhLSuEdrFiSb1lvoyS3U9yT+qAIJjkd
W893yavi8wtOJ+yAyvz8ZreRmejiyBjndl9Zs7cXipDueR5s/wUVZ29aytvaKkpXWVK7zsA5rAqZ
XASannVNED0U2Nvj+RWUs+7xnjR5Gs4vOpcI796pCooyc8WvD+Ed4qAT590jpQmae+2LYTvAQaVN
Tib+swagjwx4GfgynwrbcD6tKoMuoJ4HbH6BNiOBA0r8SWbU/0wK7MWnnuLnejsv98i6cYZCqmdL
g9yQCverQ3HSl0UXhXk5yHEpnyVJ5WenM8YLJ1IRcNOvE6XxfCtSNix1BKMKBQWmFYl/TbdIB8gr
KM57PSzDfbgm5RWNxls2LZBNuDaDKE4RsfNXFSAAiuJmykBL1J2YloHioI4+xsILp5BhBGRH5inK
JVohnp9dRDUGhLjtACzBHa+jSTKp0Papc1mtSyl+Q3JT31tCp5xZS06cskxecw3UaK9Bhz8wiOMX
hAT7XgGph+0/8/3/uuGpuUgZBPVsIo9bCHsSg8Lpaaf4+1EsQ8tg5VwE1QaVKGx3Ytl1tORgfXjO
zT5fhvhEKHEyhbWA5XS4h7rfv9/jzgaoImquHYNgIgoBGviy8JSORmCE/Iwk9ghavWM4wlb1kZJW
hu0LaBM0gprHkNUhP591NcbawlYkUYMtdtzhOFIHPwAlb7t2kTWN9CC6WReAaxkrwoXMyOPDQPb+
g7KxahGc2F3BfJYUKA7yzsoU3Z23v237YHmvYd7gD1bt99UlLIhT68oA5NS0FepNXBKhAFIt1B/x
O14NnqamTBpVTt5Aa9CafN3FfPgSAf1VM82dLfr8a+fRqjSwPaB65rymwFd/Wscl7gz6xdPeXuuH
5xTLXeETQUvlUcoxhylOcfOMY5PDRvejJCbPRAqjh6zo4VlQaDrrWfPpEOi0Vsn71Fkx3b55GoBR
Qo+fshZMlx++IWtfrBQ9WIMxAsEWYIPXCaCy8Tc7xB8Wv9geL6UYxCEL5XZFzmb+RZn7540cyzsk
cVssseu2mZyjwWZF1m35uDLuB5zFFYpK5cizPDYELychUMKIKwnDBYWvox1U4cFwZYHo1kUhTbnh
wQbGLmnOU8q2nhCm8KT67jvoG/comKVWdef9pV4+QQRlUgQryNfqoZ8+tNyGjcF6tfyuJbyUD0nM
KQJfyPAfpXCunbzlld8mejtWICC4RP1TuUBtQNo6ZfN0uLBhvk/2POMwsR5sXxa1YAuWwUoUODM9
tQbHNyKxuxxCcBveUiyEsxQeSWm4YgVc+fAFN1laRLEQCBdspiymTBA3MQLn30gQVGymnTt5N9IJ
pFFarXDO62BmJUclbNz2oV8UgRNYI9JPKKkdr4JYRWPglG91//XoqZ9UEHeg/a2h52sqow6VLBaI
XLb0axZYSJYlqJcwXiwtM43dXCv7BidXDOJ5jlKUjr1m3Ad9KmSmwqBEJgEDpSAX91E24votpxBC
EMHLKVx/sarEdLFPagV0pgtps+hr5JmOmxUz2tP88hRiO3BFYMzNapfBhYTFW3C64upyi1p1phQd
HU7wbVtuQqkcL/GkK2AGCD98zhI1lnRFfuK+R76GzLHFAp8DiEW9sal4x7WZDpWh9w/0N8OEhPTd
t2cdrVlrWnfwXj5jw8biJqF2KzcHzIayb6VUdIduO4gMiGQOpeZaMO7cwgM39mXPY3ADmb/BmlkS
LWYYbMWoYEyvSUtPcmSDHVhce159SITaZZaRZPAzVU64kdFgJrReuydTpF7fes310B9SWt+xCGGQ
bQib70/tNXMRavRpr7iIkanaoPZDDKUj2A6gVdUlOBfSktGPOB8rlkD/ySc2ZUxoRXs1/sLA2J9a
CE5NcTgGz1lgFrmDPVf28KaJbyOyIREV/GMWd4EGxyIyGWNazkn54w+M/Hnwgkha2qhkb3fTffzI
Fu458yd16aIVAoeYulYasQ+acdq4wmmuV2iStmYxTGbHNMkPRJpO1ITw+Qx8KRxrN2nFbuwcPmR8
Lyg357Ff3Q8zqfwRosEbwiBWzDgkfgPKAqray5tWt4sW+4LvnM49qBaaeNKsqvvMBPV6jFrUPKUj
0Rd55ZM+IWKiwMcPr7EKdaXaTis+VNEVN2FIMB7w3Jdn7sNMJAnnwEfiqEa9CJyfZHC+6ofk3XBs
NZT1tEuwuo9amfmUKvuo2U6duJgYYuEcb1EL1Ek4nCf2OsuidTKkKFg9ngQZ1U1iix0d9RGoQAuR
iSoP12/u1N8jGIUIkTClMP7WrorysViZAnZQFTCarLcG1x6zZI4Nh3fYpDBYxl6wRriiOEkKX0u8
jdhAZZUX5RwENnCj/XwJi8/knNYbYSVPXHJnJA067Mu+efc2r07FUhZV5f96+7FE9HA/6GZZ8DZs
7lXCrhZcm5ub57puNHfRth4DaI/ZxHB7YSbMo0XiABVOeLzYCQhy5l2RP96sLtn9RE+jnDFSyDew
zcDYRGQigbktlNH3YdhxqpX5ioLpMCSiHDDWNf+b4fQ6tuBDtAHoDieuvHb2c64mIp6BNLwydJv3
okrMBAkvaSEjb7db2e0zQ0NXCNGLdZKS9djF2uGhU1TIUDPVclMkt8YXGbkN+D8b3ddV5OymZhnl
sa1K7rVCEJ6fdhkRSB3TQ5JEBCuzHDj7XVwTdgGGqOBN5b0l0vnkJqU5+/UHmUxbXDbq7pnaKgw/
mhC4XugAdhjtQr8hkz7LI90jJJBYFTX/dj5EWBL93dWxOnD6ycP5pXVDY7NNGXycP7KqBRJ/xvJf
MQC+1H1/URvceycLECBmGGdCmLPWMztMqgrpWHVkFl6f9vYWFSvWIFwNsYZonVGNV8WS4ULaNnJL
+lODl75+cowhu9e7m/oJOzWy1mda9v6s62eGHUYzcOksQePGMz3G3pf60TYZqTg1mBj3uGZ1vG10
nBjSlH2TnqA29YWlW5ShUBYQksAd3LIUKReWYsegHi2Ea4/1IIlLA0upUNIwAyr6ERJlLitstjLR
K2E7CjhiF6FdN3ypBN08PzPi65GqQ0/Q3X0jmegQIHGXxhzrcMT8rVswt1DoYPLQliQygV+LYkg8
NSyxP8J8GnrLx61ERecizCAxUyLcwF2MWsOG81brR5D8EHLKT6/mWiueSrfBfTmkUg80p/OHjZZ1
0QPevP6zVVHATRkUw35oLIP+Jg+PWmd7X6nkiHRsdZOAYz3z3NCaX0ltrsn+S8CwewY//rkvGEB2
OJnAfYdrDEUFaTyb4n9Bv96ZFBxlQFC2+79i4vEIxhF80k2dS727h2zOcH+f4LuOotK9kJYlGybS
sVSCOXcpv1t5Oc+3vk/2/+M3LAxIm/KiJ687iIaoQY4A3zoMpKIeeb6tBm7ipaYLjVTtghRhcAg1
FYuIw9mIr499/2x7qNGTy73L4jhNU+a5jLk5N//kD9x9iDrrhe4EuA956po21RTztogbUa5vjpLR
bMAXNS8b1LUYJ+FkpVwS+r+PJCzKgD7z4WzlJ5xxx2yEP21cPyn9uQqBDpqQO13Xp9EmRyYsXI4l
ow9fjZNVsWjl9E0kDodjhwNZ/wwYMs9irDAoP0+pEEQHzIfIlpdDa00g1ahjZ/XNec+q/STRWMIE
GCSeBk4tBzwViWD4IxJhc6mzBf1wz5qHtHo1s7zXDTn6CoHmvpMFUEtRi58YD1xflr8mZrtwKZlW
vxnrfEMzOfZ1hZ3b2A9rG8slUmcL+WkxDG7emhIajmchC9ihn53vXK8LP5gLFTZepdqPYR0Xly9b
rpqRbLibmWK7GLSWEdsy+oLyGSIcvNqFhpWsvqQnXmfrc4nfb+nPacXlQ+fwZpHRf6wTejssIggt
wHNv7ufpDxQsZfu6CFmwm6DWKdyGRZmAR47UOc43WuQwpmjlOU2eC4zn95PYNJDCVoGlUFzMhyNI
oUiDruCvJC3ZzXNiE1+CJFHYCY3L33/a8GkVUWL7uvX9DT41W9c1fPHvSEWNuyMHiS9MsS9qEu8v
OSBQWTd95wJ6w47iis721wdDvc/dNypiZXr3+reO1cwVgJQZBGow/pfYe7vVMM6zfCjXxmYxhjfK
UsFxEjSOH7hp5qtONT330L5V8gpvjWDtZfdVpP9GwCGenX64E2+I/Xh3+5NksxQXbhZRQjr2uH9m
ULxeoMTc+STP0zynN6GkMIjhMZbgg9nDMYm8d0VIc6/zoqxTdoaUdiqZpttXnti/g8wsMaqPghJr
pI4DSt2eqiVQtDEmTG4lOhKfbE7kwk3NYBDvpgU7IlNFrEyvtEdaBNtT/oWoT59Yoj04iSbRZDt7
kiSXV6t54b9uEu6fjHZkPHGYtrFzmUmNruGeqVYjSjN4RFBksCTnkFP1JitbnZGLgfjqGo4x2k43
b0groEhfNyIp3xHLVVs9x5Px64fnLSuhqsXE7BoHuv+tILWrfSrZxUiTJjuo6K7mwKzbxJCsIN/a
+syt2fzSqMxJAfCq1uJq8paXwUDaQdaiXSOYsSsuieAa2chuh7qhFSW9Fq3+Jco1+b0nKIbxnwao
7x1VY4AygX8OKnfT4L69a8MzOelrOWrZwpyt2nMQfp7MIZbGNWMvusMFJPIMGJxhqCcwAN9jLg/H
Q3BSi+oClCpASStdTFqu6X1eCL5p7hwAwL6iJCF4mi7V6BQL39GrddP2SgpWD03sMHKE7dZR2oXY
c/UHghHDtOQAunOGE39CmY3GYR+kAe+N8g8dMlk4zs10a+CC1oumTXwm9oDpSb5kkvKSCty4i74+
4zoyhaN5+uX9NwX6YZHhlPagl+boTa12fccgeXY/zDgugesbfRuHgc0B9quDlDYQvPl7rC849zY0
QdpXMQPGZKz7CCTikCDEYqhoBl79oruAEqdtO+cAjrRB/dSRBVJFvglq9P3N4nSbUqu+ku+fzl6e
XMTBrABT5NEfOHq2GuULDlwCrsIDDNPi11CNHGwbUUHPbTwZrGdUqRgHBAjLh9ZL3cgaP+bYO3YV
L1ElEH+VDaknsLUp1Iwd/b2YvxuEABYUM47nXL4niDjSlwUiFijlRL0o8oDbV1ZehRTweAps3RzB
/RNqrzE6YfMyBBxC/I3nVs4D3NatstXxGursS0JODIDtNSbN4Zr43Ckpu0nnbzwhq30+zJhhQl2L
C6YSCI4E3aKmUy2s4SFLCWOg6QbIEuWwgyCex56k6QWRZZW4wLO4SD+mSt7yjim+u0NepC94d+uq
DejtoGZdZWw4ojpcj9/2AcgXWhZDHwmEpLeNu4oog9PVAXt7PYOMwvfvIGUQ0zDapT8WfJUpxMjw
6bWnCgqLdQRwFCFZwaIWehcsuJiWairXi8oR4ToufOH2nvW/gOvnw+7rWCfoC0dS0lWySs+TXJHj
LAQNYRwa9/yLhh2oGF0Y5Q31wGV6g9nUyI6BGx0u26VA+ytAug7sTyf1aajZrYpV0b7hWU2sTwFL
YbdCz/+TlctFJm+BoNSo8WVTf0vrq+wvYvqJQTeteGcatnzXmV2Zny6P/yMpWPrFF8zS8RwWdAVt
E1qglRZwY8hid7TFVyvwnKy1pwAP56x42DAbn47MaozMmXa4H3o+oTE6DKE9blHxavPuS9+Ozr7u
nnkL2sQ0FfktdhdxlMmpbyKS6FK8Jtc1Htxtp0KIdYypWbC6NRKRp/OXnIWheyoqnbI6ZNX50T64
8FhZoBAHjsg504l8he6P3c9eT0FaNMvSB1kKFMuaB0TpzVTTElpLQ0SWPQaTWWKN0IxN+3FCEczq
IkiLlsTHra2v3H22xtjttOdSLFwmpKRCstdPCauu9xwMgxGc4Up1rtwFz7MZrC1FXvAh6U/RWJIv
3CSjJZ6fk914asK650JA5dhamYlDJsmIbpgp91iB3EX896PJzRp1h3TkIq6zYYSpzg7rqh3dp2iv
PbVj8EV1WW/DmRdpZs6kldaPqYtVrX0Tu6LGcRqxXmOWEdl2uVENJxM7JddCc5+N7LJCGNjg1bcf
0Omlg2EH/1dkkfHe4xz6M18DpmwCVEa8AIRJrJPvaIOQ03s8Ab/TqDWrh1QOdmTcwc08/spxRSKV
re1OD+ORZsBbjp7SHvwEJ9oSIbsY2uvkFfQPJgPRKizw6ECF9GXk3RVeArPyqvFkGzTlxBCoHRhK
gHaUFsa6euur0PXmEZdRdVxqOWmCK96+nP/VI6ngJr0phfFcWTh8SDOwc+N8oAlEfV0kFF6OW6ih
yBmycPqy91x31OVpgxfrM7qYAYCj1bb7xoUfBScTG2t0S7c0vJp71AVKU3+OlM80DQGpF2zgGhSQ
pI3165+GOKegNzwMysK9mddP3VJdLUvODAcZxYmluVo0O2TW9YTjBGJwP4yVST73cTpIVI0bzj6/
ca7QyCZ2+9sM1ccfkRVusIh2EArslrlxjzyOL7gr2fod4vT0Hbs4NT3Xka59Q3stMq2u2bXoy1Oc
4VeIvJLoiQqa5y0E20dYYQz3LKdzcVwvOxQjtm1skBzAllttwWha12vXe6883kyBwnu3nTIIy7Kc
VzveNJOMY3Tqhu7IyCM0WYlNyj+ZQHz+0B1YIuMrWrZqHqm7+2Bc9rMGWwP25+vVBQxW6u7GzLA4
Y8v84AShPC8ht+JPfExDnnaDczowER5VYvTlVdoR0lYI1G1HWd4CIJ7SCI2tb/eOruvBNmaHlfIb
Ft3Bfsgg2j+0vBFBa1kz9NlXsj5TN6baPqb3AKx518Q1odaekv0Npb+jVIVkalYZRFcweFspzkpv
S7pf7pked4ESlyyrxnC/M/u57oCd46Xj8yp6lkEKXeTHfk/gsd+EvjCQi/Neuwts+urgOyEmSyuG
gYqmVp6m1HTKy0TdGJg6eCfcrycyTvh/VOF95TVltc8YykG+G1oUQ8shMfRXdLomHL0YQNSs/93Z
ajzQ9+vBDGxLuu0RV9xcC7/zX1rgRCkFafLh+0/42z2b3R46Wn0IrM+j5ky7xCmFIVDzru7FHQDD
Lxpwm+mdA/krsLbORVoW9zW0TpZ41wvsh0EQk7dmpkHl+6TRNjLsT4BAsEYzjJzzJyvBOta+Skb5
CnRI25wVPPwZhx439DwBx9HuHCdlHr+WT4DrmhhQ9z1oYPJ/+XsAn8nbdcuEF/uwQvxflmEhp2CP
6HaDSky9iN9gyS8HPvJllqx6+YGhXkEj4IlAkbljno0yxNT/rYwaWEWOZAvvrs3P+FplRA9jNXLM
fANtGNj6wMKLcScTgQ6AOOXWYn/R9h/CrxGYMxStJNQKEZBPxKU4SGeaxLWkiIB23Towp4GFm4Y8
IWtcNRpdmj2le6uG73ybsLL0ywQsyECtYNQtktbFBjGPyq1DLftyYDW5PaRRTi/Su6e2UMtg6URG
5ENlkcOSLa58RLLLS+YoNBIRycCYvgiXrhC3te3RK80DugViUelwYLPHGRpTjyiz2rDvg18JpCsO
6IBnc5CO+DUlX4MD4Rc+eHtAjXIbohaJea2+o/pcSRHxuqdYtOGG+sC90llgDbN2kNwBqXd41KX2
p3Z7wlp/xbozXc8pBrghBPTTZ9cLapxaq0eoPPeVy6MpdQCPBwQFbE0zPzSGF8VqLFQZeZbPabDA
9d0xmguZrzOTJIkQM3aSYe8VteUP92tTVtWPkYsDu5NTaNNGOhbkSAlIkh8L5OQc+YneBptM8Lyc
WG0Dkw48U6nVSWUSgM7Q4AlggrhruMBs4HcBz+x7gN5AAZofcYlwx0+/kbMFvXOSJVq7ppqPocEO
C+DhsnG6gz6tQKKIJ04/z0q/8yUczlw9qAhVtLnmx0PSXs/LOBpiqG3SLmqTOhadbCMfUuoRpKYz
4iDd5patpMG+loMrpAPlsf3kF8XyJUzlc+GmhwziQw9Fr7p7dhyC5G5Fxpvi5GnEhLMyG//9bmQA
G2Htbx+tDZId6U9+EzeLdFFJ9BnA14D+ErAQFhImXAS5f3ldilI/o6ttWlNUNd8xPQGWlpBsXYvt
hcOlO/9ITk8OvFf3JTlvFDOpGyT51OwUvYtLMmnTaj2W2ulfIFj6RMOAlM/fJ8DfB+iLGxRNcakv
AXhTXvolMb4m+ke9BVIHmxzCL1FqvhawDoMD+3X84QpRAjqUzMhVLbWyebEmucfRU0BI16w5D6Rh
jlwZlJswXy0JpoJ0lULBe88PGENctDD2LAS5mWJhhaQMdSG+6lRiW7ClJuzqW27sZ4UNNNfWZMZt
YuBSlY4hwqMP1uHMIv/q4jS5vIfMXdZTnqpEZTVkM4QDsY6aAY522xrNSsq4q0CrUNz2664PZ4/Y
wrSf4u1F2pWcEIGugnWLylrwp+GYdjMuqDcm43/sOMJJ6ucrvYVt2OGHSPwyrGoc79mMl/YqxFPN
O/MPZdyYdOCDJs4y5YqlFLK3YgFCNS7jfr0N1lJ0DPWa3L7TO7HyYvred/T2QReKeBy1B7/DH/SL
rdZl3n1yLS9IyqR604JEWLo9tCJun/CAGSR+rCDud3EnvjIWkKMfU7wUDjqkrUEab+NkUP2DfMf3
0TMOPgLXZPSmuo/76apIS2WicOsJcUqycyDh+sB6Rc9J1zN/Zq3JLYLm5XqlVzH/Cw+k2eXSvjKn
aZpv8i11lFqon92k1ZlqZzk6UNXEL9nQuV4kXGuFx8GWOouDNik87RIR8ptEblMUmSch4grO479y
TVCY1DUj4BNBnUODXU0tBVRjWd5jmqzSBw0wQO3VUrmmdEbra67r6dx0YVeRqcJRKv5aRi5sYAgB
mXo8BP2cxicRZF5EH1J0BTXQPiMx0kxV/JD1XAWSE10KBhy06/VmMA91yToryEwz9Qb6NQbayyNg
bnpWwnfjX3fuFhgn/+ZBOGxg5FhVZ1nch+y8IdQgpBuUIL+m/i035vyidhmT+QU34Kt+VZ78CSD5
3sQKI1hnAErIJEi12WOSjVe5bZWZFMu5nMBiwIuUm3BZRdNQQhJ7kgM6qC4FOudNKW4B/rkXOI6W
WABxWdmQa1mNfBmAJkVcPW2gNTeI6R8uLHVxFH3I0y88uU0V7/CmmOG6HgfAzRKdgt790IjzAoS9
+byf+hy8oEbTlc2C7HeN+VyAxgPGbD4jxl0e3AapPgVQEuemaVg0YtEjju0kHB1I/nuVN2eCyrXW
+A5wGxkJj4PwUm+0aU567P3/Mgs6s7renpEd5Qz92wJPvfho5qTca/MG1GwIatTt9t46mdOQDAw3
1cS5+qagnGbc07DXDQ/vnWsfQbwwJw+c2J1EC3+CFziXazGXpHUZTObDvX/Qq4lXSQtrHnx+egT3
hScCdtDkk3WPckFliEZA1QP5YAgtUr37jswi6PRFEQ0y7sR08216b1fOb4advCNZ/95FrTv3zbxD
pri4X3P7JUaQKlKSdKYnBPCS+/mtxfA9ysaTE+ElpCVDRtjHDhCmib0Ds9fMNfRIS/Pv6nUCP3HE
BCQT+RDsT9k68VfonJ21jBpHvfcV5cA+SZ/YaoT2eipKRDpes0cqQZ5Mwi6UYrVR+cTI3+pai2F8
G4014cQTqUbxsx0xdNw+SKoLtvcE6avq5XYfgD3N/H9YBAf1osfBfcloE0NFy3t4lyJTCVwHubna
gJbkipO37/f3LItsonTcS8XIJJykqQjAB08sy5u7jOVphZhn7Ej312d+1tfSQYnyGkYpOG4RvCds
XMaRft/ww9ZQ3J6FZTpBBiZnWMwmHzAlkKU2JoJRoDOvs0r/4dLjCDA4+lkbed49sdplCDiwnwJh
7tBkKmtOFIKV9qMqGKDrvcRS+40fsL/1MEBUvdefKsdCojrxmErBvRPjAnUnvDH3e38PEAbEM7Cz
FH0AByEhh4ZfBmQ6Hf6nk1gX3C71UP1WibYDvifOHPLzJY/SFq5yDQS0BB26e0/yVUC1rmm8LOFW
J+xpcbjZ38ZvElC6Pq2VAh4zJcnsSFk1UqNc20OWNG3u78qUYJC5cQWucEtZdkgCQmsICOPFQVRK
KFd3QqB5swe/nhhYsu0vYf+1RRVzfqx1++e7G7lr5F3GWGYeU2bug71kUBhva8Vfu4GzFDVXvwYo
J08dRt5cl/r4GGx1y2/nPNj47GCzot7FqzmrNqtVDovUtgUyeQIR33wYb4xT2FsjHYNofJETrxsr
7BWWAnTS6zQWAF11RHW6FYwTKL1+e4Ln13AM7p4MDLPHVF00gizRAzHmb7yPaUOGvajbmJ5q/JhW
SieYnfvzMSS+2OxrbX0VGw1ZtCL33IBdfRJfGhocjutg3fcIRGlfwQuz2B1BVDNrkYjfSjjchzZv
dBCE5CsMpFfhpNXZ8G8xAztqgTJmEw+FACBYk6FDPIaD/rZLXdqwQsjIdt8HHbmwdU6Bm1RK9rje
hbprTHzh11xcy0iYbdEgjG+B6jRfj/DEO7lt2pfEMSgCa/IZIcXb7diw0G/gqagYyKFn9q+a+bPt
vUgJEiphIXlMEDpbjOkd/A8dwIM4I7tjuC/vqPpmUv8+C8xY9Uare0S+NYWaG2TEKo7jMcB+A1HE
e7PRbQhOuUiLTuBviwQrysbtxlEkU1akv1v2HeOnMn70hH6sfWdr7Dcm3W9tz9Kr6/kUaR3ArfP4
JWsTWI7Z/1MGB6HpjN5YATCRb5xKNVlmB++WfBQoF6n8+8MHB411A5Y8c5mdRtackiH7c/xLED8n
zbaNdS9tU1XHztjaELhoApnEDLhc4U8SkumsXBKpOHNsau6aO2/efyppX0Aq66SKjByTyubMeyzx
CoPxj1jbzZU1K1zRvE0OuMTyJgSIaMyKecIzu9p6Vfn6nntvk/KCSuJzIvFLl56X660dFi/7CBto
ZUX7DQ62S8DQp2ao4wuqEZ7HVXCVhp+csR6tjqUIY+TcRx+nU+sTqqLAidv8XmtyWJb5Fm+LDLxy
KBrMe6zcgqca+mQ3AKeD/Z2YNmG1706HDVzKFUX668AxYsP/CTU6rN0ibsT5EYh+tg/dYYBhe84/
8LgdoqCWyYkea/cZNBrnGj8HLnlkxYjFBURKVWFGSNs0RdWkqWP5/ntzli8Wb9oKaJ6xc/hH5aDP
1SM+QRFT9yilIwP4lhaotnc9WbvGeosnUaa0t8e4WL2vr/fkWsAYjCOXiywV3CRwY3E8IE8L5CoB
tCQpoC6YXZSvIVWIDtb5/JLpWT2Vl/3oGji9XxtnBLPztwgA64kcrH4WeoBJgXGY1OAXH9WN6qcW
qfEa7lXBdC6ukl0WyVpVLho1hy5quqW988jw68y4JqhBQKNHKGhtByZiXtapvSw7pD3mPa+WkDY5
tmBsPf1HvVOYXZgxDzoDRk4XhFvBn3FlaUoOQc0SMYV1GldCAeN0MiHucOcwCNs1EDfx7YqnXydy
MVJkEMI9zNiiIAdMfWRmFAFqbmpH8TpQ+Ghssd4KF+ieYANlG2Ia465xd1SldwSYrukslOw69D20
vpsFxlYQdM+WP7MMRi/fl0lVYkd7A9yWAveR//1K9cVYzHqYDwkKTmO/tkLwPXEJWNUQOTbeVe7I
GolXROmqvohCvrmLRZgwW6ALe2db0D3hjak5B1t59YczB5DLr51JBJFIWjW0acUvUJe/bat6e5Fr
Aa3L1FxxQ/1DewicXrmyZXJFTL59SIq8zTpghoMfE2aZm3UcCr5wGdcqqHLnusazY38JWyUVFNlb
LLlrQ1t+xjUCNPSEBm4he7Cy11LEL9DYOXSRcTl1qFBIKMnV8xv3fklR2fZGYRRKHeKeDVIJAn46
dVgeqbdstTlQQbv1Bwwat0Aq/+gb9mHHPXF30PLwjwk/hZs6i2b67JNyhT4Q3ZOrMBMXjSXBQlKs
nCPSpG5cu92Oa9MvBTCb4/efEaEvShECBGfCjVpxUt+esHzlXUAruF4wpwC69sq9R+98rL5XyIGF
0PEGwNurYmyCR+c/G6e8ovYtSmk5WP8RL6Fsr7WT+k85TK6pCWnoZklfXsJwGuWhpd7yYofgBxQz
767mCWsEQQ5nTISX2RWLj0eRgr3LdBBDyYhPChu+796n11bdaU7/tEI2+mBkoCZ6LTwIq9+qtQrW
nnMvbNajDApazFPY+fh0V+9sfOb6R9K+V1Jct0VHl4wBBU5H2SNJjOBrefNfauBMnaQkB62wtqnQ
lRG8W5MVilhpy/EZLycf212St+rvXMwTEQpWi0qU5Vv6vVLso56V//4FyreoYBiAYQrvspYFaLMe
LN8yMmg1wFw7fjfjGq/fNsHk7PYAPivxpx/0Z9//Ej456oECTvOWra/BOuSxtZCSC3YMPcSacAM0
3QKo7ENHTL8El0v3sOQ3n/bNPt0cR8sJ3ibUZ/VfTcgEa3Sy8Jvp3i21JWQIXAjXbNN3WMWL2Efg
il/5Alhk4GIOLvJrW/3xW49eeB4qa/SJrw0LXT8RyXK8GbtTBgUa8Fq9xIjKOk1JHZEiTuymPtYf
X91aEhKLrmJmHL0ePSooF52TR5H950rsiyNua8C9r5z/dpm1fWnReohZ+mj37L0NDXGjv/Ps4/Co
ViEUGUGrowUIR0kDLKznpqgfvlmbRRdUNM9mkPdT6JRmdoZPwp8ovhVFXVn0x8xFfWDb2+jM+E3H
8r+PyUG4P/tTiD8frpyieu3VTBcUXNnmFjr9qexx9XBIHsY4FGjddolhZy4Hgjoo0Tw0GpwdZbKU
WR8tjUb9s6+H3VwaZo45B4hGRozvzkqaMlXmJ2edbLssS3Vxsf5h7fVSY8Nxb+pIGtg0PcG7EOJ9
JEB4SpnwYI/8xr9SseE0Ehc6E7bzz7DDSwOC5meRh49spOlhjMClh6uTZdv81RMItKduhGVWgxlx
zANjgwvpPsnnsFzarB1eJGJNeq57qX8hmenB2gd1QPHJQucly7UfptHTSQ0gw5qpiEPfLuWgxgFZ
DIQqPb4GYIYwm2Um2QNJlzvo93GXzMaePcoZ1OngkGm+FKgvjuqjfjpxPQwHghXXTl60NunrQQUu
4cqnXPkIQ7QCNHLk2UxPL4oJBUXUHad/kIeC06PM9FFFhYPn6sPr/Pab/vT5BIrZlsIIWH63umvt
GuokO1JGSPkgW6mQFtqIvMyNDGlbnxfDyMa6FrzMHgMKIZR6mlLBRrR8B0elqR6BvzhWLUqJ2j/V
zztqg7DlVnnOOSdD3GDvm7NbP+Od0eIgh4uOF/FANXCmCFT4ZAnwNYQdzAb3ctASCfIQt4gl+MBv
rXtoINqtCjzdBgXsbScuQPokB8gs/mb44Lg8FxT5fx2yVTAigh3j69Hg/OfVnveVE25uWdkQx3yq
gUpJUhqfSF2oU0D53mIH52P6vf6Jbie9Oa3v58YXMKIlXZL9O0wDy07w2S+ddvskc+UK2slcuCPm
z8BFshUWb2v1BRNKpXJ5wO/Ybz+F42Yv5kHNs/dh90kqeoDX/h4bOgZQTc5utp1pfS5VPj5vb0Rr
yUY+LRWhn6nYXAlgN4YnfLpw94gmRPIfAqg8H7gjcpQdUWAfit7W3DV0FrH/tNI3FOPfAvVNsSud
ZpH3yif9y6t+6jyOX2YG8KDrDQN67VEvyWK2CNuezDe+D0MCxgpdBFdD5WUk4xXBQU5V8jm7TVHu
dzpGFKzDJrCcikrqIm9Rsi9qFL1TgzfLOeHSTGZVMW6TXpXpro+TVJa9oNnGKCHM9gldiKWFjRIA
zTwJZoqn3DzE0ixh9Eizbu3xNeXXjx0feREma7bXetsm3y4PUHW5FbpuBoxGJlMjUwgx2vWRhNz8
ozWzgkyRp6ehs19IJAK7CKzZFDZURkW+1eoQg1jz698PdpeF192oet4+Qk+neQNGd1jniRJhrC1v
hvYwnkHUzdOh1/dPdeoxyeeAiZn1PTFsohfWFKSN+sVjqhnjyZibEoNulgbsvr1er9aUfUZo4iHA
QMYkdlJpBvnYmzW99/1vTxHlLRud1G7O52ZFKK2rvHybon29nPQDYf7PNf4XjC0ZTsN1RgenOiTL
NVYpq7opTWGEky2ReIpD3Mbh/YuuENErML12juNYOp0MnjgjNe7HXvFm7J79rlEg53QEqbtUYbTf
RzULbTBklRaV0G7Dna5YQrRkR0rj6YAY13I39uG8xQQzW8MSz/Jcx/NV8V79zHsknOEcVpkwnhHM
A/zt066US7HioWxgU21h8ZTkCmHRkunErpZ3ZDS+2JCUfZqoL3VnKEy09bsqLRWj0IZJAJeaddM3
DXBFkBy8W+VtBd+mj7RiwDXd48+a3ElRq5IehqEW3Z0IYdztyph/ivCcSHMdHkuP9TQ/VS2DY/EL
8ZpMFwK6weODpucMjnzQbBwW7R74f1B5EGb37jsK4bX+UHKDa1Eo3hWOPg8dYJb+cFjLaNpenqAF
p+nUCIZxwFkHKXO4dIQ0/7vAsIsz+54o4ObGR3y5xmbvs2rHhALymzzX1REKr1EJUTrxBLavkuDt
M2lwdMDTjXQCL0+UvsxybB0GFJEltJ90tjMyD2LpPfcLKHjcZSkv3ChbkYYDWyDoZ69PYldc9wnl
VsNEal06SPwCBknND6cd6FmGeRbuV7C7BXCqviLiMkTPvC1CogJdgS2wNvxjCI7O5BKfuEoQYmuY
Zqwy5wMnp7XqVaf42+rffMLdQ1gXvHlqcWeasOXLg0nRrVwe4FrMZdvO2uH+rCwwFjFC7zIV/VFZ
jnJAeL1yy+G8yw9pcY40dSpC7QBpXz+yKEoCKSEtvz7+aBPGkB6kjTKEKdX41QwDj/+RQxOuFM3G
Qe0p+GuMKmFrIS9ot7DAnGU5rPsCOMnDQtAXQEIqKpFCXamwWxzYjj8DxAU1mZqStUKjvex6lWCS
PvZUgWyk8IlWYbCNqWqfFEWfSbvTRzgYj/Niwkd2wmyi9XS4slt4/QNpXUL22ZiIcCT0XEivDhSn
/0Wen2tWKMEg+LEA6D7vcwq9CBZhJ/qN5tJ8pAx1XposWuW+143sqELT5MC+GdLGiI1UuES4LxS6
OynCHN5U2jFy0+womhZAmbonuJRkBzATaboovz/qWjPcKEZRDzsRfCoJ8yeWbqLON4sQrDR/HFDZ
EgrCg5wuZxE0bVdo7Q3VIV0gLYLfsehSI7DuBvh+tY6RxucEOYvDubiuz+VIcg6g8HStbWIHXc+m
i1ZtsbPb5NXximP/8aDFje/AswnqwmyrE4kVdxENUi3Yd1XquWvYoz7lxec3bSsPUN17rQdcZ8ap
81acd55Jfxep9+ufKb3dUr/0WkgnNttH0/9xjr5VW91cdUTkBaWKixczN+P0OAxuD9pEFeGqfrnn
Rlw2OReStcc5C8O0LVY4yQ5SEia3IceO68uI1ETV4wQprfKLm9mGyattuiCysId83p9Hki86NxOd
gHltMg81mqKN7j6FMcno/mOQDbFBQf+MZ//a2ps5IWAHKP8DsBU6pFrX8hOL4GN6+NBsGLXoMIWu
K+gtUfaXJIStmkGNK0Vj8CES8bT3J95QPpydqJDaM+6zmbzo3N8TosYjld1Tt2TH1NDUHgmk4RhK
p/PK24xqZBG06rRz/oKx3h3d4BrTyjpxQWvNOnCel57rlKVII57yWjR+nlnLcT7hfBPrv++lgFc9
qQVNXxQEhEJYBIUWumLERqFQRFE0c2x94DKp4CLYf+y5LDJaZBZFtTd3zA9okeelQ+wiU4x36KGx
tsietL81Fbdu7n05kAJFqEoAkUYopWTIt9wPbahRhBGpUhzyB94vbbMPWA4/axQ0e5DYGU6ukPq/
cx77NmyD4pQugViGNGa8SnNjBakTgiXsbVuXC5VL+IZ9H75rRiXDpPdY96cgoS1vi+CGlQgMCB62
QK9NhdWfvIqdgepM4sCEEeWutka4LPSb+Uzq8x1yskTGu0F/IEz/+7Ihw2r2FQksBAvypZC8IIOi
DOUkGU5uGPjfzqpnXSUTZjK1FczM0hxOn14AAZ7elKtfME6ATkCzlPy9oKBSRMs/TUt+E5zVmzax
RsCNSPCQ8DFgLsWhvbC9lK3FXo4NxHVnb3Y5UNxYmwH+0PJ4S9MVn6c/sqftly+YkgyS9HGx17QK
MKNimIGoqJbpvfu5b/ei41Q+sOKW+S1TrirqzHQfiHLm0d7xWh7J6wwbThomGz1tHiy2SCjm8xIi
VK0n/Xu5n5D1t4MrnXMy1bH6F73WAsfd9wD6sANogo4mM6NcDpuKQ7W6BGS001SLbGDUUdfYXZAS
QHnPkuXgk1k4ROag9SLfIeeJKXTmHLdDoYmYKa0FE15G+tXgDgz3y0bfpxLjCpBn72DSR0bDJ8oc
hTGZrJX7U3xNTwUbNeEqxEgsBureJvV+/4cQb1U8r4ohiOPkQSJLXumRl3KEaF07QA9TIF5rF74+
GDPRJuGe2EOBvQdrvlQdSE5QUgScU/25k8FO5LZQ9b+AlGhXhhu6hWjqfp1nv3z7yxtLpHqYwQvc
+lJuVolpcQujCd9ZLJxLIWkqBJ7kEZKZ8BkKth6ILmVx1BHon5tL+IvhLEV+n6xutlcujbC/vqOG
fjQTs7d9v2t0tQaeY4zCEbM4873UmW/D5PRRgcfNvsbEvpwwnhSIN/Bs+HkGfDUv5WnhcKwMbHT4
410a8UvF6wXqQ/Y3Ca25au8JPeY9m3BLXsO9yxoS0sl44dmQv5mf7KMeNwimbO1bUAfrJm9Agr4t
sJLt3FiRK9cxKJZrYtJj+7XCblRW2FzEotx+hCpwpISXJmHGz+dkkfWS2lbbsgP0IdpKjwl24LYw
khlaSUZ3jQ6hzCrGJfvRQ9BGUWmDMuefU959LMacPNpn4II9GRjhYDwP9IabY7s7dsE5cCnjGrjQ
UAKgUdkFo8lnYTIesuiPF9TG8Lg4Ewr4iC+E3gHyUfQbIpQwQe7rC7YuHrX0bfZUNCYVXBl4Mmsp
R6Cg0JcJ08LQ1aoaxP6uSesfwpk39dT5yI1jtMi9wZ6O/zrk5SirB/lfh1hQ98ZDoOTgj/3xxuYa
0oHMgjF8HsFRBShHXUHpZbBaWprAsRA1SvL3Zd7uf+3LQCnt3J3qpgEd8iGY+fnCNWQK5mxsQ8Gh
skovojnB8SENqkmBDnHtzsinjU8cmxMmykUEY2hzUwvnNBmTiWurz1+95EIRmMpYgpnXJWYUZAx9
fobIyxov0PUSrWCnnZl59GEOpKpI5s0lvTASg2G5tFn0pg+N+0sllwFNtDKDnrXk4M2sjzkCtTeF
B3WhpkwXQmPRu7btxDEJqAMYvflP4JnDRz7uKcFHVpNXjwA0QTF6bEhrD9MleU/EfjZrLXDpuxQp
tn1JFGHs15vX+Ew33mndt8LgsT8zh8J/Fd4bnA/YL5QvewphxQtYds8wQY2k7md9wVIy5S4SVb5C
YBNws6qmcaaa8nKs/pF1ilYHcwSF3tf/vpTPQL5cXPsSXZD1JkSrFSk4BSN+QrqkDIcvsXh1NOMF
+hjdHrRdoNJGDNyRIGV3WupH69ahW0RGovO68qCvZ1B40uDoyxd2DFuSblU2H5QCEEuaIU6tHNUt
KyilbPQQTUyIKb46m4MWXWspI2BIzK72dHO0hqDe9eUoCqRKepH+2rTxoGi9nvOA/WZuk77t3G5h
gx+jr1KGRcoPJCi9K2AtAdZZTN5FcDVhjb6yH/i+n0VOATfy3rvixwhJARzVnM8OgOdpLMKvys29
7ZyS3f9qS3RtINfNItBJ3vYCg+/MulAZij9mSILWpf0+WL7ebSRPQspFwukTt9YtYpEAVeUPpDsS
0g0PWGN8biWAtkxWiz8+AtmepRm3b49rMWYDSy9TGMy8mKr/22A+gKwZ+B94SgzglBC3oN2UcXID
HizHrezlP06HhSwQ2gCT9aM9elEJU1/8AGSMyJWCQpvBiYDfwRrCWtOvuI6RKp47Y+aBrvqUI/Rf
hA1ShFpgW7Fm6OcPUVFRGjYVnzguB1GToBaLpg5HcS4vvPMRrA6uQ5ySwLLvmwxfMvL63/S01P/D
iq/dU6BksFqZPih8fe8IDO4h4Puvl1X8lcH1RIcUopdgFj8QoMLfZ/0e9CY2Np04A0MePbo1cR+/
Pk66nxFyC7K1s8EBpZoB+RjmcfLAK/d3d8SC/YnPCMO1dm2nc/ddDYh06Hz3EZHr2XYhDbxJP3Wd
bp8SIkNN3Q9fpVrAeGVvWu1f+dyCwQekuTGKSJvK/EwgwjxH/rYNUznU9UdS0zODBMlZPCJjeVYx
vBUqmC7txnTJXV9FkVOmsLCeJX5h7Ujxlx++HU68qZiYdX2akfhtaIRNi0I7jEExrlQ0QZrfJCwh
8Er+j2L/RkYDmrL4FodZ8p77UbEfIr5Iw6gw886yFNYlBDyEAXV81+PXjs5siI9/s2Jzd/HShT8s
FRiqsPSz+3oJgRLBRkqyQaNr+RnnzFoPaHZUsEWaHUx6FgS/VQARXATiIdvt2IUsV50nc/Mqj8sf
RCJzyg0GVkqOGJCkse8A4xytAJxtsHKKG1ayYcjw4OX2Pt+p66cioGTcwurfZczkbVx2hJh0cWZ5
77E+gP2VrF8tUPXIlMd/nwO4kDAmstrySVazC1CI9qHqnp0j3qEyVBfcV3ZMYK0M3evHg2QEQo/P
8v5YKxi+Ejq71Y7D12mK1I9KhaCMVcbARCr5fZi55FQg7Iqmb3vkZMSilZLHZ8iNsrt+PcGX1sVI
kAHyAyOiD1tsC71jSbXbRZNKpp4WB4qOgQ1kymIi3Hk9wbMlBMF1+Am6TbFcoOWtSf986JREKDcy
IqJKViQd4pPpxR78MNmdIsZR4FOeIOFmhQ53N2rXqx4VxNrzg/2xdDJSMHTfMS2+EOOWbaliDo8R
QTt149RB283WIbBd2j2piygWVVuglr0CP7fjjfbZ9dmSJWnasG/TeJCM1L5lgl+mFcKTu7M2d0y+
m1BjFmSp2zyI1mRmPL4Gd3vx7TMb5pIB1CeKwcuypB6szczG3yIySoerUqy3DDy+5fwpQoSJGZ+S
XqJlZe1+zMYwckfwjOmZy6rjrAD0nYA1RM8BdorMkJecV2LA7wx/i5+/woU1omcZPleeNPHKJnin
J5CWeBX/LD6khQsUp+/b9OEDlujA8yaJ1WqyEPItngW+INwcUrNjV5Wfsn0zlgZMWY0K1V+J1qdA
JC67gejdNQKLt63+UfH98frummusRV5m4qx8cDUrCyYcknlxWJWYcAh8vDcgN1q5QH0V4eHs3JDL
saBKGVbrCdlWjySpJfq439CL0Rgu+ZoPve3Y6td75huY5gfyJn2Wehl6fn1h9MUtV96XADBVL5eJ
OxFTEogqN98Y1vF9I5QqMI0HE5HS6FRr3Ax9dl9AKyy89YRYvNOuLzPSoPMd/DQQ/ZYTgKKTAP+j
kmPjVXCJBdDYWiAEhgv8dBM1gEspMcxfYQ0MfY/p5Q5la4NR9wPM+7cxp9MqBKeTZua5RAup4cAY
zdLNDiBZaLOJt8qeNEwFdGeBXscJn/+wvFZBiNG0PulPJtsHE4GwZwxyU7+O6kGzgmpGxhwJ0CwC
lYVb6kYLIkLnJ47RnvGkIgzjrigrQgKIIpGNd+izlnkGFm1aAxOPpj4NJ+VKKmuqHWvtBXr88SIq
auHDzzVFDQQy7L0kJunHQh/J218iB5ZcO1JSzN7fg21y0eibTg1MLJKt5LBRh/coaW4C/9YQMAIb
OwvhnyGek1CeZqbkKFkhYtkJ24EvWFCfF/j8NbRSXDt+Gd5O/fadpnb9lEUTRuvMVXhzWZwX7SZ7
JsNqgCDGB2V6iAcOC3uBgc7wtqf9YQqPodElH3ccja7wtqqulGCrbpFtg3zWsHfcVbP26A/m40/K
xtBZrsC5aRRNmxNG1J9c/BjPgVAtX505pfunbUPx4PfUHN4K3C37LBRLSxNOssnufG5oimyY1Ehm
21YKo/HZdeerPpBUjwioUvFrPcF4GR48do4V1buKOvC0H34jz27Qb1dyNNoaSQxBnEy3W88CmPBT
kS/wn2TjvctIxRhmvKRrZly8c70GEN1yypoF/KIBnW2muNuyCfF5kSsrPO9+PkCnRM9sKqJxL1mD
ZpuWJz/SZ6AVmBA6lrpSRw3vuLE4Gp31DtoNamYJ2e9x5gHZtYWAxn1516TLJ+pP0zH6DwfyvjKN
Plnuw8Cseam/KpKuAp/SECEnMl6O1htNltEkTQ0bOsJID+Oq19Vf+QydnKNawoi2K0yW5Rw5ggoA
ZXyyc5JOw2M/6xGm/NSOp4vCeThgXM/P0uDYjrAADvxMSxI/DYO3nwVvgnSSa/Tu/EgSMcs/t0oL
PMGTmbWiqAH4SndboTVPO94fHtoxK5dXGs4YFMvvstGMkkxb7gzxwBE85f13HzDkveyTUwQFlmYp
a+3KSAedmCD0CB84As+b/m3x5ltVPOlKdzN/Y/99737xnC1eGxOm2obwhRvRruMz4TipPsKTmbz/
qaYMghrYNPQciApQhqNYDcER6mYhxWtFXyc0MUfIwyeca/bWv0+Q7NY5s702d3n5xVvHE4Sodgf5
vRmUUYSTaTgRvDre+6Hok8AVSXW7pfWMDakC+W/2C7LyS2viyV9FonDBFzt44Xc12xoo4chakwhH
i8cBuJbhrrjs8Hucz1jna/W3FCUnAx8AntOkSTbaKswgJJcaqEsCBcsLow3sNpGgav9Rei2KgLbC
bWMEIT7gA04EOnTLdiFmfAfdmRFtIizlztKbOwXuDRU3r5a/DLfsIEkO2YNbZV1oizSn9Lz1JVVN
lCjCsJfE7dyzDjRYBl/J+Vx128MiweFi4WAieoJnBgeadsBIdr6fCJizeElRuSbWQp3PU/eFJHr8
/xzl/lsydWcgcR43pFJCVY57HFkiqzn0r+w8qzOsPuFXMiLZCrk+975HjuaipSJ5401oN/W9qtLq
xkDsj67qi4cxGSPfT8odKYVNclvuWWlWvDRHPKIBkxvs2m7PF1u+XL+njpsuWlgC0KZ+yK6iGFl8
S3MrhK38hHpEXZhnndfnnpfcoExO7r+fnQnoPLcRoT2lj8qcEYFWC6rjOFGc0+6KZ6c/484oB+U9
V5UX6QuiwVGbKdiMZw5mq77FlBfA3rR2GGiAuqsEi425N2CM8CWwmyEGRS8k0oKpeCan88x7k9k2
kQcrf8IWTvnNc7+boc1Fo07EYyleuTPi4EEUQVIPnUpcBtIQT09ncGCxkwEJnsJX860inMJsTcqd
Nd33VH+/VMLHRZY79RJHFPcUl6HTCGUAEov9VyMtv9Cgw9VQREoeu1RNbKL1AGKOnAMk+9thlmn2
mg/6P1Zgi2D2A0THFbs9/wq0lISUGTGnJ4XHoXx1sLmy8qg/I1uNpnV0Cl2aBv/hzeENtZeIClcU
m2A1yQZIuchMScdTUVgr0DvE2A6uwo/CpvJOx2sfjDqAfzEFYIXg03mcmXulV0l3OUO738HuEll+
LXKiv0B495YMCC0vri9fjQgmQ91OUXU79xhoMTDMY59cj0nWTUXr2pa8Ry37T2kT+pm2V3ZUS3Cw
RQT4y7MMbwyxXUWfsZDWdoYWE9fhj1bgylCqtJBwbENPBFIFhnx6lEe+cepCfxtGxR0sMizbtWRu
RB3vbmuQxFhasjS4g3rXQiux8hUGcPbsAJqMmVb9zPxWklg5Fzs5duXb1TPlEjetYmiomE0zZ2+v
7639InelScLLUKCJX5lY7wM/H0AbiKU0kFJ2TLmTqN16hsuDqaMr/PjPmM+CWsMNqlJaaQY8fMlw
2oTn72UyWCKbfoWeBWjDR3DuMHF1ZF6fb51jd4Xt6LZLf2juAIp9M2DfqSjt9syuIjM9OSMWd/Q6
vn0wDif/+xOQU8CrIeCmWzOsBvLp7PtC5G5zoF62UPJEFN7LQYiE0Sg+AXMgnAj+/BexrSIkogjW
LVn51METzIy95lNHBmu3tTMZKSt2c+CIaqgQ2liekzAKDbDn0mWvxzwhgPmO4t+eMB1WQYSJF2Qb
cmPH9kgg8TSP0tXrT3GIrICQY/iHRvL19M2ftH9sbfkQFKJQ56xLNteKdlPmeBXHnh3sQgKHESVC
sqMObbQSCFmrhvwxsUbK7OGthio1DNpI7isLQpiJYctQ72WuEh7pEJXZCPA9wReTNcl4O/fjevZi
54RKsVcs1I/KbmICT3HYq0mOfmz0Iz6hAvAwVjmPcIoG2MKg8VZNOGGH0dtgGEqF3mVoKn9c7HGD
KgGfn+dh/UWOCQdGojHrpoPfyjrLfPtLiNDoCxCxen5cOEHNgN0KrBcr+ZV7v9esNMFEQGHwi9jz
R0WFTGBKkuvAYdPJBN1UPIdKA5IRBaBO4ycmETARau1q6KxAuZ4O/rYACW2iymDYO7DTX8oUXYni
RuwP+MaOoMXZ+iXvUaYB0KFM9of2jaeLn7AawZU58SQ1+QWwWnU8/FYbyhCoV3VPx1qvlZK8/w4x
Mjk/Z9HXmEx4mYgHppyLwc5Lw//AmuPg7zxHJRg973JOXX8t7siJIbD9GTBAjjKKzVM/pyGk7A0t
bz1w56OhxHkM7FkX6p6rK+v1lmjHAhi5rqg2zVa/iXtzXw0Yijq7bj0vra7PmVvEE3dtWTY09QKF
fR6ChhIGa9VpshJacKeMuvusbZ/c5tRREj6itnt/3mPX5Xee/f8tLZrGhfMEfAj3Dx03YBrr9S4K
Wahsi4nPAKlr/2FZwNGNd4bSJFKKtV7SYCPZCIfKi9SkCaVDa7gl7ezafT1/YFt5Ju3kRSSw5FVC
icdh5jikWGcvBaBk3G2QhjDTyBnlpAuYpfh616gTNM5Oj6q5mPNIzmxzFkENdwkd+x5/Jf3rJ9mx
4WD1kfD5BVcpm1+Uns96fqKGqicLRx7hkgzqV1qnp8cFVYllQ5XdOa8Wrvn2qzMi349zVVUxF7+t
s8kZfRK5ZLNKHCJnZGTFh1K1NrBIs5NOuQGm1mE5Jd5QoA0ruKeRgpyOva35JuvoRYoDtYZIMXNJ
ztVy04HzYR4yhyHCjjTJruSpBIhPfZLMoylBa7rZYymtwnYxFOesY2FFHIgFKtc6LJfcr94vdhzT
qTRU8f7HOnjqBnU1sswg1Kc3XmhdvmSLH5lozwbzIE3nFkWCKPJX0JEGjIW6KpoCfcsxiFmpiwqN
gm1ZlLr+lFNicR/xiFX2o5Sju45Wcyeo0VAEl/G7vxjNkf+WN28hOUaKJ2Qw3XTSuTdi3wrRJBiv
nbgI1Z4EX7zE91ipJCoDhtF8Q5w650VlCd/nWzS8hXJRJsf2J36RjvEtGePzyd6hU+PYkDv7wsHn
NDz2Y4cnPWWaoKtnRVLxfc0oxxdNWJ9fz1gHbJfviuGsPkNgdc2yLMYHvr6edRBn1dg1fFtIanVX
e+MaMCJrgk1iu+s/f5iZnqse8sxw3KWt2qwhnpEVj43kB/yQ2Opf0Zaxuz4X9s8Kutnwzy41vvr1
ApM/WXvt/ZX3Qr/fRRHL+Da6tlXWOVydoItAyxtH3brvRbNx9YQhx4PHs2G1fXSJiEobgN9vMYBi
6nETXnbTswblP/Z7gyw5L0b4WuNGmLtSogJhExw3bMmM1IBGNnb8SSMs59fT/ITzKVbTLWTCQ0wE
qU87wraaXRkzIXEAHv3+g++zvv5DRGb4Cikg0/41NKmOQQl5C32suoy85l+6LKaLjSDBKO+2wLx9
gf7UNK7nWj9d+KD529gxlK3Uc1BTdLjiywW37LA0pV1jzWwBgk5stLbR1JtF68NRJ6yuaZcNd+Zo
OCOz6D0bo/M7Z2RjWoTYX8KjT0mSoYyu9dVMkbyMSdDKL/V3DCrcTsejYsD+S9o/zjmngNXg/Hgw
as+DBQYPkXSHLc8yG3M7DIdflRW9UVrD5dyUhY6Q4GH4ut43mZUP+ewYgEzfp5dSqiQS/BUaGP1+
UUfVvrsrzYhbIay966yPYSr563PJVIeIs2oHJZdsXe+qk5wDSZ0/oVDPwXdWYN0SLFpIzzh1yzuy
OgNVW3LpXLCzVuOoXZJLPsEmlRuAPO4eap72bkE5vlh0u78fscM/ayLLZk2RcjlNhS76Kf0TOGK1
ZByLSxXEK6E1sEPTGYiVW53Mguegz5KcbNE97JrSlLv9KnKzm0Il97uOOmOT2EcaXgXvCfpV0Njf
OlOZgQ6qPv46bcGXetot6Zuwp5GN2P6IGhukPMKdtlq0/k0iX9kCvFuO3k7qWfX9UZKXPTPg3NRk
VABc09amD3zRyElCfzpGlqr56xSucehcJKetZkFDfJUQT4ONGAKNTDPPvcPcIju4YOKmjkpW720O
rUTq+UwEGhfvScN7jo63Ytw8lNm3TJcraEchxV/NHC3AbNq3SyabHbWco7SDnLtWkdj2bqxA1l12
2jMXOuQq86Va1QYEWXaWF6ClQLPlaAyXHhpn2/RpNSFlFcc9Kt9ZaeRslXXoitm5aG3IWCJxT6TN
J/wdPo9i0lEdq/ODdlf9fkc6ZU/3qDRF4YVDDadMsdxZ4OJ8KCtbZmigKwz4DjQz5bBSqReO5+sa
NCg0gTDU1LG71kwuIpVG8YdjFCURqfuJUWYU8ECd/qG3+ZazB0P1FFbAkeD167xwn1bUvYVnPeRv
3qbSFvMTr3v9wWh26/Nsd9g9exBz3/sCEgsshds8iYzSqDyJ45VbWtOn6LKkuRjd+oBRS5RwFmBU
H6n1S+6vjIE7RDg16oed+UkM4JO9tOqUkcWx/d9SBxSaGY07RYfH2ac1HcWir6OgQ0Fa7q9YTnxf
WAi1m7edO2BenKKk/iCFFmot9lmTfzyIF0aY15Wudkwau9GKbBx/sqH6eMD1v30i2Gy2pZCks0Yl
wKsHpFK8NcTg0ld9fN5BAAbz5G+cr2zKOptcz/xeMsokOQEiYG2H8PraOJOKUZbY4dceAqhywfKQ
pLBU0imxPc/XVFBzVYNjNAf5PB4NtNelAmRk4qu7+3Lc5eeoQl4lytYNjTVJrCokGKmft/arJNPV
QqtlEXyM4/yL0x8FolaDiRfKQGkX/wXyP5zPxaur7HPQ2Cgs2YqBZF7XgQlNeSG0vaTFJ18SI3Tj
WMVH1aZm+Sr6ErltrCAPKdAoqTq+CjCt4gRnyWsrZt/WtbZx6hj/bWQMggaIDd4YBEE1R1/0TJJn
KAXaqIEDYTOAVspJQhWchxRNunDNEgsZXGo9tbk7I/7giLIEeaEf6UXzry0AQK5ksb3VxF8P1Wg7
qvteQVz8zgcm+ZK51RNQ6ysLHypGlm+6jzKm3IIpTSnpxYMrUI/93Eq0MxLDKp7O+jJuU8H9wpGH
guYUwWLBBPIwYdY5mBczCwygsUUrmGZwEzSbQLrfEci9ahT3/PvnN/LqOp0OIih4TXe3PtFuHrWF
gfx3A/1gweV6VcfnWLeXwZZEAWrMcNFwyNE8DZPHNl7eZlXURfkdKde/4haI4S+A3cn6bVgWsC+4
PeBuBZcMpRh9CgK+D08dVfuFGIS8zD9uPVnboq76l06aV+lQnI7TD1lu6i/sfwgw6OgPH1id6vUc
gCFWicDtKeP0M3tOHYVLkLS0HXTsjPh+l+40d1Lrztv3PXTV4e76MIa4Fnh61PK0GfSsGr6IW1Br
otXthv0tjXSWhNvZ4Zc66leMY95P5nUDbEJq8RlHOa3X/7BZrOphjMnQ+Rh5DsrQ0okAkV6f+wq1
Q56EF8tnmgiSFwCWt/hyuFPuufHFiN1+osW2MoSGX7tdSno28MIML9aoSLgSk6Z37GH1Q40kT/qU
fFiJtZN3ZpudUFtYk0uO4o9upg/m+BdR8fqSCjK0Yo6yis6ibKxRU8RSkRxYRwxMaL6v0sva4gkz
q1quUvNSJIZ9cepKAYPkAIm4m4iWcaPuTBAr7OvA5ZrudP+0E1h/kcxdvSlxRtUdWbwkXj0RXRdD
O66kRge6j2T4zJXwSiB1w6207a48REOOqODNCE34+ritAuzpGJD3saYNvVplzXmxrUrb7a/Wz3Y8
5yjdf6GJP7GshcVZIzaepc0F1AntCX150dG5ZUub1qtT2R3VSSRFaHzA7py8i2DZtzSzy7Bz3FFr
MukGjwDDwiUL51l8Meu0QINN6vg2WUE+1e4miKOzGlOiM/7reF6j984S5kr7sQuKdX4Lf0c3fMBh
hlUXIs5DwAHE+w6r3JD3mA4HdMquxo+8N1iVpa9U2QfkjD8X2wUnJ+zyzr8p7exlwYHGPYs01m2s
PkJG94YosftDWx1zLwBDlddAvLr6AJovjtmlOA5KfdWvfpG9cv7cv5MqvlFxQMv2pHlOqVdofFV2
abbBf2yWvGPsbEC718+pejkFpouAf7giwJMwJTftKTCjy+ZEhLnjPLB9uIi3PwTBGKGrM/PsjewN
oz0Ltf2RDN26akx42rJNZjSma8MBncT1Mb707K/3tT1RjNobxeWAsye6235+b7RLV20YAB1dTmMc
Pm4TASNCMhw1r40gZVjAgIc4Vp2IkDPh/hklvB5pS5uz93RyG/6f0+c2ykV6cHclfwKkQ05DoplS
iDpAPgIMLQxnWDH0LUyRYDUY6IGEDiAyTmvEoCHmtj42DoOwHnWCMWFC+oQlD3rHGZcoKNhz7dgA
pd7xat6NVDYI3epdGNtGHayPHjjOU9O7Mz5NiNQB0zLE+LjHKG/UrconAwQlinhakZQ6/Y8JAYE9
EJeoEb/Peie+cBbgIdgXNxm6pTF9H5FuxX9dybo6W10Fa5RJf+YzwoD5ySoYW4nx8HgAwS9MJSiU
RUtzgJ2ZP6xoe1A8TKEej3GDm+hlFa1BBkqEEXoQbxns6AHgAfsW/2/D9oJG0z3r/3fgNU6HMcQN
3D0u5gDd8BJ7kfwj+wX2J/OoA+cFHSPxxnvoPieuD3N3Im5fZackZ06yG+U5CnvF/jisZyWeR3ZE
VEFFOjJ64whuMWkNmJvWLwguJabq3cXJ/KTcFOaOi+eMBVaNc6ToeDQCpGQK1A2IiNRbph5DejWz
P7ptsDjE46BJozj+DNBAKr7HV46Z2YK+1W2lD9l3x2L0YmCxQBl38bjvvDKm5216dtxFFu7aAl7s
5fJ/jjTcP+kNw1zSYlnik0QGWXuzzreUZ76ipEMMb8e1JsQrrDsIOSVsf+4DRr6d5gt9zMPuZjia
kpoVSUOL+Q7WOTEHRcQqqDhaDqYksUMCPwBM0M/eFnQZpfvTav7tFubgwW/R0Bo/QOCGaMY1r08m
d6UL9jF/Do4uDkWu0Fsf7LpiYbmQOpKcHIXxXrSBtaV3VoC6YBh8zuyXW5Wv/KbFZGamLgLO6aIe
VSbV0V/1no7KlrHC+3ezRNalfzSpozY8GBzua5O/6BbSx4wxqRShfTcZJhDlN+6IuCDaXUyDnYTB
2MagLycd4fZBZf8F5r31ZEiXYWbXJosgDK9tY3Uz3r852f061O4x7r+dc3Q3AhnYr/+e1AweQSpj
OGoJfR0taSbznXJsvg/7fl0XXiHiPcC4gjfhExyNnzoahIhcoPE6MO8PuqnZTyMjC3NiTo0UefvO
d9hztnOXhWNYXtAFc241I5wzrqoqUmEY6ULagm6P9bnvGwG255bgbN/AUf357SywQU1sN1uiNXLQ
QvNUqvKcwDsKN80sm6ILMcB6/af++pprrQjLD2MNnlyBBzNqu71wpG2/vclmyTXDBaXrKUdHV+cp
Yzt2MrK234uibo+qzbLKFuihZuK2/CUTYGdXmUA+uw97bZIKgSq0MJexzmzo5R9SCDm6+/ndReEh
6CncTCLLHkqrYzYBvDGMn1XpRUUThF0NJfuo+lsU9A/Wmh9IX6rUFDXCQYx3Gs2E2AlpY3IpI9kH
p4DE0KuWqyMHhJS5yPJWDf9azCv4d9PxbCbiqd7laHosDx9IE/FiTOKagOK15s3Uv1JrqIWUGDvD
Ra0V1LeR0yYL/LLkrqkyUPSVnCGKLSGyY5vl7IzGe2lJBEy1MUfQ5KxkRC+mMoutJGZTnCYiFZiO
xBDQIvutIgMXX41YZPlBeYr9bmvS38p8tEo06OrpiJnr0xOc3LSF8VOOiUk2w/wURWilw8OPjrhT
cW39t0ypCvEc7Ka1j/WzeKp91ECble0Z4Jjt2kB4u1Gv8g7glmDjGzfN1FrzPRAp77lAlqvZ8vTq
et7f1J45ITAaywqNwuOxvNvebmgf9H7Kx7uZagXIw4XXjM+VitLL80t93Yk7/8ML7K6T1lLAZnpk
Ipoj4kcRSYAo39RXvBDz/iZQKQF/UGYqvoYMcc6IIS74LiyUefGhxEWwo8bAIN3JXiN7wEbbYpDL
0NcZgebzB4YBsN9bkvBCNSlfngpUdbjXToX51qUzsfpZDJbKGLNGvNghAJCNbPbOGzYe4gBr8LSH
ZwF28NaywFE/ofkTHzC4BBl1cADfISdVEAGiLM6I2uJmG+OYWKSwfCZdmuZGKrSOK2VlqHEt9UIr
jxGTY686KxanCVWjf3lzYN+dRQtC75sxxNSwxDHpCnjw2dHLVlVoJGkcrlCwgjthZvAUJL+h6hbs
ngsu9AP1oFqIrQd2+Hv+1f4VS8rJMZb7fxYJaGRwpGrW797LyPX3X6Y26GTPJpu0f9kjEsU3IctE
TL4Oh6oUFiN4UQmVuu95rbKJ3l0GRXYUffBWgr8zt8+R7YvtROrRm7VlV33MaXdmgy9suv6Avx8j
3xYxHcnJv4QqMFYnknU0fzCvytFyCMGYM/lWLbi4g+weeY75o1Dhrujx4kz+bHrstFvFul56A/ZF
Sbh7Z+TL3U0CBUSAhcVcq8gn9jOvHGxN9USZI1GvkuDVM92TE0K9XxpSdtFNB/MQVC9dWB+AqD0d
fHG3bSrmL2hiqqLAbZS62uW7f29JY07urjyvGXc6dxcBe1ErdCMLihw1Ai/Z+CyFdIV1OpLrAfLe
dP2vX3wtiLETImWEXnpZ5sGL4CovzyryuyUmVDx1/YlpAHSL6+v9JVpREn6GBrYBFG7MZrwl1UgV
oz1pVvrwFj9i0t/i97o9s029peoaFnrfBjipSbXdDrq5J68XZdvJKp1giLIQ+RQCzRpBcgVfdLlt
I1sIN6D5bRERoFCZw0bXDI+/GvKOUXiJoaPzqjGGYcn7Ylem4dngPidfobKXZiCfGzurnhpxgPg8
lkzGkv6TbJ839zDb4JWNkeUCL+LPv8krTai9qRZ1LSMYsG+HSAcU34SUlu9IErOBScQRlJlzzaJN
LPv7FTXIGCOVx4R4GFVhGAp9hgqu2SC+jPgRgBw2/fqGOJmO8hDiCOeyGjI9MwJwk7Gjw+0Sz681
Ajhu4Hjy+U9MbJeJvXYpskN/D1+5xnd7nijGeZNzDJz1PbL6MHtPHKwox7yYEQ7knYTz+p3MFjIg
WFV7IUQs2rSELC7ni5qinKmd8gcOVpFRUF9BTCwIXGEcz+Pk4erQlvzSZTNSdNCs1ZkW1/VD1Tt6
gpOiW04CUK/aUej79eHgLMW1uDJ9ToJktXhhn9CX96jxtjDOtpSrbf6xS2sGt41dWCArxvCklXU8
RnVdJoIzq/GifeK8w0Wam8sADGWbAWINL6zdxVVDtfgS30b+d9y91z9a/5dOfDKpTqJVIfDUvNSP
v7kcS47PA1JaC8KeOsRngPTCJXb58P0Z9uFSH1joZUW7BRTQrg/OBxSRhLnnFghksd2eIkzQpB8Z
uMM+B+lZXdr2BIHEHFE1b9pX8oRhLfoL5F9gQT99knQT1tRMeqqO3zPz8/9WFLwC6c9QLZmV1xUt
aTox139/NzJuEiey1I9lyOQjeUbogtmuH/GpX1TBO76clWKx7CgSPXClJA8KBZnUuESfA+upWVCB
9tQ3hl5Y0r+hdzm2gdPlTEety0i4FQSRe56Vw/TogOBn1xlg7/aFrzd6KxFD10BRmk9T/s9dL6mg
3hfccxumVZUw9HRGOTnf+VpgXvRkPvVMUqfktVznl/Fwk0oSba8+7UL8w0xRnv69cqC+JUe0Xx5z
Ua6CR1heHigF1ppqK3Q4iwDUnndxuL4Iw9PNeL3tFWWAM+hYpCqWpFzo6zjUYyKX6Hsf0QE857Db
0AwZAD2lAA0Xtk4HZkyRhqLtbfi49S/9JGS4jqIOxEIg7cyE/RhJ9Diq/bwpe6HkCdotkTCb8hXE
h81Z1IcokcIla/bdXQw5HYUmb8uCwoj2z6BKYj1MNWxBCDyGL2TwbYXrylolIsA6ZBmRUwTyRcll
j/1ELMZwtQqVSoMb0xbuYbf2G8avmYEZlophRhvwmeRFGyIL8jSn/fJHzkMcbCri1tezJ9T9eeoh
y12cC0RzDa4HJ/V2BP1ZdSxE2uKMDDzf0yJHebrmYMtbQNNLoaFPhgEz+NYDyP3mSbg3Fe9Jsos3
vstLPNIDprBVOEUVOrKq9xram/bPSooQiXjSN5s1g+wJPmnsQJXDfB7lNigirB1oE5kI3lMZ7fFO
JrmYlmD1Y+aYt8E7XKydyjDkt/l79BQcsbQ3PlO4/LLSMPz5LvFNieFpIyIePeneG7EzAq8dg722
yjqRnouWuUjhmQ6T1u0Tgot2uu7tiXXUh3jvjLLR5R4KrZpCgIn1pCYmMC5fr+MLeSFAVl+2RPo6
VPx7kIy5YpdecWrS4lg3/8Gs66MhE93oH181N/dJpe2naWxlaZju+PQdVdXlHY+bqjdm0zS/KeZE
kZC1eujPpvrSNClPk1dKueAG1+f2QJxLNhRSQczI8mDu4BXprYqAs37YrEN7TU/w/9NxXGuDyBpq
AbbAsX9v16eKzPOD+YJ1wDYI211nzebApeWdqhDg8C1zYfh9aYdCKdLxTSGM+JhmYc0PAFqGLuuu
ctdhc29om4Fjhdf/judC/RR2FdIwNzIxZ98a3swBm+BCzOpMLKKzWKHjrmvUqAgzDXiNRDZvI7SO
tVB9jk4ZuMRIIVxyr8tGLUMmevor80qOWrjbnqfYQzvBuo8rCXAOa+CWqf+2i/3dMWn4a3drqfuu
8LjfTp28pO2/iCS6Se7vv9s8qXYK73unUq9iVun97FpVVJHcUdbyy2ULDVobMvzzNEBTyjhYFWnA
4/d8MKwF7Upeuzdau6QxLDXwOEGFnKIHZPHm9VRlC3V5c/KIxZmrI5IBXGL6psyBHKUYWglzlMR7
WWXGPyFc/+XSwuGv4ITnwKQXTSEsJu6fq6d5/bvttXLt6RowrhCFL2mYzsQvc8zpPuhrKZYfcnou
yYZlgokh4e4lZMJF8GL48FSlAnr+F91r9qPtZ/OIEpj4Tj6GhlBapaK3KreSbemqF77Q/LmZdkPY
yi731KoLCn1arz3bOuZ3IH0QNpY3k6Wr/701QjAJWdmXsEZ9Fs12WHAZQSP8rbKJZwbuMyEZx3rR
vc2LF2RizTxvGcBohXv5YchzaLMTc7lLtHTRqC8Nkvzs5rvGG9iwxVc+SOUJjgcOd3eeueq7hMpz
utFIYiNIJT5ZRckSnwnB9gyp+ToWJKRzlaFMGItekGeobichjfFCbUQyje3ngnbpD8mS+AiSd/xH
eq48biRfk+h8yTkQRQpil6Tp7qMiSXR50m/98d0s9c9tLSGvZ9bCabIGc2s7K+FI7ilLG1rYIxjH
7KzsyZZ/hyJ5BTxMzsvq/yv8bLjzgEquWwjz6xmy+uFGY4ibRxbF2mOKDQcCxVH+B/ZSm+D+AqH4
SqyfyJmiWscGzpuCR0+v57J4E0vGc3F0Fv+60QuH/ihQI84ke3Bh5L9QsxQJJTdmZ2i2mR+HnL1i
04lvQKf1Qhq4lUXz4OhHmQ+aMfxKy8B00kZu2r1mP5OTm1uMk6qURHSZ7K/1upFpX9G7m45RvUPG
XG4JI84aNiBUL5yjNh28Vy2A4yM5tbOb+JECa6VoIi1lb0tY8que8VeYLcM2uzvD/0LyC0s71uu9
LdlCKKBqvQ5DfK7qG61oeEVqrlA91xe+7kYyPfR8Wme5mTjI2Q3wqW8qarU3FF3dNsuyxl4DmLR0
gbjOR7fpTYd6mNgEC3tJj9jtd8Ll31OS3vGtyYggyODQP3vJKzF4qJc3G/3bDmMEx9CwJtj5UqHF
/1gysHgNMcLt0BhaNEv1G3SAcorB/y+R7wn0eaAhs4u02cjKSXO5hRyd6NYlq3riwkg8LsBsKQ8N
x187KODutWnPQ+89SgWrJAz3HPL6YBWWKB8Dd3K3fk4B0tv6iWVXWTn/EDhLc7iEgh+BmHM0GNo3
x1J5SLFgyQFv1J35Zai0MdMA502kkCC9lRVIcllZyNsnD+C019uW3HvK1BuGvG3gpOTj/8OcrX4D
hh03HWkU7yF0WA7l2VuP/acO7ZkgUSaY6F9OMF337FtbYz4Rfa8QUxX2x4E7t3p9JaTmuSXDF9oY
UWJz3hXKDB5TGW/xsixuGMgkRJAioNqpSlUb09WHvN2EIiOYhLJ5tuuiliKH/TMJbdx18Do4X4KD
RaL1sdUTntbu/oCfsfWrbVw6M64saGsGIGWaRMQAm8u7iyfRNEfD2VtLcuzPhP1JSM9FQe+Rjgin
6v5vFmXBshWFZKO9Ablb6ht3f/3uMMBlUILVJJw6GLkexOPlR38bHepg31apbRICi3pqv4EzIUq6
+m76KN2NyvZkLNCud5YGxmpEdO3JpjWRbabH/CLQXLeXoflvL1Qe8pydPe1Mu5HnqUoqGBbryiQG
rVglfXSm1n7FcTTAPTJoflS+Nh8Mdm1Imx6llYW+1K+VbrNJ2nfi5Hdad5ez86cRT0CDbqrN5i2J
RW/zJ+WGVePYFy4GV+RDHv/oVJudJzkz+FaLnwGae+QZO0Z0v40UYTG5LapQ2hudCu2sc3U8wnUO
sh8uNlKq9TkSVhgZbm1O0KxUkH/kzp6Zeyo5rdCM23ml9lZI6bbufMRkY5tS2GqQ0IuFTVnN0k4w
4RGUx/4rDVfpVVk+SfA5IjfGhlWbFQ+Sst7Y9yJb511s30bbI0yTVxFPuJ83mhKaZu0tMT8EpGii
fLIStyVKW+GMhSElSE3Eiot+jjw9ZXj8y6s68SAj1UdsD+xzh88z6kS62ztMQzQcDf1Ti5z/7qx8
1NpBkmCZLeUdgRcL/d0vCKewHI+HZOpgp6nrJaSvd3VCoK0miyRRG9ETNwtHhCCaaHLeQqqRv9JK
scigPC/pVRGge0nf3AoKsUe6xrEk8EylIUM7kUANdJX/e7He/HuAnfrkRahGB66stHx7tVl0lo1D
j8QXE703LtN7u0z4K6MDpofSJLMm7oYFfCZtdUPJPETdpdOU7iCzqxmDN2T6Sa3pCZbl8xs7yNd0
s4IykhoR3sarT5WHXhQaQd9DRPSHEPP5alZ41OaLqlUxq0PxdBsT9WkMB5fwPepp6OJcVg1edhpH
g7C+C6X/1iT9VNMY0ZXHh0Sua9/6rCAyB7kaBBlrx72B660ht5e68qaaIkQq0OZspRgX/5vsIWR/
p3b0Ds7Qp2LPJnJXK6vAjGIjPfLmTD9whSN1IuRMO9saGsXHl61Ro7XXzO3L36j8FygQkppL4gwt
IcVmysFli+fykKerOt4FDUhQe2kB+0wpyHp8wmGUp9TigUpZD1ltR2F3KSAs6/XY/WX4BK7XpNld
gAp5iA6snDcKXOl6cWG5TnrbHDP90mh9LTHEaqwo6YCuB6QGxO4yUnRKZImz8Uzjx4zni/3K5okU
jknnzy3jU4fLufGvYQZWAbymGRuJ2F7WHLOKBJTx4APX2U2TSnviPiFzSg5lxdlhCK08GvO87Z6r
oZkkvcied7+bWZtu8x9njdlxi0btpwm3LcYTaMyEpPKj/dzMmvYg7n6Dg2xMFGQVfN6rdOoIJCxc
X1JIO9GcU/NwYzq/7ifNixiPkVe13akmWsh73xTImiPYKYUBJszYxxhg5ZKx0HfNSSiOf1hDQAW1
9gWoMHZyCqwjfSDfhehSK1HYjSYFJpxyv8exVo+oO3A4qhIKo+zzt2b/kigmFWPRLunpX9rj4OMo
PCiSTRDhJ2EJMYdN52Y+nIAqcrfeqWLLXRpiafkMVp21pmyWgp/Inf1cBSJfaJ8Cgabmbg6m8nrW
vaiEMwDDH+7TLg/1RDpcvtEONGENoD0egDQMHV//rwGH3JpqTRRg6qEMGBHMPzpKiMVrrtqf3Gl1
pxIAY3z1YpFmTjdBJ2LvJh1ih+72GfjpNtGSz45x2CZVBGNsltwX2txfcNXMiFIfWymgJjhfPsgm
by8o2Z2zuDleJKDvdVqR2Y73yvbRn15a5pm6q3riAZ9jgsBNU142YdylF7K6kAYXapaSKvbYWUIb
cy/8txBXe7sY0cNL2RT0ePk5H9Vxp0wwmdz/Hf3jW5uZMZF9yCkrj4bAi9SCaQUiWdy0QiuUuMGq
azYRT2CvBXTqTeakbV9Vr0n0wUkOXjMFYaTbWJhrIyZ7QGLbZqidQ6dM/R1rEURlm+UztqD63HDW
tMRxzzKF5Kd45zhSIM3WT4/UNTAP2nF/j8jLLqigYCLWUirsqL3Hxt6ToNwHgz4cd5hOb7UsdFgU
FHWFcmQ5hDfDEVs528m+MNuSSv69MA0lO11Do311IqQ8p2tfj4WtqiGl9d0+Gdeu875pxzl8fcq9
d236p3kjCDln04hpuseQ5onLOloxzZs5G/LNjaPRdCdrdPHp7BN2uE28uXEFKmhEoQeeRANxjQ6X
ijKRV+6xxVrtTihFlr5X2/+qFADXCL6CXFSLarrzYLxynlCRsxGW3+n6JktH16Warl2VgdXyT9bF
SjFckbhATROj6vQgQG+koRe2RZoqya0M31tn2+we7s8XDTs+bTvken0owNH3VrdE9CTZn2LmCzbb
PIi09MayNvqP0ecllZ9wpTJEJwZwaKubTmtpFrXWqz4tFjPmbRoHiVa3PNC6Ot700zbi5A4+guHP
imRLJJcpA+mSMF+tI8DlKbWuGf8AZPOpE2uE+b1R+ycbzr11S3oR3VbgM9QCdn5e7o75QwRuJ+7f
unB4hz+YWl9neYsH+6wWtzeA6IWaMcFSzV53Scfe6ZTtD+7/5OHCqopZwsWINcQ1jtBi+rQ4Z8qg
pNuLPuB0nv5eAE2QadkLre2Fl7sqW8gavXymV7Br00ui2cOO6FR7+9jEYK3J5QaH7u/VJCGDC87Z
FfIsY+/yjt+dI/jzzAJV893PPD9JKPmAPrZoe5zhtqGt/gq2Wo+jrqupgKSEW8bfgRaZY1UnsUvd
69A4baMnyk67HS7OibW1D5i/c36mp1GNZSnJkQN+KMATvYufiGUK1m8R3/h6EP3tCPSbXrKVJs9a
DQ50/AKFrrMZpRtjJ2ar2LIQUoPkmQnSMn0hgHIehLG649wvVCEMsIsg7reycvrjSXuS2gIpeWa4
9VBKSpDPqcPJjFbvBT+REUAJLOzYthvFQ2Eo5PartMaCvXHF6GIuKjt84oFwL2p9/oiGyPpZOW4B
Y+PLF+vVY0z8grSlSLH6T+vAaA9K5LUrS+fhliWRELuVwFWtFiYLsxQjUYvVfxyWFrQUu4jvRUVw
+jc9b37vnjvUGV8z6G2Ib+dm2xixeLvhQvmPwQ274/E1R5KlXpzEt7HPHUUxgvFuslRM8qypVO8f
KPOcrTUu0KLptAvAI0V1MxPMKuqZ26PuMMgVmZ3n4eFdu+pka1OP6IEkSGTzW9tvXHqNzg2ztHf9
Bz71vyBIhtP1oEHvGxONmHegbfV4qQxGX6wvQBUuPn1bHVWM9f+RNL9YxP+9GrMZ3oOqicnWYpFJ
T8orEGdvAHIh1DisnKqez6kufkrzW1OajerPsgkdAkDsUM8NzVWsdZtUerPrqgc5FzgJMthua3a6
ZfwzWtE1vGdH8tuJgDUbqmn5DdZM+D5Hw+ShZBoAOlACVtNXwBXfzIsOocgKlzP/o4aB5FWWx0rA
KVuj7dhvMnQzSyXDMu/g8/AlkWB+n09eUEX6xNmBVeLEdMCkx6vlDdrSvsNb+VinOicQWh6SLI4O
nikuRrp4ZKwHoJ4R+cTqgMnJhjp8K5+JUMKjzrmlyF9k/N4xl8fKNFoAzOLyQEg5awEVuZFOv2OC
mD3SB2kGjQY8i0ofhjM+pk5uu/Qa12sSlsdNap2OBbfJuIQTIfEfmHziEYrX3KjBcP28e9S89Klo
aEXHiPoHuwn9oP+bOWGdu8uXZL1ImmYL5czltnIgm0M49sO85tNwQfcYZ2xEhasXmC8Mjd8JEy56
z5Gnh1TnXnllvacUGOPrcvKaul6sNYuDXmUKDoebecF6hipDWOkunmLrTDZea60YRSRMAlzYBZgz
2q9B2cBNNvBUdpif0XC71yTOdFRTtHi+uG+R1uh6zeHVQXVYJ4lSiLuTHwtYXK2lXF3fpcjolX9e
9aSs2BuzyFCszTLW/K2NYGy9j2WOTy602AoEkwWVeEkdpNS4s2fScKzpsuTBJim88uIJfKQrwTgL
kPahUZGpm6qexsRgljlmPagLxVk4vsyvprKdXXZrO0VeBt18a2aIkF1qYDYuhOOJsRAV/52/s+Lv
LZ2TwpTe7YmeKKIX+0EwkJzCza4RbQ9WYJGoCpQkfWY4KSC5a1WqUi4VfHSxIIHYYUST8qR23fRc
pmXr+wQSy/vqK8FXA/yppr8BLa55HFDllD1LSa3XcQODyu+IIoWmsYGfhVHSVaNSJHGTU3YjaNLV
hyyd18XHsBx2bAB8kx9vk9t4a3WtZN40z9aqIzABsmoN+OD+dPwwgXBB+mmShJiDSXuEAIzx2mi5
EsquEPXWltEYgr+SOjDieluOxj8pPoxxgIG2YYzFSWVh2+L3MARnvvlrjEcE49+8ain2iyjZ77pw
9DceILs4yENVDaPrgrhToLjH2vRbpyj8xdONI3cGRx7MRTjQBYiYnAnQgC10xFpBDZAArqpV/tfV
KU45RUaF/pMrFZFmQsToFsZYIqDxk8pg5dVIunI67R+UT/4WL37uNNLsJ7MgZQMtqxQXglrY+ZY3
0gQTHN6hQpJF2D9PqYkN4BxlbW+ZBzMMQhi5RmFkdoqfKxfxawWVUWLHniiSgK+MJfvisUm6/VbZ
6m7Ou3IBfvA6zOwmAlnjCvU+/mr5zGf7A61jy644JH3WquG5OxZpG39SCoMyHCUSpjz0QVfcaNJZ
qFyrEsHqmwkgzzvgh0dz31PaQnl4HK4LqxRjfulC6UOYBow0ZgkWs/yIS0ChgIBRLII6uGssTcNv
nQCwSiuOjRQ+FMrEJnmWa75kLxzo35wG1BpHez3rM2u+394w4isJGvm1CDMShBsFEy76Yj/bcizk
TbCIfd+9r3YdsWtc0O8CHLTzUKcqWyD61UabmnQUC1LUx4ne0VNq7rqlTmN/KN8v605oGYIcF+Lr
ClMJDS7+n/UwdsDRXtlLM+CvWrD5/W5RYtX09gj9/d1Krzph06MDcp3XVacC6Z8jjefdpBHLei9U
hyvIFh17RptjiRAODubgTOQjKVIR111JhfbMaJ+6nyXnowMJAawheGZuBcFGrcjztXn9RLy8z+4J
1cQr7vWvZXZ6sTNgfLOvX91dC4b8RZGiB2Y8WZfL+DnD1HQcFO4d2ZHE76mpWDJQ8kCMGTs1o/Ij
eNQTzbg/7QQfcdzdZVhK0p0mVcm2Kwtmeah8G3a+zfg/KkkOoXBXbTwphORGHXv89BkvCygaoD6w
3FXYoy9+CQH/FmW1HBBRTBQ0RpHT6hK53hIznXAZD+BpSIwjmNly+YgkEuRfrraFjUFCtmioJe2B
R/03ojoYsCP7uQYsltfhdsxCaWbzbZjf5W3hPGQn/xw=
`protect end_protected

