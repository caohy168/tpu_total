

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SH282qh5D/kKoH/fL9MUtXXRvtMeNFMCx2pU8KZB//alIp80aFhaRek2ArZ9/E4m3OyzHGccdezD
9RPV3AnXzw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j6QIHzGLO7FS7lF7LEbZH4cso5bOPkVOKKQ2witjsEOaHNVfvu/6Zu3Q+AfEOHn1SnQ/fLSftYN4
nh6OUS7WfZlW2PzOoY3+VbT8fL3rpXnOaO0Cy6oti45poDjkk4q456KC9MbAhIlgClKHehAMM/Xz
dXBwjzX5lqTzje0nuPU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V+KPErSLd0mzTM293tJRpGywDtPhwbpFcZGZSu7UvMpU9f0Y0w7MVPMLeUKGz1lAlENU6JsERb83
XZBC/NiiepDou9WMR8fSzjEXJLQwmOB0/F5KPwBysr/p65/yc4f0+3GVcW1STjC/yO9WqfYMYSRp
Wctdu9ogdUZPgXyikRhe+y7YwUIfiEyjdX/tPjQc6FQXgbvuaAjcRspYr4UqQ8/gq+k/zLLOrPa2
OXkR6Ea5Z8XWfQINsC4AW/1inFBDI1brpCk1OjLqpkt51ka+KHCDdC6iPmieU8o+og2+A3ToxSqu
JJOwofriNQ11wpp/fuwqEDRpbpQJMekizvih8Q==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o0P6uje/h37W1dxtR2u/dwylAXRFZLs/WhAXEi9WILpZr4a3ge3eW6J7lqe8lqc2tP3C7KTA/1UO
h9YpPWjcMXuNQo6pne77bcDMRvK28iOyktNcVxICAnfiRoW646P6EWhp1C502d+hSZ2+rZ6+rVYj
Nz2N36sqibRqSeBVsQFwN/8jpD1uP2qPabRAHbtvxP0iSI+XlbTtNUlOs3rrvjWy2enI55/xYx0b
sZ8e4SHJ35SgQbzkoDwuCZCAo6AaxgF23D3DMr1qLt29Pg3RF3XR+k0B4DKo02hh09bTeqr/A1JF
0sHAkXQznJF3j+7xWvScuMNvNJNAcOQ7SLC0Wg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xktOccc/l2sDLYqO7dioQQLDMG3llFB0kQWh1LklBEVxZ1swJ5MaLuw82biqs1Ff0U4gZIW8hYSS
VM5ntQdH1xsrsCM0xpdgjth1KtREL1xHXrVRAhISWEdjkIUfvoILdkzdjo7FfTlmA+uDg1xYswY8
jykKdEXD2preOqLNVhGQFXRqL4ycv+Mycitt6ae2SiwxLzM6Uxn+cPabX0Ak8Zp1CUkYrarO07rt
OJ3334B7zVmyBNIGCzJ9fhM/fmyMe+xV+vJmblPKRCI49dZbbAb4Qdg0MhsFs1a7R50U/J/HUeSB
Y33awy8QP+XpOjD5RxLNIVgV1ufDuos1mqR4sA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
puScNsGu6Gw7WDj51u3CvuJDM8GEP8BAoZDVeMsylgOQkWDA62HnIdByK7/Y0j2YMUoGMe5IPNbD
KEar2/rEs7TGHVgHHspKY7ptTiKYLZVHcrAMe/oBSOTHB6JNSoj5s8935QvKhjG3xtqjxPA65OVd
mg2LPA6d0uSRM1W8YG4=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fyk5FmW6BHfkBosRZf/OuykufIvfx8pSLw9VVWCTXe7xeTZYUhp6RTmSGzX3siFoVMKCE8QrT3fS
31UN3uzNq2sZjAA1jA8ycwAiFpIzNNe3cqqrAwgE6A71ff/A7ZwYr0Cgh6tjcesnkhFeDh8ljBse
1yDmANOPN3gAgmsJVs29MYhKDvHUjJRnrFVf1JkKo7d6lZQF2N2Mq366HdmYshCLueY4lWXdxDnd
n9PAj3T62PWy6zbmmDy85Yd4VHSYGtdyyHR4nfAU0dct5QeCU2B+3bb+fE5/lwUQoPTsk8gtMz0v
62uSxjgSr1QqlZ+aU8laZ6rOod3nxjo6kXRxHQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 233824)
`protect data_block
vnyVj5vuHSBxZIshQY8ueM7UxnWTM8KUsEUbzG7oAMvnHrqp20KPE8GlIet7Ql0lynVnzg2bBC3C
QpqYf3yFtcFybfhs5SvZe/C2i1PwRefMQzWoVxO1x+DDKKSptjDnpFIq4pnR+cMvaq3jrKPDvyD4
v6UQJHzmjN/suHNyejggR1nBE5xmvYqh0SiD66+b1rXN6cn1vG0BPbzUD/b5GkH7VFddjiFEoQcE
NiUhSk5fWKQOivEvdi7q8xIQ/4WV52/mVA9jQQ4vIFGFYiJxeP/ytZ7DVAYneWYuUWR4Bxgvuxip
s38g4r2V0QlXSciFqFsJ72bHgLs6u3MxCC43S8Jrt0TUD3dmBC2lBbV4fGhtzTkr2rTjFetB7r3z
7TnMtw/QTkttxw/oquRK6EgQB6jk8Cv0vLfj+2LIC69x9t6cHLMqnIsbNjKSkVs72ccem3v/Lr+l
hZXipb2/o0bZYcuKENTVEdHkjUx8JAGysvTeGXizUaW4FRYUbjMYFp2CzdEGf1bltXhE0KAsy4jB
EM6iJc7u32urHpqPyl0WJ53iHY+oSMyrve8ONGHUCJva5q+dMhcfDSXhASVIHgITFRHI/5zheaNY
ddLkBRbZSbZ6WwF5XgDniDaHg92mBU8QNUB7FZGGQ4TlRMmeubbgG2QdhdWe/5+Fi0MnsJkA7+x/
ItGqklvLj5hD1DQymBZOxxF6avGhATXztGDS98D+4hZFk0HrRwkRvz+o7xwH1mi/lGM2EVgysv4f
xYWsSrm7JRn+PnwdpGIl4QLgWQBLc1XpQV/CB4uK5DERsWhu4cXKcjwZSzmLOB7c8NtlNO7HSpZt
Jzea22dlHAucfVJ0d9dnvuRps9bwIgcgceYcE0EnfbmFHftuaebS5lKztGPA+8ItEZCGadlmEbOR
3/WWXcKP+XrWBz/OrXMFrXdo8co76GHdU9rcJ9VpIod18g3+MDHG+YJr12qeQW/tQshfLLXgglu3
LixrnEfxQkNeD0A7svb/iWCqtWsOGfy1JyMEp/RGo9j8wxKQdP23FQzjM3fD58VpWYXoV37rZRws
Y1B0lmpLI8cQOQCH7EW5Hm3DyDF8kZxUwH4V7LcHmt3C8dFfzv/6XK6BTXQ7TDojY20afgFaOL2z
FcSCQSI6w7yewiNno49CGRFbCbZ4UkPbuzEWCIHtSomI0I3kE+6UexPY2Q5jiskxsQskmQnuzDuE
haFaAfZS/kn/o77WM2/ovnQsTRU3yKySuBGwrIWFcGQvQA1N7CFv8Bxz4AnnVcQiNoYGBsiId6RB
6yu3wMmSq5nQ1IpCHDZjfucEQuEYxnjn5kHHAftLGzGsLbatEVQ14k/ikvOmGbmOEBV8Lf+azLTW
KAuZnnVkAMvfE2Rke9cIgPT0KroGL/T/c1KAzmTl3IwOO2MtHs0LZqSKBgETbo/J0OPkxaYalmmT
Et36oTvfUMHgfSV7RMWpkBrweciTgW3IqD5qK7L0CZ+MSktP5BfixQVcDj9ZUersUdYIvPTZiiU1
4AVt0IsS/hNc9crl8F+MeAam3NlMXCBCKJHW8oK9wBMeHA05mQiU/wtiAFXNl3+GFEs35/O7Ocyk
D8r6LLYZ3KNagY1olUZuYg4zci3C7uQrhpLNW5/jMgqPVsgLkmM69M1ElzQy8RcBZdIn3wdwhN91
zEvZwqQ5LPGIUAH4bdt7YJPdOwjN726yCxbwDL//GkPEo8Cypi2LL9tbiJRqzwGp8TmmUUmEvE96
FkTiWi6VwW3/2QgF/OTBMRyKMisdiMWKjQU1ZJM9R96Y4GiBsdogUGeaYrfOR/E1O/OtCSwdHlUj
kWMDDCkYrxBRQpdCKwk5zKStTvxezaCfGJAx74puSiWrfPMdP0wDbZvtdsQvQ6St+HMz7Yodbjx9
vdqv/CtMQDEAAv9lZ9wpFOhv1AonuI6Bp2xsW0oFOdcz1VikyApTIQrZNZaqUGXrZ3xqeOqEn31q
M1TcDKkn/2tISekwV3mdrvK3YErNU5E/MZlxGxPrzYMh3zLtT5pWaghWzNNamEBW88quld6JrOnI
14DIiu1aKD1jouoxuJYJ/jNN91GDbxzuCPEXvyt9NxWovTifQ6TRyE88FcyjVmecGezJbURj3nRe
jYHLRXNcebv5ZjMWWev2OQ29xqyRDIQKsnEsrmh++wOFlIi/4t+10Pq3wThE1R/rQ6NEl9uinIfR
Mewu3f+oNKGn/lZAxmNeUqkBfXRcbo0nIueOy4s+gCmD9j+QwVtZGE15pv7nNH7GAOq5Oh70xumu
lhgTD7C5Almdt+njHjw9ZQ2VtJz+d8IFLOs4J7ZCe1YXBSVF8Suzio9Qnx/0mtUs/hLcElB/fqYD
j3z3Tt39wJUtKhtEHRk8RWL4SUhXZzWsSlQyt0poa/hOiJ64cHHcIibniS1rF0SUAG9XjAYC5i5j
v85gxUb9oQG47VWdezA4T8guMJbf3OwaPXGrY4jkHsvIwx8WgMS0y3QzcpBPQoSvM24uBPQfd08e
ui4rh7Pi7n9tvU57e5b9U56MuQso/kXGs/2jbcvRxRhPbvK2aTKUxaHu9Zbf4qd0u+EGHhwgIxJR
Dl60aMN3HttwKGdjPF4koPOGqfCqrDwR8gJavNQ8SkkJEmMtP36OcSqiDSAEnpBJBeb35oiI2md1
Ff44yD63L+hU4nhY/hoOGoJVcfNzdizgxVTrZ5mua6oYxuRh5zExYqXHuyQCmDL4k6RkHA3qpnNG
fwpMXb4mYCJepanKakvC+ry/FGQ3S/mSZtpVeHp5WtvvheGcOzpB6NlZ/eFM8JT97GkULbZOEe+5
JeldT/tiZP9/xOp3/HfSlNYEXieUhKyZsw3T+soaHuq3oxQyTE5NMmqP/wBrkxgAlY2o7mtwiiOJ
CfhrVMMbFQ+l8VuFTtjbQYxwC22AXowMqrLelCN/09ZJq8qbabRXf9wKOkaQjj9FC232hLzaFQFa
0lswHOhdMTFaogBU0BHtkcJ35F30rmA3sntLloy4B0yg9t5uQGfVV6wrzRb5nojJZlumV00oJ0nO
5abkujMx6syOX7ue/aC6Zqs6t5hws0RUwpIuPseJJYxS+bScWxZPVTKkH11MQqhdDPduXFymzDqj
pGHxsaQl2QflPTAwAacKiyuCGoW2O/QQfoJQXEr2v/WQMz4gSukO/imr5J9ctKcDrojd4jh3W16q
PyZFJ1pnqcwSSqfU4/SAsIbrMzDdjB+kRivXz0ux2VVUFl1m+CGbuGBp6rPF1hHLus+LzdNUP8AS
Zxse4tXaIFRp9TKNw8ak7AQLEyVx92ZhCix4fLNEom7VjnNhYRzv1K8V6lnOL07hRi8z2ExgSm6M
DngnjJL1768nJSaVN28LOiwPPDfvj5gHu1K1UUk72taQ06bGSQTKLx6cY0/v9NCpRANQNQygVvpC
UAK4+CMrFg2PDWuvBiP+EYENdZyb9C/1aiissRtHzqe7cJ8wvW2abIpChPC8dtV0Jo9EYBycYcuv
V00rnsCUIouY/KBza3BIDYiP1o54hpdxknop23x7P3zNyaU4tW16MfwTj8xt/VNgdbTW0lvQB1eX
N2xzmMx4g5o7IMwu+28LYNe5h6L13EV2HbaKo7vPp5qfxxMNlupWj0x/iqoPs0g6zAm1RX0tcs3U
yNXR8vrRBIYHxE7j8lfth9+A40OLVEoWZZEYNGFjl2J53xGCwgezwl/XObaZmKUDd/LXsClx+Zqn
CpudixDqQhSTZLbjYECnhW7xcFFSdPKI9IxUf/+8yUrawR53ugpbmgHCu790w3BaJqH4OUd7sFjL
E8Y4XuPdlMiDvCU5NIIfM2+tJeAS356SMcqKY+c8RBTxq8EAd4CfePBlzrEkZ0TvmbvRA9dL1cWX
7+90mKWcv6LoSP9EDthUJ4dVttKkn3WdL/lEAEpNoztp+2fBnNirriQjuM4KRd4TQyc5LPBvwLfB
OhqsrUVt7vU/WckxA5Ikosa/UalSTM/yKpmxIYIwt2qHG9fyaiphqwolYGjpBXC4C7Vo1ufq9Oez
S3UC72wwBEmAbzdAG/sfrK+1OdlTVUJwRLzsM1i1/ENbr9n0jwW5ykMykn/DFJkWlfsmp1qhIhL7
aN8lzEVRnW/UkEcrM8Bv6OBAea54IgKhnV5XTfh4mwx8Bk3EOnyoMP7t6d4IlHQpfri9whNrzvj/
kbhbZpxGwCHgeSg2evW8UyhYAdcbWsQyCROPl8rx/5XxZPbW031Alx5E5ZIZlfqZLp9wObvqje+c
hmJ2EPfvIOj6Gw9Q2kAenS7mpAock+qFVP3fNU+dzlB9VYx0xJmqniIw1TTwObHv/3xijiWoMxQB
Vw3bQYHgs9pQL+5/zxYFTsvZeuhf2c6cvB11j5txgSjKERDUgm6lr5RiZGvxyK6sevZv7l8JYTZz
UWTHVTGKTa2X0Kg4LHHvU0LvDfY5M32Q7kSe2SEcvEIvxtvxrwAh+RbJoBxcQbY9jckxXDE2UXX9
N4B2GncLQoKLocvGeYavSczdkxo5hdfZ+nl4ar4hC9VNSQow0qbwP2mx0z/UE4C5n2RKsup+iWAo
6KwXdok5lzrGD1bej04IOkES9qGoJpjkuoMTVk+4QBuKgqJncXTmTrxIFWVXfq4o0LHcL4Rw94eV
l0m1ya3tCsaYfqMN1kbLmLhkYtccOcGsux/HbO8kZa6obAqrK0ElUNKWjI3hPrE+xjWdAWl59UFC
J1mrFf0crJzIEj+QFMkzFMAQ0KVUKv+MUhfdedPu9xu9jkFYrjUnEkrjPv3ZuThG1Cc25gUxDUzR
eRZM+p8AdtOW+jIV4yGAQvuhAm5IlePcqBoKsEPhMzVuk0SReVQa8CGmtfBltFDG9StlmybWfynK
bsRJENX+lEEgM+meYCxi5fY4dmSMPPA/c+nyBChkbqPNjWWCzdwEPUgrGqoNhfhZABEhLfJz2qzb
ODsjIaHoS0BrLH5N+FFEiV+eI9hdVXfq2SL+Xq6kKmp0BE2fu24+KffDDXhn8iCh2sJfKHXBIL7B
4vjynck3NfrO7YrGRAIA8JAp2L6Ism+VaiRWeTET30Hr692b6bD5EJ78Ev6aVFo+fyFsypxFnFx+
Mmm3oNBBHL+tM1DmI+UQB9PGdCVJvoqWOx+6qehuGGEhKykvJGUkLjWFpzqW73M7H12MIxIdlISN
CbWy5873cRZCxCc0mVjSJH8f9wjF8MJ89MRvwQLrEk5f90fjUtsC1LUvFBoEbC6zjOhX5pDfK06X
IJZ1rwzp+wTrX6LZjgbYLBp3msrYKynTZ0JeqH1+LDxNgS9Dvya22oyeah1TSj5GnkWIPuMhZt5C
wTGbScDajp4qK9sJ4vlCm/l1t/lnJoeyJGyhi3hab6Pp92Xw1tm4mNNWCXT2tUGXTwkhz6lSuAMj
nUhRFo00vnNl1e8yJkUi7BYa5R1rJAgwZu0/metjsQfButUskQqMEn+md2tcLMM5Y0v983NAkYMs
I7t3GpW5dTVSOvPYmLqzQHBRBb/WkSHUQOEwWyFOz63zBHbOTr109bd15dQtUFIW7Z0oY+SUOxnC
IoRJYhbOYyO7MeWa4K3wmr/JJBGKk6u+7RDBzYWy6AFgkIrbCm7Eo2Z4dhtX+FIeMHDLKSkkzJ+0
mEGWHWolmZMH5CMs/+ISp4NHZGMCGnEgbmerI5v6byr0FJP1pSfL9S+em2Uu9VFR1hNUNXTTh79l
na1NT3eFU9ipMRH9BqwCJYpf6Ww65jCLnUAPLDFSh2v8z1Bnz9n3y/z7gaSlYW8Cnf/pRUpwiFaY
sVzCWzcBHdiPOpESyhRR7Z9nmciE0++6XLNpk5TPTHiatISrdM7WnOMidL92byf4wmXefb/ArANQ
nefLexViJgjSPK1xZ79K1mUqDQPYLu/6F8QVDF3Ex5szVnAi67NFrqo5Pe/+PoCMZvVtiNqbpI34
OiPDJXTDMMochTs1yBgsjFSmf3Jfpy6wpito0cgomyEKaEYYCo5rDOszIpt1ZaIDaLNF0RzH7i4r
Bhi/6X5dpdF872gsi+4d5UjVBAUH/Hr6VmLu34I9Ck27tIxIiRyk9Nf5SGngJBqyvvMWdCHa8gkV
ZKDVHOvJAYLcwCEx4PxXD1KowYfp/sZUwxtVvBrUNSFMT4kGm3eIzPz+khdoxJHT4n8yZlteQucC
gTu74wARszp20ZQeVHxiFDAS5ugAlB4O+NIxujEoYj3q5mN/BkScEnicRi6ffQ2w59Q5uBh6Nz9q
irj4UxEGO1RM8Dx3cC6fzvjNeL054qujYOboy9Mx5t0pU1ThMhFxn4wTO15cASmwcgfP5X2BAiP/
ctkPlKInbsZ9WQ0tXs4gG0NZgI6TefiWwp72Z/6qsZirECzMUixvA9rb9skirx2TjWulpf22k3Ip
YkOf0bMEgyXXXk2uydlwOpaA2XSBmdGqkEeiTTEeFUR61Qp9z9uNsH768AiNkyAvOBAWxP0RPCWB
ekRmgsPfaauskDXm3F3J0zoHiJbeSDjvSX693zITo6zE+ON3/d79R3nea3AFVMZ+gcX0tAVEsSmE
XXiHLmapQ03AuBGuxb23SnMdMntec7dNKJf34f619JcjDJASudLJa13tKwrhtTt+Psp8ql2BNu5s
2ZpFf2KY4H2tZ+oQAzgf0UQ3A+fzgP2qBpMHIa0xYs5Uz3swV94cud4TgBaOluYN6Us1OHfAGLKQ
JhgSbStfAPh6cfi6VnxgqTu5jVz2r33OjCE9rkW0Z+1C5qLzf3zcyn0ungwi7dVRs70II4FJxysb
4Gwq+eyqFOmILHzZWFJy1qU11n7rqhFnezHGLigPeraTMUwlAZtVaflHMSnkUvrpGIfIkUHbkM/D
5/xUpw2MwZhgmwfhNE9Jav7PI4ZaLXSxPQobtJpMSbVWUd062Gk6pXq4HtcIkYpgidOGn1a/S2O3
gPuP4THWoJBblolbQLL3hKDCJP8AziaQT6VHi9qHi3QMs0kqaVL5VyvtC/UKzxBx7C2HVRSVXFNc
oyjDJf3tkpd5ukFw0hS2nxHVxdtApmGDP1P63EMbZKw97ZIbMPmEXKLIub9A188p0yxS29aHFnX1
8QzlI0qduO1+vaPfojjvPuaA40+Z8MgQ6sD0XPx5NrvYf+Q19oumppYX3JI1Z97Td2f05fMZNhty
nDkxXkNgYwpXto5hjt20IJ9hGexQ/Dg0BuVuMwItROCw7nguHfpNnmcEU8NFBpAyt+drcGBPwOxh
bEjGSoAJAPMWMM6YTj2+DsJVKV9IOV4TjkAug4M+YfrwLqEJ2hfWQqLLRaWQuhXHfhQY6GT+ALkI
zTU/zfR4a4TR9K8S0l4cRWALXkgaXBoVvhSMxQbk2+OYAdeA5l4538hL/PEXlYLjleRmnjPi9jv3
N5bRcJgVHCBwQLsi1kUArC5xbPBzrGb66PLwUrgZn7Vpk2dsFKfFqmT8yM2hJo+9woiY41SiHVuD
3PuGcC9YPt/uYfrxVmFmOhirX5NYPRNPuCaF/ESWuDoxGXgJlNhnsE/JlRR5eT7B4W+hpr/NcLWS
UZ7aseUKTatgAM40LCLNxwPfF4el2Kl2KT96o1lHXAwF1zrtU2AGwb2BGodMsu1vIqsWixrFxqnj
XM2ZOGCUCcw4fJTHajiOGk8YGiAuG1+hlyNrrQegahGs/d3wKyvUMCSQ5FcOuukKLMLBraa9xAy1
pFdy8NmZfW21+4U2FZKyfYvmtj0rOnhTTs3s2wqiCNnTQh4pqnA1xdl8yL5oniri7ZvmD0Lm9R/o
ODd73HuED3kjFFdkIwykcG6pPttX9ZhDat6Bdl8kFMSBwqmDRK9ONzKz2wX/hoxTyRhkwF82ALQn
iZzmw8hnpzOmt1UkG1imAsgL2fet6l/rgPb+St7SulLqYagOYJ6mVTFvEHzgRzcr+IcSCvXJVmVI
eY00BPM9W6NqwJTpOGjqsi8yA5FVFmVj1KyryCcTXW68xCM5xw0tyvdhk1/QIHNQjfpPd1V3vY86
W3b0g3GMpxlM3TsMoaLKt6ffvNdFfbai4q5mk1ZlbF1mzTlzL+aEf44OK1M6CGwiBTAaAwHzGAe2
06oqrsqNA8dQWLArW8NW2FRGZBKw8ye28/opGDVXO3qA8oD6qxevalJloBK2IBOvcD4Wte8L/tv1
VMZo7RC972FROLSHymLogY+zH12FJZEuJYgP4+S+1MqfBJN7aiR53JL1YsYfv40VLoeR/pG9DVPd
g1C4fXoYKJXayd5OX2TerJmc+MtHkCTlWu82bY9d7Q5pzX5WHQM74FESjmyb9n4IxM0ZI4XNpqMs
O+CkpSdWvq+GUj0zOxD7kLLB7QVcuQNokhV/U8mDLvtsxicldd7Vt9QZDL4siKf04gx2qv4N1jTo
A+epv8O9FHznnYd8JpMJ8R9dh78WXjEG/xXJ4Fz1BKMHo1l8T9QJ/yC2xL8baSz3due005Wk6SZm
6Tee5Rsoz9mKhXsETlUXYWehrQpfi+KD0uSN/C8/th/EB80v9kpsICncVrB+zbMyBc/1fx2mWdRR
qLycIQnkF1PiYeLzq1BoMLriz79iyOTQM89cM6E3GpLeJugKZfpO1jJWNBqBoNXfNAShmeq16OQ1
IVAff2S4KgAwrz5t0JW0xCwiJGtRdsDyNp6/hejd01e2/bp/z6/e5yFUbRnWEYrIhkJrXrJVtXli
Qq+OZEKoY1P+iiMFsqHHa2DnzxJH1R6zby5jAPCc02McmoGpm3kfNY8F9PKP+paKuo/xFcAqMXhm
C9x/Agn9nH/cFttRoQ76ZZxsjpE7eIXB4XIO+PKMhzthsSn2ow+VuXsFOVCuTJrkgldjN1kmvXJh
5p7tix6Y4dia/kI8fPmV4MXW7YqyFPNJVibFrtbHzqw8DIkPrJ+D4DKtiXIbI4EBPCyjMiQOAJHZ
W5tggoxAHQx+K5mUJweNZKMBdReNdWLIy+i0+jGlwUHYkQ4oD1WPvGLH4TBOKSd/Di7b2LYexF37
3v5D6DI3z1jsU8fRX3Y8jvtYHh24xmcLBy3SumbTpgv61aL78iq29FPDmjLQvoVaV4SKz3XQ9OLh
z4sjc/HCI+fRfEuXJ7EdYGtXQ57tljoqr+lu99hwDmATH7+sSP3kausMDZPvKlsurRFd3VmOe0CB
wwUoZYEIxHpywdw1bEmTYwhiDqRSQnta+ELxv9a/79RvDT4P/5jB/TC1xqMG17jRgqhnK0BEvhRv
0n59oTHyG5DLgVinnFqnOT16SJlXRRKGSgt7nafz/oT9Oitffd+8slBModWJiB7rfhhheKYbsMxs
Ks26+qQGvupWm9iqEubYBaddol1W8IF2/G0JeEb1w3+Bgsx3chFvHDRoYTmao9oW5xCIuagPChkB
ux/+A5X89RAAVZ/mJ1z+4pr2QfXnmdebSzl7vL6i4UbPqSRud3/JDKzGstpJ1zo18UfgqD4wPz3e
rkrqt/LQ6Khf9RgZmT00lUEqwDdtSGAWlvlsSPjdcCMpKnEOw9JhGKh9o1RpQEaDZv1goQ/Mv/jo
PyXAwRc+kUTdoUjyOz0IMJyUfJWhcK4oVoRdluY2yANX0Vh5Vr37n/tCgDBe0wB+XBjztfD7545M
qQ3DKlLAbjPJdRz6mfkML1eY4KYRXJso72LsDQbkJs3RW6PlQmvwq/ZrbfBW2vp46LBaVMmng2Qb
WLty2Dhh0Y+WxSjBQo9m2+cdC4bJ7xRgUulN9ZvonbEuZ34ZqMJLEy4zO/XNs45W+ZKWT/7gSaMZ
IpVqti6MZQF4TeNlYgpZbXHT8VyK5/K4/p3ge/XfdGCpjlPMjgPik640pRKBB4Zpiq1TTcyrB5YM
HYJMvs60Px4P0nPHttv6lmxkh2ufItY9Il2VTFNsVO+GrfCbxHrbc/xFD3CO1q76nH9Vc3qvx/hA
iBxCxXFW4BYx5aFyZAnJsFldcEX/iSleYtvc/6F2HiSxisyEmO7ZOgw/DXFHCulPHmd8MmNkqxFX
Rfds5ayZQdUXTN501c9uDsPFcRMtsEQP+S8+H3hIFOBY3rsZP78nDm9JGjODbjG9scryS/mJcJFG
4AcV5JRUKffW/HBwHVLNCr2opIGlc7kLsKk6uyXvrwzrfvQdp1luNqRvihK6HSVRRRyBc4LB6Xfh
zcotz+yQuYx7P7r0tVjA5XPk3ZkNT/zsQ2UkF3ejy3GsTVOFf9ifm3DVsPI0zj7sLQUC+j9NpzJP
rW1c/+SyMvL91w1gaxjYhlBY84WujKRTqM7rK7+bd2CwyGjSqPIyibEwRn9Tp+rY1o8n/mMm9u07
ey3Bk+AUt7R/0Z20od4bDKWxgY8Ty8ocAvtVlL94Zeorz/yn3Mg659jjScLLF0qtkBVBLwvkWL5G
RJg08FaLriqPM+3bhFKJNKyUpGk4Fmf8wVj6zvX/0BmTdKzlMroX756k6PcJYBp37zNXvBDym7iP
hVNSoLIt5DRIUItXnsZyvL4g+yDhjBBw1fOg4j57/9upatdNErq75omhKkX4CU2x/dOAegysij9V
muoHYAoRL+jZ3r/7W/6ICSPiEVvAg8zTNkdnH3xgTRCjJUa2dB8IWKFfQ6dzNiHOasbHpIb1nwbB
Q/1hM4XohSQYgD6p3bj/u5WhEApoQ7mr0LGRKM0lhHTLIkrFcxbs0aWZWj7WzZPSxl7bhvSh1iPO
A4LHSIae69HW7jAVX3XmsmolmiWjPmefPorxJTu0WzUKvY2O5ydCkm98BqfhayeC5ndyRfVovY6D
G4ug4XP5ao9hw4Fmxx8bGz2O32PnrFJqQTXk1lrc32wQr/b/J5Dvz4SVMVJ8J0zysHSXoMc57LiG
kCV+KsWUsR91zGD98+ojukxOHn+ZPtSol3aKfAB8rfUqUPYL26X+omw91s6jnADx0dr0j6vg16SQ
9QoxwR5t+uMjh4mfqmyrn3j5RdMJnAgWxrR3nMePDIqDrbT3lZrcGutQjtiFxXOwAy8sBQvEPyi7
QNfcp1mzGVjOTSsxD9gEW9CNoEDmmgfETFntvteEP9K8e0qXhr4H9rSjUe7EKu+gb8iEXyAwdP6x
32Hc57rUvYf/whA5B9OsnfuHHUbYo3LaX55C5Pp3QcitJrb0OnyVztKmon/7P2L3oLFXzdwOxo90
xDUOtyAFqhvvaLltf9Wv8XGoWJ9Sc0Fgt36yezI2eTVJ2jJ7x//pYYeFs78XTP2MYgiqljU4VRxF
4UH7x209NT2AyLfqhZDBhzfbNZC9sxg35+fz4dYLLoeHcacr3L9zaiBqijOiaX6JZlRr5ZtZErsq
4pXC5aHgxN7FmrhaSsvT4WSvMVLhLqezf6hezGFYRXpf9460urCBp1vHgrH55FsJUsQCNQGDL2C/
NcU69BS+FyCHFdP42JoC2jJSQco+WlyiBDJvBofKBTm0E/c2kUtduJBLcn5wG3fqMt29gMPEyeZk
4ENvVH6gASz1AxETPHHz55bEZw75DzdyUWXX3OIZZjwdN3xj1paLASbOYbRg79Nd50OBouB5Rkzj
RW28ayiINrW+ae3kXDsbePuedNTBPtdFPw9YdZUX5F4gm5bI0OqyCQV3ZsoWf0GyEM7haNWhiKUG
EJCRuK9VrpJpSrp6mReRasCTw+KXELDIbOrUJ+I/AzUcOImEgWzkEP9EPMhMe45cTRooPVZPU8iz
IZ0Zfaxlw6YvI5olxAeICAPBzJFbQu4imJZPMjuPI1EboUbRaksy02ASXziA19hzKJreM61M2J40
lnJIEldrcMt+vPNxGLuur7Z/+zB410j4hn1wrxRYHmdfzzUI351EWvbWnQBkyrDoYaFvWb/YLRon
em8NOOXLje92OZ8U+tQhqbWTrzX3GAQ9YkIWnI3TSsXLVr7gkRA0GSIFV/opLGsVropVv14Lu3oF
jYSoYlad5f2ad9XWMkRU7LH53iqckF+Mru6UgAaNaz/X2EZlq4PTAYWvJY/asx14o44tyE/dkeoq
hjC5wXz6978Httj7KFg+3OPTGt+UApihdMimqaL5Hx306spyl76ZgoX/94Oonu43InSMUbqGUaJN
IK89L2spcTXHpIPQSwP2+ZnvMLW1e1M6Ew50Y7DqiWnlm+ZEO6Foc8Icqow5aV8gQaT9GGzRSJZ4
y+mi6VBW0+6EeGK4q5FK6uAz/dd9Tb9KpLMSezkwkklbkK2Fwcwi0JwFrvlYJSpHKNsUfvBR+qLs
YcxKJXRUIaaOcPEaChslEEpHqRuE2w9bWCwsPkaWVY4bRcedDumpvDXtIoY/yWxRn6OfHZbOGNPj
1BaPaupboiNMg6SmsI7HKaK3Rw9mz8kkYic6XD33zo36EaRP+fNQssU0pp4VhgHq+OzE1zf0LO6b
Y4Dwvf7E3tdQXJy2aOvWWKWgomrKwd3jXHujUoyqYkTGmmEJVbBavVmZ25TRhprdiZ9ZF0dxNLRn
pbm1WvgEj+YTPEXKB1BnUnU+pTGTpvVvlSV/kNyKENLkkMQ5ExgPFSjIorYdZzANCCX/FZXOKuFR
iFGJlFyj/i8FX/wEBHicy8SX2w40FimTw3CmxitqVQ+v9kh9Nhwr+oh2dWO63x9k6MHT6LcVhzgs
ezUxZej82DyXLMpzfu4qkbKe9tsJDwz9qB27gxxADKqS6SN/ypAt1FDqqVSbM9xR32A821Z+9MyE
BRD9jrQtDbcY6howJftrEMX0jqHC6armI18NFNUU1GD7YS5zR6HwxuYsbTFRSqTUesbeJmgbZv2R
cIHNM1jQlFA2wG7a8ZfwTLTtkalUdg92oiN+KbASsB/4Iz7B5ebUZFraIQrs5liTwHQ60IMlRzLG
GGwIkTarUa3i3Ax0FGoHFwa0VWljM6FuIDnsRhFDPIFr9cQfjJamYhZlynLJwOPwki3N7JfMNCZU
nXoMISIQLCY+1m+d3BMgyMOUwuQC7cj3KzPzshoNlxubYzo//2mM6OEBWpaRa+kkYcddM/PzfTc8
v7KBWHfs3NJ9DEgLQMGS7ZXyIGE1SVk1uJw22WJvjTUc0nvhqT4LcXavoP6CDdDMt/GD7YLeTmuH
LTYR+AR8jSWRsEJlJSkwManMMtE302gAoTX22F2xFm1DgIyo/2tDz14OMFTXIcX6Zr4jpd8sYOtI
eQMth9yk0kZMZvQJ3j4tmTvBWW6YWHbJ9jE/ywB6A/NemeI1c1CV1sU63WHFA3Z9ezznYh6YqfVn
uQF1xCYY6ivh2jExG7gb4eV5mpIoJL71H085tqeFSjD6F4sJNyX3Fhjg1XzcE2BOFpGfF9wP5cI4
rg5CxSyVjoGhv2QC6IkTWbi7PQWQVJ9nKsI3m1WxpvSwkFW59kBfhHf46fWqg2ln/Kjvfw6/8Go+
+JsZPBXO07T8yV2infNLA6VWs2keiX08G3vcHLsWkRCsiqvkVdR3X9VJZR43GFXNPT8Lw1nUIAFM
7JZhwKNZqhvzGYLKucORMIPYddieCLS6EJ+sfuWYMznbiFMP8euosjyqKR9k91Wsw1/9i//qWZW2
u0Y4RdEVsTeRT5lRwb+ZI//yWNZrQueIkOZwN9Es4srhhUs0/qqgKznKBzZYpnHdHtnkZsRVHsD0
gvHHiP+Rb6bYPCvluUH28MCSiXbxg6ZtEIJGdYEgC/hLFq6xYqHKnGWEjg4mibhn/0JblDGd2E+K
tKtIxabVSKCGUtQ5tjltDVvVL2n7WY61nv+Gv6bBqkeaALY3Wl1TY9gDJUZ2P4yS4u59Zr4yrhV7
bdeIe9laGfcQr/5avj0aZLexWpzStl5rrjW9XxSq40QOYxdBpq36LvbiiUU0nHTrT6uleo6lMtFO
lxYeIA6GLKc8iJD+6TSedYwVn8eqxjS697F4xbU8elP9cLiQiosobM7qYVfmKHzNnyHXNpQnjwhh
RMALgSo514ROMgNKk7yg5Vxrj4EN2w5jsepIApy2Arg3YN91nvY0g8UeRRPCy5/8CudvIGpGkQXQ
QmnowPpwRX8sgN6DK3ehp3Eb+TkVG4Km5PeiVG8mqp82TMkytHCs1gVp+WAQU1uTLBSJmQeiJN30
913Nenf/CchbbUpXgnAt8XEzV2HepF7f/8l1NgqfcSejMnRfvCJaB+5MDJQZ8OwJy4VzwNELpQEi
VZPmZ6nG9EtGuYYyWf+/ny/UbmzUKXEWZNGm+1Y0ytRLiNsTvzUfJPG/axNQcTAyPz9xXt/G/nXr
xZDFMhWzQ5JikbdFM5uvbCF6GdRp5cWtsmlbIoIc9Bv3jctHXahVUZQ+Xb8ysZKgps0rKu1INshl
0nDVT+B6dhbCJ/8o/HY7wJidl2JWMGNXWHcleaMzmvtxtke7DtZV6OzJpHI+KU6Fh2J2ZpfD9w+w
DPLEVftZrSG4/Y6UnKt7oZrdNveFQ2z0ycoobf2PrjZ4QCWth2HPwx0GcTBNyn69ikOlHkZWgG2O
KUsk3YFDzigeKHzWck687ngn5dlha5QaEqiRNRBxOhZl5BoUjNK+ELeotCfgCEg/4NBwwUv2YV9B
tdHjX9pspfcVuNXAvZZRb8PLb7xrCECrlo1IhSmhnJfMYSaVMHn3kPuDAt8gWpmhxEUC6LOtBUeA
rWefwQmv88cV3xPNec/AqQmomycg9kSOUdJrrpmPNxznhdWhlIMBkmJx+3ZNT6PJ7ColvUS/t79u
4guaq/JWzS+BL6Te49BquxpDY0mhl5Lo+D+RfQ6mjE5z8LChCNYUO2o4a9kMmBbJ3mQdideu0Dum
J9k/p/VYhEeHhVekJbaMvSaFRbRWHMBq01UKMlLYjKmgJPFcZMraM8OsNY+NkHEkDEgsFQ4oJ1iN
y4JSX0vlEGuGmTcTacVTq+fKEN9YFRyKJZtNj/zzyOh5KNmS1GpzM74Wbr+D0mwF4LnFzFgvFCaR
6uc0Z0j7KJmv196PJsz+aWZ/F7K2geRwHw0waq/WrfaseK5S58Zfa+5T5ffoAGCG7IKR3en948Hf
VTY+3YJmrr2hk/57gg+uKSY4dMEcqIKnZ8/Sq28el/sTHartTaePMVURTefHoDQv2n4M4/sWUARu
eZE8C6wmlu99dmioSSWMKcvgwS1n5UOXsi+ZonapH2BPFUS6F4sK+P12OY3XNTNRy0nhJxzXYTMP
0z4NrkyS3CeSAX0tCwKkTZYXcBMnKognmRhMkgBgr4/v6mimOM9mpN/CYxyw4h0axnVrq0ROVlfN
8uCKBbba5AQBO0cA3VLMTWSLAIFpI3yUZsM70xP8fkmovCCchlfGX/GhJGz3J0kiXznoUFkpmwij
xgWYDZJ2mtn2xJA9aHqqJVGSHrfl/wDYXEd8BIYAbMIVYIXgpCwcdPjfUjaGx7A9cai7WcSsSiE0
7DTm95extCvNR7qbWkvvbCM+PWWpTYrFcJWRsuRgoRxw8EXGOhBJzUlzDhuJOqcq5U0Vqyk6eHFp
OhmpHZyfxB42t8xcrDJKR8lu91P91MSD0ydW0pZ6UgLJwHPRtm7LprfApGTAhzuyqpkiRq7OQjhv
d3Uvd0LItewN6NAFiACzzpYMKrt0TzVLP8NS12eHWmRuvhND+t8Ww5aEDnhDFpJOutz3Jbm4UQcG
inHAhL4qLathA7/Ppu9mAk7xeXVJObbl5RhHtNjfQeKgso39JCtZalHYbF/LBcDP6PLHqVbyxKfh
6J3Np2MJkQRrIjCkHlNado0KJdN6JNo2AlXFDhYBFqOlI2UwJA1/Q8zdbMJg4WqZwxR9iFrKDhHt
/ZScplObEVW8EKqaAcgkQ3/qRhahihajZ/pQTsanGSVTLkomkam+Q7Qh+vAE7ORkMGFK/gTKJm7L
VX13x0tLlXs26OthDCEPXUKtaKwCTmFTcOYbFBN4aECGLFpllG1cJEd/Vc423RkemITwRr/XwlGf
lV5wobLdZa1uP9gCh/0Usd9b6K/oicZjT3oRdWTg0FD4/UssxUgiYt79N0L28w745TRp+lEIm9Um
wX0RuBpT7zxh/ykSlu61LDsHIOvTpZa2K4rQQt13B2P/FU15oHNpOd60NDG/aqQKy/rqDHR1Dmp+
E3Gs+L1JLmoXGtbDduZmLtDDB6Xmnu8nNSYYApx8afhzFmep9awHiy/DVCZdIvowkt9sCHMOnWOe
og1TblHx7Yk4tS0moikRRuLjMkTGOyOt6yIyyUjDCFKoUQlNB714AnKlEDasglUQ3yGX3BUedlT2
BATpsEVNlxB3vpeii67WLm6WOR2cTPfmP3giuRayMhZm29s8dbp0Q3KH0vMPYeEQgkQ9V72s3X+Y
Vc4ikOwW4okGDlYj8adAD9/v0pcyQDzzIvl5IEJwsF/M1fahsMwowwzx1PkgaFhv864l13FUgLRI
kbAyzh6Y9LLRsSMdfDQWS+Y13kaOBZmeb+b9YzAWWWlmqOMQyBZ6VIc++78aMz1IKg0giHOE81Ov
XIZEqDcq+xUeIwYul4jhoaGurRqWhA5MAu75g+4zXpRUGbfuNyJ4L3gXQi45/f+EbQSzk9E1qZ93
KE9zEhQdyv7u0xvLPaQT/fw4ot5mcbMT/VPLExHZqpnCxWcEaLvfqkUn01LyGgjAtalRCZE6mD1e
Cdjrip7UvAK9r3eDwiqG9PlgiVvQvHgLz8XXZ5wmc0NvFxEVOjRQe5moG6+HRCztd9VJ+k6+GtYp
fKtQU8atxW6/0drjynHHFz9/zOiUSs1gWmljA5sL7j261HrIugUBsvyjDsDgRuXatewrTMz6vZ1a
1sOA7LNmhws7e1txl5U5F5jYpcQU2OSbGy2vfZ/MvRfVvLj1xej/MF6xsuXKG8VcT8b2HcSYtoc9
9+ZPIT16h3f02WxX62L9Tr4WJKApNiIJknfPze9/CZrUp7vlRxp6z8oqJzBZJ05+rSKTF5mjv0/4
Eil67RXAbOgl2AWu2eJSbPiRlnC4Zh140IDdgZ8Grw8igA5abzC/Fpdc41eXR8vr/87XPs9fehWk
vCfjpJ8s9s9EEN1eCIrhJaJPmH2JvhtsUp9T/1/p84cEbl6TmIyoLs4IcTtO4xy9BfZWjQ840PQ+
iDfGNI0HwlHlqJ9dCM5bebHINoBkJZcD0gfh42zeNDarqbhilqkMh4JYCBTpiuCMoBYgOBbEx7PJ
MKJ9cK+OSBOiIkeWalwRLYLOPBi7XlS1dAoRiKOFdQAgdxzyaEhtjf53RC9jSDeea0APIA7/7dZC
wkVGfbLtm1NlC+ZDrQpfGf3oY0fjeirCqq8j4gAu/MvqrTie5jppFRMyHlXpvyidrTzJ0ISgsbBg
YLHaIxX73/naK+0EHC0eM1ZhBwlS29Q1bXjiKj/TPY6KcWFa77SvV74zrIAEDir8lW2WQiDdAMgL
2e2opZEJwRNcZn3fTTFnvKklqJ8M5h/mTvlcdaTw+kQTjNwC6nooQwazUZrYZ808g64misC+WtXW
pfbjQ4OOim0Cn/b9jrr0WSJT24ChPs+fboT7eIUYyr2lfKpivUaruv7+lICT29ifjqpN0SnEh87Q
gTbq3azdITlQ9mq2EheHzDYrB4dHuLXPagKSjQyxJxoU2C7+Ab4m96pEqwC0xULa+ZAaf5fnGVWN
qZvmyqawjDqr0ppW25bXdTxHQVuFO68LrI0WRoNbvaDXtGkkmw19HQ/Z+e5r3sZH6T9endKdXtpo
ZZMCVuTUAQl7IwtuGUM+khUCRz46Ym0qGwEaTkFxqHAf3Hp6ySe5U7PtKDmSMq9KctW97HVo3c/M
hshO8+ap+yVHp1d8uf4Lqmvzn9gs9j3PQBWsrhpDkGQFCEG1PAkdazDAMLa5p/AUYI6cvWWrRxNL
uQa02D9eDyh8ftAKFp2Kru+SBncy1rlD6Vle3TIawukWST1OC0awBJbmCMwILWrbkERTqLkIdn05
OS46+w0CjMo82WxmQEbaNNlBxD3y5q0MJc72fozoDltyp7T1x2mbqbU31IFR7Fgv7SWyZxw1NsNb
MwB4h3fax4YWjPMAXHrTIk+3Ps3IFzo/uM96GptbA9I53DspQ9CbuCJI2dlaWt8GyQRp8hpZEUZH
KgMqtFYOPwoqTJjaRKGqD1KMVJJv1ciu4Ka5jYNKjiKeqA+SKzsvofchHmy7W7JPIBfTYbaJxEsY
zCuVmOC+f0W77qBm54NCXwH2O7Ny69ftoMNMSYMoFX/Y+aUsDHztJ53HBVtPig98G/sAzckDhZEL
XmLpHR3wxpLP8h2OKdS8BBy/b7Xl2PIk1PtyC7u+optT1cT/Py7t8cwU7I7os0KJ2O6Z7dlvmcDl
FiJ4XMyWCawUH5xm566CWV89QRH7G40PxVm4igaQ1FUwZFEotUQT37fIF7GGZSU9W/lnN4CAXH8+
RVpdi9KpEK0SbjQiVSddB3LuTZPy3s45QVN966Y9Rsx+khTap9A7e16ui5FACEU1d5D63YRHS85i
a7R2ddaRS9tlq39xoO8xP/HXNUj97SN7Rw3MLXCx0hK7jiqd7hU+0i0z04O/UCct/AcKR4CqvCbn
WfbYNFRsQ0E6XV9MxBfXHgfYa91BAF3oChvKwKZgsfp672RFd/+d4V8q1HD1KFzTENNsn9fitpsD
SMDpwornChgEmGabiPJuO6Vk/ziYuar7aEFKDAPmUpmcOxO+cQX2UllRifKCCyU5kLiypcFPBtFX
naKizauQ+nhkf8AGXXv4ChnlY4lNXXs3fvMgheSPiGOElKrmCM5XzQ+i5xBMpy+gOrmX4Ma/7bXC
/Fdqzg1grXYfxMS7w17/4fjHZ1LpqtcNHYHxnDb0dRdhR8umH2fNEQyoaOWsR5portODK46epY1I
DpU5Tl3zWeepR/W7UF8KWTGqyyARZNsx0Rbb7iIg/NKNtG894/2VjABNa5h+ni934BAqUxmdUVX6
D1j1lQSBVowWPOPeVrRg6pAHDPcnuMI3Piux7SzMDEYY1d1bWWA5rDbhcfrzs8YWsSc4FxpzYeFr
iiyc+HCOjarqJfgMzpjVapRU2Q1Z4lhrHrN1/X2sRgS7I0m9osxVjJYA2BuSZVatSmr7/1Drekwq
xEJk1jCvTQYjfrFUlv/Y4NwIp1uk69eWctdPOcoWxHou41cdbS/fAISaluGJoCLTdq6N8n1+93J0
TR/jMAhP6KcEHiQC37zl3rC9Z/1XcfA16br095RJNut3BcVFgRs2LHHU7l9iKgEksOtxpObb7w0Z
gqa8kuoiLR1rRCW29XBu+QS0/ANeI1yC0DWGnXcAL1aRoSPXCFMLIwrRQQ9AOkFu6U3i93q/xmf+
LJFvyktSp2k8+yfvXTu5hEVqFOfhkeqRNNcsz0sdqJVD+JmCi07a5UrPWC2f68Vxd3oGQAh/eg27
kfJ6WHVAB6xH2QOZ4CPaLkwGRYNbsNBtnWFjekwYVxY7SKnNHbYyBBHOT1Lz3ej9mcGRX6y+qHsR
NmNPzp5WDX7BpMGDySAah303/28S0jixc0B4ppH/k6rdFLKTGtVH2nzPDEH3TaoHAlJ/2MJQYWaj
xaIfdDUByfU4Ye2+1+Wn+LxGxOHol9PChnYKFh6KRhtZo3XclnIOsG0DbHMlmFq9H2Knc30eXW8P
/MQF6cO5O8dEKff4w1KG0fF/gLatA3NDtae8wwfd1OFk1+ZIsA/Y888iAwP8Pbltr7xrJjHXFXNK
aMTxD26oocTx2FUxE0bUer9Uib8eQJIeiIq4UAJeodK9VVeELq7iTf2RXJg+6KdiVyGJ0rBhe1oz
RZd/sxkwtyg0yAVW79M1rShtfU6AEDeaX1RqHtjL0jmnXXHbLlWpPVYWfMI09/ICYRenurx/7Jcw
nAXZfwqe/rc5C7rpZfm116pH7yDs0HsDaH3ED2BYcX2C4OIBXsJ+TiOa3v+rq/ieAqNTnvUYGhSV
Y022wo1qqfMCUp/Ko5Qbz32wxH4LZICdNN21a5/Nz6TzqrCweoT2tqnbEAGucDrrjrsbK6WJd6hr
M1hvBRBCHv2teACWokNUNUYbAK7tFQ/NRAtjLLcyraOzdKBmzAbWy6aBvAK8wXjs/isguF012dNn
j8+RhxiGt2woKqweo8F0p+D0gRy7Far0XHInpN+8dCpeTwfD1xfx3jl0EZHj/EQJncVeo5fEwJvR
/rOXr4rqe2/3zzOe0mORxwxAWceK5xZ59lODoUzF5DqaHZnIDtabPh7Su5veQstiikYi7NPUxKDD
hiPqOYawG4uPmjIDBwicbqI1bytlhkKdsPIW9aVdagPOl41aPwkA8gHFUB1NFfE2HuNXw0N4992A
CFTGtjdmWyPYF3jOm8TorZH0W7+OO000NhkFvt35NmV/CeXscm32NU3lt/aJHEta3CeU2tv8UyL+
ujiVL55m4SQ9BriiJkG41BMrcuzPybKZQb8NuacjtZY3mjIup48yKrlJwqwRbKnZyPHw5ryh1BpJ
2rn3mQ7gLZuY4NWbph5iz5pRvdr1H5TJlP57alayZJPPuE56S4zq5TnitO5aLTSZi5dX7g2T+GDG
zZ1Lbjgyo2FqPQwnEHtm8zTiSewn1z8iwBMjLLLeKokts6cMxShHxFtwNY3KPV90Kxix2fT0sC43
XSPbkX/y/u2dT+hFLgtSVdUWwwszwh2NYsPgT06rCKFw6tjRnyOqQYQOStNXaCVYS/Wy+N5cN70N
jmeJYQBpS4TQPR6Sd6L6DNZ0SWrIFTm3Scpl8xEJabWSs4JIvcTnhquLAsqcQsXvQqsXpX71V+ij
0tJbZW837TPl3vzWoIyiO3L3GfNAXFldS5Znbmo/UbU/30BDzEdPoEL/T9+HJsoPXNB8WeZoR8Od
bVR6dDLvLGL2/NvwpJtqM1m/otzGJx64bb8XAqeztmGsYow503msgPXtbHJ9LtEIr6Wns8DbTg5g
b0oY3oOfHRx4R80fkSsTQ06ozxlx38Whgw0pS5pJxI4IRgPdGsInajragrkjLLuHgKdxKPTo9rAE
RuGj6tI3uIdLXJHyq7kI7R5bBBTvcbkTNnYFiNI2a/43MWJ4SXP5teeXNsn5urzxF4f6OromTEWP
mbPEY7dVT/3kiHjTuhFgce3XqM9U2WEPnya+Le5IwQtmDrGIxWlhihXTWqlezpO92J/oDfrZm5Q/
7AaTGAyjZ31m1qdCdBA3L6gD90ABaTrjlG1zppxAABA8FjI3jcPPjVQZSunHwIyMQH8RG5cMMSQe
qJ8kL/93T/o5VGwipAYngIldLtzm3ia7ukvMhY7C8GooCkn1jcJl2h4/bIwjXezeGJ1YwXfV8hbv
Ut7yjKFqrLxR2Bh2yPvkI7SY+Wg+KqeL5VD8Nu3slUaERhOL4NCQqvbIsvOoYygvfLbXixKQAMVJ
JnkIqF4rp+I89hgCoP8qMirA3Mboh7gKNoIopa0TIxgp8x+xgPFNS6F3OfAHQO7/wYbzpxOTdzga
b1Oe3uLlDppkvt99g5fFHb83GD2v408vh5d83NKUpBfjnpAIAvkxIUuP3cFm49cUasUYY2PPNaVY
ZXzmgPw1xNKjLr9NqjIQl6epMkhqsGRRkAmv8hlE4Zx4vnvhwahMJaoDi9NB8Y63wm/8b1Ch7qPA
nsaSULVW2NeSD661hhPlsj7U8Rc/FsLzd30OptNB52Y7Y2JhDE/lYd+y9yTMbg586aTmNNZ+8tKc
hxivXwLpV8AmXCkrePRlR3kF4OY2j4OQC+ur26rsV5+m3DQR+o+X9TbeFjKRZRagMYx5GPsp1s4x
y/yPsucrxOS0dvUCzQ9sfQWznUIeHEyToIVIKeMjigRROyrDhluOMOtSmqQNHU1JI4Mh/Fqp1+i+
J1kyFIKm513+bOomNphK5lalspP2q6SufSX4q57poshWsV7EpC28W9BhKYn69IRlnYEHI1GRZ6jA
JbIk+1Uj0wl8nj4FlT7S2d/+xVUN3C3vcrudrSQtkR74EslhioJL/5VK+1FDQ3TYFXr32Ezn28RU
YJLzBFfq267CRP4nAxQ6X134kToN1JB6A9Qguv/FceLk6+Ef0YjTvrq48jhdBzw1QgBrIvv/f97a
5Rfi/sjVcUm9wphkBpPmcJFNgjevCvOppTlN+5pUyTKTxLNP5/ENEhzHOQ1lJQf1iQP2VJUlPsOd
1tdWYFlhiX6GxJNj4BeXI7Qfq2dx9S4GYqkopB7dH6dXDdYLWSPBvmU8MYlhUqBToyN2CWD34ecS
Q8vvRgw1NgGjJtueWWJJ/udN1vHc9mqonZ3/VOexyEwIail9lRCUV6juHxxNxqB0zVh11BalYrzF
p1vvjbrujQ7KZEOVOsnkdn32zwvUXehRQ0epzU5a5DoOnuiVDSO7m3gpJWjRcPV3+FnC72R1sra6
wtS/rgaqnYgQ1+WXL/GqxFjSLDv4Ce+/YxuStRzW+6Av0f7DEgCcgZbsN7kUcvextVv2rB5vGo0K
ZxV+YLlKXfF4PFNpPxc+CoF3MfqQILTN4DoHE84WpxWuH7nyOOW/FXb5X4ZkrBETRfOaonO1fH95
ymqjWq0VRFDWmIUe9XGQf/7qwD1IcEHwVrBfZZ9wHnbJQy/o8ylOiuE7f42yjftjesSzfTjQjXxm
DJ635ynt+bLGja9Dd9ZenCfWHpYslpAuYVm7hL82Phglx8pPn6FReOvHPG561Ky/c6lv3X0OXdrf
Gyi2rJR9LIM8R0BqiWcIKiLOc4QnpDLFQHBVyL8WNJSIQ3TScve+PgrMjyIXXvy3s0bdJdoY3Vyw
WZMzY0eMgLF2e7GpKA2MJfkpLxqWdBiYZydfgLVhnbdcz0r1lXs2hjQ8PLSf1xWk5dXbjWLlEi5a
ltRdQaFB9zBI7Qa4Z5nF0r4wy4CgTdSWgUVj/XgKznBmQh5Z/+rOQTOQmy8gvG73hSqZkr1rp8/t
6mQ9mcVwfsCPkoCeDODSglJwW4LTSdUCUr46bNLIo6NkmhuJFrduqv/P40OQsQK+6Il2qJRaRvF0
W2Gqinhz0o4m/cCb9TpG6Js9DVR3qodtY4qa4lcFIElW9QwVpGdUBKaGTlnR8DjxozebLVjHJs+R
ds2bvzTNys1M+5knF3ZeS00et6iqHdt4DagHBE3ppE43CvvmHf/PY7lAH4sE7FnmTZwablZA1PC1
f+4Vx1pHjGMQrjEidA/6YlIYDh2Uy2aMpJZfkH2IC5zyTBAtNirYVFXyB7YsxaZmCzoXxbZb0/fG
xpbcooTkm1id/gSwf/5Q4Nxs5yPV136A4feRPcw4DtxMQKY9a1Eh1khQXzqIVbOkbsQJdXnZ4mCD
JPahLeaYy+HpJLtkRvxhooYlxTg5J/WZT5SB6SpfqfvbT8+6YeoBbpYVr4mrJLHuxbImS2Fm9/UT
l/Pqd20WllOjcFm+V5lMp8PbU/a/+zDoFfUZUo0WtMKBzgWKf2D1v4qNsQxOTPkrYH8vTKEIRFP2
TkqfP0cSDK4F1e+sAelge3kWqYLySgLSz7VNyEDAPzcwTTmXN20rcVTaKGe5Xnx7TugWYAXRHam2
fEI+wUUGosmBmaLhFa6y5mYSsZHlA5b2a+VeL7CD5ANQzUmlrgge1z2AvN90+EkMe+Uw3aKXeaZS
yb32abUVskU+cpg8ER9SxrlNrx3UfcauSHsj7Mf/gI+JmlLrxMwM+o+LqjcrbpgFxI8SK0Td8L4q
D9e8MQdNzhFO+sZyGxUjDHTiH02Sn3gB/K0mEuWQujhEhG4OQ5vxr5MtT20/uw/UHox28m9CEVZH
ny+gz64xh+LDZ6f8wEs9DAPTyfzjUN2L5+AZhXhVRD7ef1GV1b5KiCoIAQKDeFLfjZ4F0xldumO/
oty2X477I3gFo5iZ170xEQLuXKzNktc/Jirs3qyF6EgxJa20/RFXoPKtPqKIbrnFleb33gT2z/Bp
tyjIUAU5RAIokqc7tJqln0yFm11RM4oOYva/VD4HmvnjiatBZjcv+gZpNExF2LiJGyDhjNpS5DQu
jfUkEafxWGpeQf/gg8Px4Xwrh8HLQ5aOM+EI8vEvl5/Olqk6aDwC8EA3mXbU4cUCBK2EE8bKq+hw
VQjN5/cscupzJt3Ojkn4yhRkKbPBvY10jIjjDXaI6lVsTOizpgnmE5DN49GH0mxPRBVVwnQan5T3
+p7+QNbrw0lUOOPDDXollJykjCyh1BN8uyBB7IZNoGqa5+PrkwXEm7DYksJLaS0nEWt51N0QFaH9
RZFphkbJc8uUuKWc9IJK31UKY83/cBOmhEGod1UiPROJixe8WAExrFRjH6Ceh1mIkl8cIyMnMhfq
EhvrxLx5RNbiFw2JLfnlUJV8AcNsRlqeOgNIGAPw5HB0ZJkq3XtuAZ50Bu0T/u5Tj0SM41q+DmJM
Tze5AwzmrUtKW24bxCTMPkdAvjulkSArgr3NrUJb4IYgC573zlHQMgtqGqTFck9KLt6GzvYGvyLf
iKbAH7h7lpbCP0rb6GfeNmic/zgQ0EQPal0a84A/zl47dtP17Mlw7dyUNDyzIiR9v7cSvei7Dwj+
9Vv+miJL1dsbO66hsZ2gHvEWMh9ktNRd+LUlO9RoROu4ocfkVc2261P29NfOqjrzMsREWnn02Ylo
sGjTdfy+LGUEpU/np47Dqa4DcL4pMzpIOC0KkdF3FFBONZiyBFrLQ0dQPzvr6CuK9OB6PcmrL84E
6aFbZoYOvt1esKkwbEYZVdiSB1n1dz0HwffZtaY0LJUKBTdghlInwbWQdtZxA8uPSKBF5VH7wwsQ
u74yPOWOGDeFJV0n5qzzbgcS9CD5USaYeDJAtIeWCwoFh2Slnx3AxnfW7SKJkYsTewAUbGIVbleH
5qbXxUvGoghNx0JTrdsmCe7Gs/fhczmhOPA8r0WTSNk0Du3Maa11+4PXlPBfDoHKbIdko5+Pxdhm
6rm779CuuzB+stQuvLnyFaJu7YnFADqmHmc1hd7Wde3W8rrk/YzSuUYianiQbJ50Y+9qvu0uO7/G
auWuMZWTfXbiwnKmD8jMmsxunUt07F73qbXz7aihShH3g2pc/nFJ+QrYM4u/rdIVhBkFfNX4j1l3
srOAbJ//hpNUqG4LLouIbJbYxxFBaHzwrd4DDvw0Pe/lsEm3tXmENniIKxBROn0F4jIJ7ye2Ck2i
uVnYC/6K8OyLAW+bZZS/JmWwK/V7nU0Q5CAorlooi2Gb4AGmIV1H0HSlgOSERB179Dw8AEzu9Mby
O6CjBXB4ZWvD96tMnkwisUGhnQfmaJxhTL6Y3yosj8P7f8ns2D0nAWjM/fcsGkeu0aGQXOYvcpwv
m/kGLcfpNzCdX2Q1MJb+hm9M69mcVBFHTI+xl812mqAQVHB747ET3IQ9mBLhPEnJ0NRFmOLTHrd4
UnPIjCZQGwHzEZo686AkJ5n4VkyZCtRIE9zqpeIKztshwSh43NGc7CVoZ5uhsgvD7AJpgYbDr7MJ
NgbLi/bXxEXCQD+XJnK45ATnL0XiQPzuABGcULgl6zNP/IgHyfQGHQI34o9G51UAb8yKgRcNvKV1
TGiWGR28Bk80DHvO73d8sRH8CN9aoDVpcCFjQaVg0kKodZncMWjm3qUmP+Q7bvqhiFZKHiafMEd0
A7QabGnjrKiCjw8dNfqspPV0Fca+aavE0lQrdSKWrfWe01IiskCvUbfdlRYP91Wkq5eEjuIcNipF
jP731VdRwX4m/mICUkL6trqhsg985REYFqmKAZzzSRLtyhvds2FwC+KkW9HEuWjNppQZ76rc/Zxw
8X041VdCklQYqVY6ilI2F+TBG3d2g3ElXFA4TMRJNUTFPQVXKrt09nrBPN7nSedHHkh93RxsTuo9
Q3pMaRhId1eUdqWuYhd/Bbz5wXWbAifTo7UA0t1dMnZQjuRn6LOLJILPDEXjEe+7+KCPwomOZg2u
NOe1CXEMs0kVDP3Q5JVdE84RQeAIkcTROqwwSV9fu3nXFNpgOBGOCae5XIEZyWuOzfBjXKcdyyGq
69B+A6LCdy1xKFUWebQ37tsxWRb4cEDHuPFJP02ApZwH4cTU2W/z5h+plrxoJDJzzZJ8B2u8bfQC
ed1elsstqFtyCEV7sylphDqu+Iku8VMczbYfgx/sRtNbgXGnEAm2MgHbNcZvHwjff8V7OF3E8Dys
RPt26xx7LcBzkJm1/d/rU/zPxq9EcJxfjAQqsOPXbAhz0XC/U8K9qFNhMamg+jfMWD/xm3jTgrje
mUZglNbrXnKUx8zFD46q/PhG9g/JtgZGEVXYvB/mVhdxpKappXkNaGH7zcv5Qyvqif+QzcCggnbJ
C8JlZdLeN/PkRAlp7xSUVK6B10Y/jGAfsgXQpOM3jNq6Wh6O7vJ1dBb4TqRRfZjO27nUTwmUwvO5
dsJpsMEonTKKBTCgN1ZfgSaj5D5AJxmrpFE8zHfYfd21LDhrIKpqCjLaFHnk3waOJluizq3eghHA
C6GdezYNZfbdIUerYVgvdvkVhqGUMrDUESyCpQ4KISA6IEui3bCMufk5buVim/slWIDy/k29LW5x
yUHbdSxl3Qwm9eLmFwxDbdy5yWgVHvKSu/9VhSBItxD+GLt3mDNk/wjyPxLIn3eVOKXz55v/TvwN
ISzds4Xr92ye6pZoekQB7+OwKIRLsQVFCfwFvESV8SVo9EgV5TDqpHcoIeq9XgnCWZlamEYjkdOe
tVycVngbUi6EhQXOCeHCpk1IbfniENaRZR+G0Uk4/3I9ZSucLUn9chlh18/zOTNdZY3+sVZgvJdF
7SdLb8nrBbXUYS/5Lwa2rRKLNIJBDnde1Za6TNfsRpUkj2NXKJCVp1OvHMjIRvYyTy+t0Pjx5BpA
vEJfoXWfVFuyvkmeGQy5D2Tr6tIAgiTi+9u4vdrbTgl7GwUfCr1gGn+hTjT1Ixk3kuWm4JY9be7a
thRcUz/AF3/p2u0pvf+TBbqGYr2aSCgsa/tZ2aAS7gczPG/tPqGDuKCHnDooyiENW0YUbpsx+j0g
585hiR9FAHB/eE00RzH/msgsiJLx2TWH1sA1edk13k7XKKTZbDhqKcXrYgtaAuHDD9UZ3iZzvXyq
npx8/E9/omrs/+6rl7soVNoNyoiBVYVwjpaRgso8XUvrpxT7zGnMe1og3Wkjl+mqcR5omhcuAt5g
GPFAvEQtmXi4WRkWAtNK50+at1QWAt2ajUkW0FuI0fD9tpIFZANtoqapbEzIBajRhe3lR7Yn5XqE
Yg0H665WPU9CStbqyNs9U5GebJBM5Q5k8OSVVwbXUKmoS+8FnBQjXNUan5ZjXgtP0hyuDZ4ys8C7
OCdAXWZ2vS1G1NbWVBbWllcY5U9Qv8PJDCtOipXeDwwhlQRju3waQRGdkddcWsYafBSApAPbTft9
rP5Nq1tGLhsCkNsgWC4Q/6qMowZFTa/OPZLT/I72ftgTjM+RUgUULA2DNQw6LR8lb1+lRrc43S+R
tSd0twrvpgMDW1C3E7GCjUIumf4benxZ7V+3qiF/cFx0Gm5wMcuxgh7FqvEwY35GHctN8QXOk0qL
B0ixhM3O41LUE7cwVaiQJQVEAtbAl9Gdpd3FMmlcuSdduXNxTROncpYTOIx4PcQXYGEJMjHWsP2n
wbkw8MhyTItAk3bvSDhqtE3QYl8pIMGijkzO0t2GLfbQQ8cnWrwwJsvRodAWwLg/LZHXxoSwZgA3
Y1H/oQRiZY89LbLk4sBwCmVb0ED9gzeARDrguD9gWRB1Hjd1Nx0k5/26mgKfZu9rcaPIUbSdlph8
MBjcHrlpoYR3vcc8y7ap6Fca8Elv97Wp7okvxsCPSWQ/LWwPJHyQXX1XQ825btM9X9aGRWBG+rRx
a//XaTypXcizwPlxZ4b4TKQRdMGUL8pie2I53iCcZLaSXPhpXDSfZm4hsECJSLNlaAyS3ow1FLwM
JaWvmmcmgstT0Ioo3MaVtcAELjgILFxXv5pe8YdIoHh7wDVhBnCYSxC7qKtC7qPhDx61DscveGoD
J2iJM9V0k1033SXE3bnFwwWnSKYSjOhqI2FmHJKYSOjKTvIs1tzgspiHZl24tNFUDMYoKyzrAkIq
6OiorUDSOkpWVARLTqV92BY6uIHvcX29zDR6zZw8Qe10bvkTE9SYHFZwGU2eq1610d5a4MvBp5zD
xtoZOZjEfvohmE7zil8vh+N4UWW3LU2IFxjJzmOO1tE5/3nIhpmYGaEAKkt1Sj7xl0VA/iWYtFnJ
B8unMdq0JCKiwAPkfoMl1r/rfMLA/CTmLpX+hKB+CP9WCFaOhUgR1c3wQjOh7aX+eja1rxtemajf
gjv3ImeTlqSh5MrVe0919G70nFtChP3eyRyLdZ1AEQiT7feR1SwqZiVkpjMNGnmYCxFXww+ia5SU
vCopRAxu+tdMnfwoL7VRmt1R3z7LNKPZ8o9MjQ4rWLEfmuYxgNk/S8A7Zr1drylq37kl2T3wljdi
p7ltujCP7zjaPGdLnPm5kwNYuLRfpAvXiBys6gJoPI4onbob+Epp+CMLfuWvtqT/3/Y3OBkoCh1V
PGOWuM8uvRxhSaJMs1cScXBD3F8lr5WMVNI2CpxafJv9aQQATCmfdWKA4qZ4IQ7vJnazToASl87U
oN76hbgDfaogvvwRcFh94jsA0A4RIK+8C/8fkjhV2EYKAc86GesDjQBu84wBUc0xdNMC8tcyRTNE
BdXOea2WtLSv1tGwyCLUXahVjQF+ms0bWh/+EiiLA68Rwu116chaZb3U9kztgBuzmlCyR00fGch4
nnctGAc7dyoLbmjq7UHvnsqAtGwgBJ0cl8Q07CvQJ18stnuI9+y42e2BOupWynG4ACXWdRzYkn9r
pbZyMQpoJjOVhV3o7OekE3zJaSQ+G08MMkmEVQ2jplDueFKkY0NQmbm8lWNoqn8FOp4z0To2Hna1
Rqd3yA8ncAdKOqSjzr9myBes56FMA2P4Dg0cSiyTaKpT98xRdFiJdlDS6lJ/O0doGAAuOYeifjFr
2cVTc7PDUQt4n7BWB2SWIuitLRZRGZlNr5KD2LtDf7FvKCpSajnldkUYMhj1RtFtxVuCO+5ONpSU
yybwG0+NygM/xmaeyFd0ExnmHPD85EMtlF4K1awom6mzPola4SVQZ0GJ3DEZe1VimxvNj9nSMyo/
wVvZ/Vh37ajLThHj/E7U7p+xAQ90l/Lkd/8cQS5Pv+/oVceg7Vsfc/6vj82GqnAqY/1ibNpDyyuB
evUiwFkBr4BZEeKjA2FV+wg+fat7XIOwDx6lig6TkBsNakIMRO8XYnx1/0oBklEg2T6BQLtEl4Jx
SLoZNRONsa3/yJTNd8qBiZRjTcf+DNWKkj7jETXYnWD6+gpSQ5MMNSFLk6izhky3ojmvhfH907u2
pE0sTBNreND8cuUeSeWJAhLoVM1rhTrjKuZEfafceM6rodEuJso3y2nlgkSxY0ej1chnoFBJaLLX
DEDe5PUpe+9ApwYPw4KW0MN8HjFXRNHyBzkx01gmEPVu2sfVKpFlUzejJgOC841i9sRVAKtMaiWR
pMM+S+IH7gkB/9wqbp3diUM3rdwDC9+2pPK35RyxoTVt6EA2HzEmF+wni9/djHSenS4wIYf6E8zX
3P+ufxajV/0FWuQolEEFeKxjDvcSzzGDVHqQ5O+sseI5JOEtgb/ZWlvyAYLNoLCTyKweeKxNLQkR
3jRnPY1nYmCQHncf67nejpM5pA4Rk66Z9ZRpQHRUq9aeZOdD4FO9YXv6B4skVJeGsOAITH6X+SkM
7ZYa1BdZ72XjGrdMgvMECfNfMf5FXOJF7IB1EkKkNZro53P9EkmBXQ2MABQT7RiLhlny1NA8A0kH
sbf9ogxbF/nhejA+3+f4I3yNmlKJEFqKhZmK+u/nkOYFAmBqy2kmmHEPT+/l9J5Rid6Tyk9QAVPs
CCtTaYGilSzEKjvBbthr61haPN1w4LX3OcQ2qOxDM4nBjJQlhd52QO1x6SEUNwkjKoV86YkBbX+4
6h+JkKGyw4ULxYnFdtu29lTOhBwZ8Bn8ZNyGP1KQWTFAyJp55WC2GRk0/jMXOmG8R41VL6phsalg
4Zs/p7Muuf832/1OpJM7hyWXPwZDHFm5Dso40RxnSCtZdHmEcdsbedsqaY0dzLw0E3DeCk83+Ur6
0xlJ2qrwOeAlMb8miUsjz4qBKUbNmIhYj1UCc/82oMhvX24DKfayJOXn7/MrvJp8sgCM5BrbqwGI
OSOpWqnbtg+Asji68RtDBwuBTF0tvWAH67IXg83V788XmlpaXU+1/Kp03rChUfV70U06TP0D6ANu
SuKW7sMQvjThrHY9aW3D52bzYZpTsZYqMC1J8tnz1wyionItPK0Qr2Bb9W4CuIPcevwV7dSFSglM
YoMaMK8m2HFmrlZ3DE6YhL/JEL5LVbrwYxo+BneYGhkLrO6EyRAxxCdU6u7tuSQ0O5WE8EMSsSl5
/3YBCq4CMh7U9OBhbkxV5YOIB+NgqEG4chc6xc2hhorzGzOC4gzTciZBrmaqo7lzv95BWGpfoMu4
UIEyagsqAkPS7r5le1+ZWoAeZ2WU3oxBs3+fisAQwl9+Thf2tjhOlSRv4B9DPZfrKQPDhfQzPmBI
iWua1yV6mjWb8MtWy43bhNQupLYlATT1zj9ZUtp0FMAskhKk7jUY3AQ5kl9n5U0vrAtrMF6tVNkV
rXkpU8Ad+ZoGCS0H8j9iJjyfTZgayYgyfRNPh6Fh8LUdtTMBkHHpO4Brs0Y7nmlF0kFpiJUrraGV
lL0+IKHCANhrwgRwag6DMTqQpdZrOTx+Vii2VcTF9CWkjdq7NVcwPxrEw8pXnsNwYFFDMwMNDaOT
L9z2QsAs4DnaTw5EXHvqKhtswXLeXYFu+PRIiV8bJMrwCvDl0AqrwP6e3HpSvGgko3SIRuiCzQkv
Q7Mjn54mCa0el2TNaJTn3O4o3s6CaLnKMAg93cmFG92PbLeg4xrFyvvy9YdnlBAsChpsuD1To46/
3oH3Yl5AgrfFAESOK0VFtwkLaq33wZ75QxPjs0C7935ahuLH6hoEUB4maY2DtXvDtecTLKMCNVSs
WWy+Ya1mktIwyI9m1WVlSqM6bAhTINoeosS2QiOoxg6GiOzpnr7sOxgNYyQxchxzqET9X1qXGlD7
6j4q/zQYS332Oc+HBtZ7RdCEpE/PgQFQrjJl4VbIMvTlSK/isW5NJz4soZz9GkUW0MIesyX+Hoxl
pwx920pq8ca66rEyaAhhuWRC1MwCH/qdyQhFcGdqRXwdJBSwJDIdPj2PzM81hclT9YPVJ9oRCkST
581+WoalBevohydKCddFAyP4wKi1lS/wzUGWgAAUnNzHMjz+LpTu/mCx/o0hNHV7PuEnTs7Trx1O
mrPAHwIQAd9hCVb6DBVW8oJL/SCUKrQ4lbbCF3AVdLjh6pUbIyLwq4sKGU1KoV/thxfsq3+3H9PK
QkZ/zLeWy6UHpX2jqy1b8faBUwhLQVki5TyocI3X124GdgZPml7ZZ/ZY8cDsMjl7uZ1gpnbmSIQJ
PckpCWpf/U/J/7ahRnEip/z18+k7v+caZ8VTAdzhiIapIB+3qcD39sEB+YamHPvB2ix2LmainVEK
7thii4gjnzkTUnjOgclGeW/mdG/UZ2uTTB+0AjAZ4UiKMCeamOxwhclcDl3jwfwWH/YqqN54tesd
G0uhgE8YqCuTsiS5eAhzviIIO4SYXIHoZJBliEdBWMQPtq2GvP2YP7GtfKJTxnBOgBSrOMgs+m/l
kAVV+Bu7fQY3OiBITSWyc5UgJZ6nZYYhDN5DNKBpBYeGe/GhKVep5D2bSEkwp6sRSopPgfjXAg4s
/eFOQGewGBaIpzlsVyTYrl3iAB0k7bycAOZZy3hAvTa0XbUkf4o9x1IzESHcqa59KbBoVzIjkxNr
eVvPbRnUZKbfbS3Qus8oLJD3t1ksm+LwGdvPucty6O3g1zBd2oOJYchA9Y9e3v7f5tFd5LweNy5d
TQgbwZxbZ+ejSPHDRalPiW+wWN2uJCIbdZZExfqvFrHoOPY1ASjkwLI2W+C78RErvYGA4o7Mq2zr
kdAB33USlUGKNmyOxLHJF1QrnpEFPhKm1TztZ614Ghq6TEiUimjudigFq0++ebyFAI3+jpWzteKe
Cz0lHK2VPe68UINa5gd8RgpOX8judfACdHru+Q7ZvUDlC9RVwSvyAzFdq++unjnX//FwZuhZbH0K
qjHRmKp38LX3KcFGxuzvPBCYNhP9KCZgLyQobEMeOjowT2/0xn7uWHoGaGcGfKbBIlaiD2LlSy9t
BsyL7qs9wee68U+thTgStomFzDnmQXn+otr14VOc6Qs/3fsrRoH+CGWOVZ69MeccKLjL5E7/2VoA
igBpjOhQPYUqZhNMATyJC0vAb9kr7f8aT9qh02XOdY33A+YlMEGx0xu2Q7nCt4a7QX4WiLtV89A5
NOQxhPrDBZigmuATcnlb8EsiXufNVX6Mm5GxpiN4E0/MpzhGSPJ5RXdk7qwv5DW1euzDWh6P1C+P
FBXR9CLyNtp9zmDg2b9KBxRVLZ9ML7pZspFJQyyc8BomqYQ03dQJQ7N6cPI0OBct6tHF0nzYpfId
NpgTBqFJ4StqUMpYIWbDfMHR4gekqQCWFoegCxL6SwXB8uCwMWdqk9t5JUREPBhzn7ZzSBcyapdb
pEI4wmYJWhcp0pj2sNq46Dr2tYCjIMTub7xQ0mHX+3iDbiom9vEeXViqMoZE/Ce4wzVh/QGXQox2
qJZraMjy/Drdltr/CIGlFOgP3FiGTC7nquBlz8PQnctnba07QsiBaBDB8xnGcrsJmG9PoPNcZVpR
XatcKG+YG3SLFudityL+Mhv/hEipRUZeWwh+TVtCFOvPBoY8f7TssfJIrt+KqoQth9v39dTgoBb9
Xe9oEY2a2vKfYzUTXRy4nT5GHb3zc5inBCSTcGP6RUTX6pI02zCDq2YblC0SyO9ID11y7X5pQeIv
B1cEVUHrHJFxVTCfvFgNmgex0NnBuirPsxfUvI3//CxzYPyHBTMMq0IOjmVENQjwBrhAWjwtUwsX
Zas3fU7w1YGs7NBIo7tRQrV4xVUrKn/ADVYWp5yEHrJwEzzCumKccV1tCinB+9I/1YmsjkbIGu64
ouMZkM6ccQ5UN2faq/hvqiKrRkx821AxnYUGzr5fSkXepfwmgvH6ZiKySVbpKERi7uJCZ8M6ru8q
t62JiqWzq28esVo0OzzRZDeAuKUOiOzMsCkszCFmXAVLtFPXKRbjkO5hRz7XZyXCk5Wc3EL27E0C
tS8XqqZOby8p2A+hgZxUnNXfPv02GS6clrqRL0Y4Ja6S7JUvDXvaH7XpWXi6m6URlyCY8fiOg5Uh
h9cp961OhpO5/tZsQOPDSwjXR9kc3HwAV3fE/ebJAzzTqV1GNPrhzYNhLVCZbG2Mnz6AqTR+Eoev
Lw4NggDuOeDjsGT2cpB5CU7noQSeDmLeFHbAyXjUUERAqdKuuxMn1gmvyc25XVWVaHRJmMNDeziQ
4KEShvz7fPJphGqWu1C0vQeiUn4cZ5a+6tyK68bXW71zrxGjul1PFUkjpy+iwN9UAVk8XT/vy1aJ
z6idHHlqwh4TDYUVEhOz15mVNtZA8TKsGxHcAsb0+8Uwc5e4TCg8ZgFyYFwCHX51a9y7B+LHl2+P
GvMEkltUQuiODkVZWEY8QAFSNcBF93i4S3HIJ/haGv4oT1gbch6tJ+TS9tl6sK+lmZDzWPcd4/H4
rBvIJpqwxlkyvVKVjpqXdQqlxhGTl4yav1KmD83HhOR/XjkafWZkTK7nwPKYvwqZGdsPd2WBhc6V
MfGOdAAuMg+VR6Jyrr6TkT4aChdWGx7Ts6QVaGaxR5W0DWM6AcwSGNd2WHSmF5OzwxMhKCMgqSRV
fbDPgaKLmgb4m7hF1mDxOAwGsxbfefoUYo6mLYmkq/LGXDEuRHPy16mFTpnOM+ibevBPdAh+jkid
Sw+Wg6eaNGyi1abaVZFXLkRFRmiunWWO0worcUd1tndIEr3Y1dSf6Bm1ex5FV+66Yc7cZJg0IwKL
YS2h8dwS8ElV3/HS9jJBtvVhPD0Bm3o/CfEwawRjkbmuSSh7xvkDdVsnYTfa904Ensw5hMseiRFx
KBPsZ7PUk7WGS+iiTtRgE8eFZ/GTv8F/3c4dVClpqd/bAZgGzNcPGiEQt0Gh9CKDGHF63ReEErZ7
Tiyh5jl9MT6w+dbyxaHagNlZ5cphnNIOg0bSsuQ2Gt46Z8vNhYIXNiE+xfuZItTdIhm8C7P4c63/
MYYkpDT9V5of/5Sjp9ddyfzKth9Mzt2hhMH4TaIfzl+N7bOuCwunDYIeO5pNr5x0aizB1Qmt4M/F
WSbz2dpmezTTiLl5mu9HwxfD6sB849SXfhUqVMFHhrBk4QyFo+aS8wusjE6VrV5272Dexu3Wd7e4
JSDo762WhL2XqhyJhzaRIFEL3JZZ3AXNJsNmxBD7otkBuco8kDyxivUucc0z8ubPSwXpjisxoKEE
hg77LzX5bgb+9/+pEc3zINhEYwg2A+FjuUMhnnYU2f63PEd6hlGHIbkcsRreKPZ081cLSfpcMfAe
axKZtiUtzVr2mgtsqhA3HIltmwxh/KQwBZtqhOr0SyLH84FbmX349QzjVwJi3vVaxFa9yVG6D2wK
wRavIuRvyVninfeKezPHaUCz1d17SqchSOxDS0XU+3uqIt/1y2V0PhLudZc3zzw7ae+6AcODkOXV
JJGSKuLClI2kZigPeM8tsVIAQXPooqQnefTebVf2Nz0k7GnmizZbQr6aBZpAcwGos6zlRfT3aYnm
RdwbK5zNq1e78G087Ed9TcgDtwminDROoKORrt5Xsi+0grpAGdJBznkpNHqTWU5q9x5jS4uk2Msw
fcqrgYOof5k0HZOiiAcNRb5nlTAPKYXzQXfWiar03ESKem6LnWYPYjXD2WfHIZ7HtLbadonWup3+
9qqWM/i9+r/ww+7rCkfBMvoY1tpOE12wXbAJhSRxbgOry5xLzGw0oW2LEA63ioR7yj7Y6syXJFRd
Z+gXQ/JCWCJ7HpZSXALvjJClPsgE5oaCJ9XV2kym6CsFBNlgUrFLqlSPg4m7iIFHT3XRUydXOMB2
uV3BNHG6r+MlM0+HDweH2wvQCY3aDY4m9aMWg5m0ZAust1WJVzRHTtOFF39G4OgBIJ+gbCUmvqOx
IWiydaAn5Bzr/QynzjzcGvewA78/nPISXeTxUh//Oemjhz2eK5QYvBZtpC9JvIIGd8saRnsjo3o1
r7KDMWTwy1XWW0so+q5/2xvGmOZIv6uYPFn21wuEzPOjILMC/FR+P4EtvMCopQip7KY9GmI28XiR
EgiVf0vj8O/ghrKXc29YT/mRLUtIVLNfGL37CafEawEdSVBTSWjta2+/3s7lGEFzeTkbCeU47TQn
OqIAFbfp6UAMLqGInZVcHczg+HvDsaOjBCXef3nQpDopu7Mxsy0D6HJmhRcD0ZAUKO/d+cEEDRtJ
hTKyORNOH7yDJwWcGOZnfO/1IeCtcn1gEQz1TPNcjv9niAwWKRoTB9DfbSyAVenjsYUGc+yKwQsW
LDpP3X0MAI1aYHsVRdT0tzF7wK8S2Tb9UvYdCZFCxh7WDTp4xxphKCFIBfRBuSePn7peR3zcqh+P
idfYbOhQfzikzRE+qBUIi2xwFGEnUeJ1Ngo9tOQC02KTqTOf6PlMgAklufsVUiAwGI/y7c2oTaCS
mRvBZdbp3OztMsmILr6xLhRkVndxUxem0ZGRv9dOrfpCngOIdfTMa8L8mKrpsnyvrYjHBWZXSrQr
gjC8s5z+KlARWgtebBAw/0woJKV0OOF4RyJrCZHRJjUuR/dmc6mh8DC3oPV/HpPnILBjXO31kdOl
t8tQhge4eZ+NbBxlQHysUHjoR1mUEPcMObHpx+ZJ5eAYuTjZjRRLMZ4f00+FGjcqefoipGhejbok
uj1RFC3YyZE28XJTaSmzFtR2vH1/QBy5DE7Fh0zm3NqvlZKOx2HPwufSXAIhiNlQpSEa8OrFlBuT
4A4Hv18Qa0s6cMCY2OF09zEzqx10iL5GhXVl8DQsJNgZ5Y1aiwvDfjmVRLzIC3uSKSn3xkC78Vph
yJEN2CWC6aPKymn8MJ3H8T9YtJdqktol2fvKRdxR3I9CUO84ShVxDCwqPVwQfmWzywULE242FM6K
8OzxTtIqxvFepCxdDztVyC+DYG/JpoqFDU6X3DxU7mEwHLpFhk+xdgs/hHe2WRHUD8IJp7DSyMxy
ZgFY4ryQTCWuMLnpU58i9HSY9OGhHrtyQgTdgTj8Aj2rFI2Phfwgu/N8Kj2MTm4+fAmDAvj97SsM
mcjhYvo9pilEWjRAULXE+fPsmrF0vVw2SflXarupXVlc87T0tiKew9+GgKRcUeUeLgNIrWSTM0rh
duDPFax8igqH61uCeZ5iFOUCCl43q3RTvw9R8bNCMnoBIm4nmBiGe/fYlaJXmJzwttKrc0qhluAD
qZUTsQbaOAd+JzcUvhuXbNQmdHX5DDjpjzecrd2Yqbm7+lAemehPWS2sezquowrp4c2puCANtXEg
kBzXDSiPkgFvVDHiO54huowQQjZ7jTy0UGxsZIlcAA+FpSTXHcocBZcs+2ad5HFceX2wr4sDXsOg
DDtg4usaP1ewlZmCoEt7c6Q0ZSPLDdQiBMC3+J31vC6BNNHCQzwahQX1nXlAbedDAxhhUkr3hnlG
7o1G+xr5y7HEPYh4OHPf+7lC/vypVplkxObIOGfCIHfEOQNOkka6DEnXx12lf/xiEy0aplG2Ab8T
G6fafsw9eBtPCwmA0KR8rT1eL69Wv3ixjYlx1G5qR4KEv3Ps98xT8YmxXMI0AyojID2RMtDt4qvr
FKlLP0wlNTFsH/PPEKla+ZWHA8RJMqIxtoPq59mmilW5qNXwnbbviW8vIApuhZLlBJkGWngWV9Xk
3eYaEGQHMZBfXHMijzuOAU59GEE8O/3l0BajdgMGsD2HmQObY4kcXIW/IoXs63Dm8V2wslzzqhT9
IU748Fm8SuibjqRNadirlP4LZaOeScYQfrtf2ZtHiLwZCESyo/GmEuZOzLQCbLy6C0de8bp+c1kp
E9VNcIsV+7j6bbY7fsmw189RQtv52zQdRvjRjzsZHgX1Q46mXw1Oa7Ex9c+ktCQQW9iHlMwSOOsm
4sRxXJ979k7nphKfzLM4jTmoRqSUVtQRbQFOg79R7dTGuOZMa7+Kmgjv9b254d1xJrziVrBA1Ko+
XrV1fnNJNojwuv7LteY6RhGh96BujrCLYFRYxmYH2kv6tM9gOkX9E+RNG/cTtOAgV+jup9p30qBN
7AAvmVYbNAFEAdSSjjlcs5Spr0FmVR0T7VJkuN9H1kHwGmdbvbhiLFUCX4HtnMssub1+WLHk4jbp
ovIzOR/LHz1J4Wp/2dflIzkTnGD+9dlvukGpdf+LcRR7dRg/N+duOI7/oYM8sRORuTmiYZOF3Zi5
IUn098pn7WD9g3KkqNHlyOpnCiaOlDA1ZeNfF27YPPaZ6olteE0v49Enf17tvdtd82ZhWSFeys8e
Z9H6renhqQZjKcdFeba9xO+87ZpIokrTf0x1lYQ89a3nEyDs+gOnExW/OxTt0Eu8t0LGPj7Bs8P7
X0bowD8IfBhoetc2lVh9Y7S4tQDwNk2cN2lIQuFM6u+R3QUKmx/D80VX+cH7B5ZsH8qmD1wzGgBy
zWFcwvzHZwpGwKETS8EitUjw+VQGERZ/K5bQO8DDftrmRLKxDVIh25sbcg6eepM/i634nrWf111w
nTmCgIuudEiImydYFRJPywhDn5ygulpsMjA5T9suOkBocP2qG+2mUfJiUgPF1xcZcpgP05mjaPvo
Wg5SfR062WsAYlhwt8elu6sY4amUeMq160sipj/YEi6nEGmDXCpyyPR7oXQQLQMI0vGZv1ky2aQk
WcaoLiVDEMBfeV/JRrjU/Is91UM2SUo7Lv/U5FiQLp+9ICT4KZDyNSNYWOAjHz+t5eZh0WyZs9Jz
zSVvHM6b6AmC7mclN3nZRb9OGBK7GEeJ+LlpWYztUsslYMMmscF3dTQ6FUpB4a4eOLK/9cPZgaM2
PRSBJkeO5uYwvgF3UPgJEB7d8y8H7wBzVgdcqCohMkGmGiMEnwy0wpYzOAMJUu8pRo7gSMJvvW2T
hI20dgphg4D588UP0e1HDANi9911nTinn2nl4Lpk/BLGGnppwwAs5IME2ToTG6EPNhx9ida7kcEF
/abUjrzm0fjCZud/Csl5AUtODlbHp1UwXNT1Z9isfdWEwb1GWdNmco1l+I/aJmqPP3OchS0w6+js
+g7dzbJnZeEbcmgX7/Os7XWxb9rjdTf+TQC3iPupCQz3YfPDOg3ibG6QYqncRtKaHRf78C+knMdk
sEEFAj68wA1VlDrtZo/Xaqqxpa9w1bFRxIm1n5ino1EkbHQoMV2Wvv3li7GO2KgJhPdPaZh1i55n
6uAR2rBfBvOW9tA/y8ytYtb4Xjvvb2zqZWQZfOKRZzInrpb/AIp4Qkb7xdbZh9sL1/GbP2gHeeIA
uxWuW3M2Hy1GTqUwJm9YnipdHvlWN1yrgJC4pgnY3KyBpnIRfT8ECtgIZLY1Q5fBaj4A8iyCS+LO
WgLYuuVMQwAr5EyzN8jAJB2FJsQn1GSJls/vLyq5s1n+Xp/GDFiC/Jsr5zNHUWtAdZAV5taW38sS
lP1bq8lNq/a8XuAxbjHdvFoDi+6tBOOuWQTqSGvs81r9q68UZI64LZcxN1mqOwLHs8Y3aQx7Qpnc
bEBpXj6+kwjZQgCxnd92ulzU6sYLq7BL2HiG95ZFkoYoYJC8yrThKXW+B154ZHukD67ngdaXf1j2
hk2e9kZvU31Rak4SHgn7WDsalr3A3MLmphDf8k7ek5qS4v8ODn1c0McM2/hUpuCNJQI7c6Fa+O9F
m8qZLJsBkvA2fihEEjZgihiyCWQQVbH/EpyEiDJJQI60atdXdwJR+HZeoQ0XA1CkQQ/qLodIoMVQ
5gGGfrclr+qTnfZZptYzlH/5MpkEsl3q7of6J0adwO4k/mOoQIb0CZlDix9DBsSeBRPMWiKhCWek
GBT3a+2s5khffnx7vxl3EGcH1dg5w2jdqWB63Hvo8a/TAXNigh6izE9n74CDY87VoMFTtdEtYr1Q
7CNMrOfV+IeRgh5mFJJmYEfmjoodsfGyWjQ0Ipom2l1nQzCW4t0JUgGulMTHnKo4t9T24y4Fntqq
9LuIw27Ikrlk3IQm9dJXrRSJsZrvcocDuehyGM2ZYhYtnn/8X4lXvZAvy+SGCCrCAeFyceQWttjf
nyHnao1qptx8eD3ZhFEPP3nEGLtY/oSGJHiRAkqjXMNXlaMpejubd7/YLVSSydvwDap6VPAKj5HM
324lyyhF5yI536D3I5xnn4asm4+JJFc73dEPIvFIfSF4M099m5pNW77rrU+AeCDRbEH1SC41Ihbl
a/bXJRA5fOZ3SjhYWTJgLAg2eMXJmY9VQySb7/YVEp90u1OLAmeru+LCAGJ+V6k3yB9mvzbJWa8W
IQYDi+aLim1zYZ1eYii4qhEKHDxvi1XPPgzWaixvgI2Dr5zUVk6U2srVvPn4HoiMaQ0V04Ril6CX
O8wCz1Sr9oB8NIycQCzB9qMwgJoMDfpzOdFo0g50B5wJwcyP+/VRa/Nd0QRbqVPGJIn4UggQXrUd
U+MKhSRCRTqKUyAmx4MRl3n3PWcnormJBl47LO/mZJ/BaM3F2J7FvGZFGZ7IOsFDvJPl1EJj4rp4
yIHoaCrjo/sp/OOvLQTNAvJUqjiKx58yuKL4AndwZdehrio7Airxlka+22ppgKO2W98EbXVhlFuY
7lLY6XdNa5A+L8+4cDEhEsadlbqXihQ+GBz528mVEKYYmUG6Ma1tnHc3HYsi8BK+MnErxq4s2mdX
1LIaiTGlsXR8ORTR9HaVF7LAqyV+bcoxEjxR5+iow6MHxy9Mtd3PtxCNqPspXa2BdkSKstPkkxwX
zqJO/8hBTQU3K0tXouSuf8djtn6m1f/1YQnulKFM99/+J2UT9mLHiS22RreUJw9Zp5mIPNDk7Yzh
cb0txsJCyQB5qpqmmnL/WMpRyRmmvlaG8CWCG8aPwSGXvJQO21X4+xnpRjjmWERbPOiBeQdqwR8a
wcX1RtuA6s9BsVPM1fWzTb2LCvelWH23Qdtn617tjBz1p6ANRApmTPZzg7fy7wbDCNrcjr1FIuyO
wFOZNPhojkJK+UmsvXgDTiXM1VYIOSYp+XcM/hv2Z7JAGjADMWxaDrfepYBLxQKXe9UWSHOcyfub
ykQ5UcJuD4r9Xt4hkp0nGOumOJcBpwNvj+Dx+/ohONpNZTs5SBoeRbdq60nJTNnryR/QhOnv1mSh
dHJYjOz6rW9+Ju/Hm0bMJXNVVqR99ZegfYVZ3LJyR+L/yjUmSUkOmAm2keMTmQg4vpeJVOhuA6c3
pj1VUFyLzCpZ9T7+70YevRjloXNA4ZZHYn6FYaGNZnztUQCMG2ByUgH4yxbycaK7ScfOd61GoR9a
NFZhtndQfbRIfGbgPh97hDYgnNMw0BRo6BIkE3MbPhYHfyyzKE7x+2g5nfcQy09F69HrEot1oYzz
Z2OjfFkOsL3OHFOLd7HGWfJWu0EJKVgqEi9sq9qpKA0+3FrnZF5kQUyik/y/C9ACxm0q1swpgbTE
M8sDvMYfsI1KTFZrT+O+8spRxeRb9D2iVCAxvZYNK0QSHAAFfoZoFs4BaHeeyHWc6RMV2d22Sqph
u0fIijRbfjIuRBgLdjqX9sFWduFs+FyhH2hdzfvhqDGX6/8qk4yhXIriY/Pz+Qovw0JU7A7sf/T4
top0ZWAxqPM/NQK1/3oURe8VdQJRRUD7QtMcUjQGKC1b4St8QSyHK+UO0EqDf7Kh7bGTtdcLWQKy
acxmkHngNR1C4gjG/S20/G7gCTyk1jxfcj66kvj2PrBKJ4ipZHau6MzhBxOOuxYjtizZrnPulOIK
epWlAmqhvlN7h0m3WZ31XgMdxchcPuVRheyWMlkx/O9Utrzx0zCE+S1lxemOvu4IDiQCaShfaXJs
ocu7kj3/H2wNzP2ShYQDqspMaWUs9D6p3IQjuSaPL2Pb6NydR6N3f6G6dc6q8upE4pLqwuvD0zYs
dUQbkn5IYNDY0HOrCWvVUXv/c++TDP1U7RWWoUkPFLnH2A/KJ1bfOen2u02+qDohZu8D5iyKucdC
L2ctaPvsTpq2RixDocMnhkUVrQEv704kHeGx+oBAtbVUBBArC0/hisi8684uxEJ3tRDJzXrFWhb8
W/PQlYFUdg4cwGLQMrBH46prTREx7xJIqsThbMyvffRZOugw+lDVN/DOMOGKxpf/YeDyFFxKlc7x
RYJhcTzJh2480IUlU9N81vMKH9PsR2yUCbOC0KB2KQ8p2NzpxpVCgFoQGU8BSXQ2nb0qRRhZb6Mv
RQlIQ+qM84VpaYkpC56LDicfXTGob5TvvKY97vO9zPAYpNilr8V+HEV/pMfmQ8D1ra1OIeH0aCXl
gst9zQblFTajFe5oZjoRO+yBHNDIV0rAIPBMj4aRkCzLPJKbUAmYt3VvoMQ4jk1tfndpUMV5MmP3
XocZDoKVTv++2yk8Ivo5urCxZDJ7FnsvXnShwcFwHmcyY4QtC7rXgPIBt5AdJTllsytI2IFB1vqC
dM4ORzsRQbWK5R+9QM2FHcwExxlZqXm5PNpPCpYL5ueon3x8rbF3GpVYLB/nifX1setfdyID3KVl
WCk4Y8yOYedcg0Yjen7xZozom6AdflVcvkTRWO5207q/BNkp//dNDw4KZ7eOruBTz2vGnFmvM48T
6f7sDPusAHfeB+jLD6ShZwAsBNEcRJNhkMT3OUyiXIn/R++BC6N6PcGYJLP89+1YTilFY/t7x6m/
9c+2vFUS0MEVXH9SwJPevpoD0UEO3nZDB3K0LMyjM4UWrbNECdeIY/0ezYghQwCnreJltdHdlk0u
etsv8Jl/TXkhjJkat6nKDOdlPtjfIoDe5rfPM0jzau685fupkj4AH3zhRELSkw8Y4ZTxC2XF2f4E
aIy3Kdg5P/AEK6LDi50uv42SO5zKC+L59lA8qNsgI7jjEN1oqZHmke5n69oXXRDTvIJoU30YFDUE
eWm/x4yhwjXqbuuXtzz1pEzqVYlul6WR+kVs5y12Ss/tEByf9if/9J39/6DN8tszAOKX0SDKPIUF
Ql0WMbJBwyiqMmy6DOmK1fXXvOstfeaLFalxWrdHlBwB5cFmqqFy+NM7B/t197x+CEHdJlgHAV4d
KGnSFCRE4oSjpEmWDNvzaoMEdiagwCkbDY9zlgZE3D9JMuDNwgFSEF+TZrXXTw3QrhavzWRIV2s5
4Pr0doYelA0Av1UzmqdSqOgP0ZBvkP18owedZcykU8qjOxx4E0YfATMAIbNKI/aCbdIFfKJFI/sU
h/5Tkzi8fhlaLivme2Yc/zIkw09luhc6bRyTEQpRjflfYCZItUu6WGJqCs7FdPWyVS9zMcemzpN3
xvkVoxAq3y3Ipv/NO9ZZVc5dAxSld2KZJSL1HYMSmz8pz80tRgwdh8b2pLcyOO1KmBVXqvWAGd15
4gnFS6rYo876k0stmJpJoBkQ3fc7kIEEik3jtyEnezR3MweRXXO0gcXJ72EVI24g6ICJsxyZZp3k
tkxmmy/0VVVu0YG+ZhKCobefKqikJc8XcsdBTpqcQEs+N4V4hLfCA4DHUq6kMe62XUbe3lGTpxIh
BRSdvNAozJs6tlRm0BrHZu3c9i0+CMqV567OBAf3YHrQihw/NY/HsydQu3TxKPQAPjSDUtd+rANd
riCj33qcbaFrQl+nOH4KcUQsUqZR/avcpOJla6kpQCh8xKE9oYAPGzOtJ2Kr/iLpfi6ZZJiV5k0v
eWH7Jzp2a6+e8Ty7jT3FrCLymmbfcX5RfAvMR2ANp3f//Gv0CnpLbSOlf3fIh1BRPNdJ1f47A/Fi
2srE0vDagHYVo8xNt61g6Y6RAaudEb3UEBKWUgQDxmHX4T0JchlIXxnheb+InF1IAhr5t+m6bcAt
Z1I1Ijbx5+ttPPofy3q7zvfvhblAIZT+cCBi8+bbbZ9KQ8LisXzL4asxk1kGi7M7nqxY287huQ7r
Pxw78Jr+RY97OiNIQM7JgcW+NpriY2yADA3NKLDSGmo3WBg8XT4cxmrAK0Q70INkRfLI75ZgY+oD
XI46+/yucvErG49GMJHaihi08Bu3Opt7B2SLVpfcAn0UBil8MgjN4RgXXfYQLvaySyYFoiO/0lX0
UL2Zm6qV2gUkZtYHqlIiGVKzViIYreFtW0YdKpxZM5IbsJeGIZ1jkMsZn83TZXw+7rFf4b9AfMYw
XJw1B12iuLPy68pgpecyKHuPUjNNyOO6I4oUu5koR7TYThwF+XREXt+9cvK3xq3uiyAMepxGdIa0
oJQ/JV095txMBfeLulq63JfMFVC0p3y4g2kd9cLTckG6uN3wVqN8mHkQtiuOSnZbo+7FberZK0Ui
EpG10SsGFzh6oN34v7LJdaYobX/5R/+lET1BZf1iovT9NHCPe+vW/vuzD929ctMtR7B6eDGDfT64
Qz4UtdLMP6T+znWSjhDhA4ptcyGa4vKrVs7I85A4GCZAplCPP+wglnaERSCXdeLWey67tJ90CMJJ
lbM6UBcSvZoFKnyjlHeBETl42hXO3ptBjoPb4I3xhGFfoMrwnGq+yeo1AzBdCJzrRPgKuMeR66I9
Evn/V03j1sWDT1lwnOL2xV1Q5kHrkTO+2cfqRxonEcyufAaHUK+5/F39cwS3KjV6FeB4HhuIGTJQ
wTrQakeNXTyngvBUZZ+ykeh+oH4mDNKT6C1czlUwCg9PrCORH/zEt0w32IJByzOzoYdETuAV8fIL
3PqjNRvtxk+j25yJ9rkptPpXL5O6e+IrxDoKKqmMo23DO35tauF0eHPaQjiP52J1d/0jCktp/pCH
YSp155jH5ahJUu0vxJAKzcxibgtMUSauAGzvFetSPUS8DQMhoGx7aQqQdof0GAshf1uta0uJuIgw
EgoksmArknpvTHOnLStPYw5bMGPEEkN+IGoFGmVb9cenmvx23N9cjqTWQj07r/OpmMLPs86dGmmU
Z4yA55c3kQ2WSwwhT1oJ1RbG151UZFeTti7puFZQA5Mj7jfbZQmYR9abvTIAagqumVOyTQeEdeAa
P6bqKtiVNq7X/g+D2CMSuMlaKMrN9bQzNCe8ffcwBL/VnsbcwOZY7oGq1Bw2AyN2f3+80u2nfnwc
FtSLlqsvM2sYbu9Hu+XLZlPnPdyVWQcLNIo3AqvEfHl3XvTFsM+9M0daLc+t688Tn8VnI4Xlk5Ix
D00i0N9rENAysPKeMMEEEw1Xbi70Y42IYPpIuutiFOfRw4TSBVY+kLq4G1bOVdGBSK8Q3G8zLeR2
qkcD/8vl+PKW6e02H1OJc+dkPG79tyK+VIk+fsWV4tiYFfct+kk1GCuEkvVl55TXAtItLuoHFatC
+Q5s2qlXP5YPnRHNqvXMYexpoz+dFNCUF/jUYvUUD4p4XTWm6JFNtWBlxm7TUdhMn552U8ldt7oi
DzHlMp/LpfJ5cDwvl5sKUB+yks0o/0wWuk1hURX/hMN6XJ/rnwcm7QEBqQ9HTemGMGJ94LM/fH/I
44xLswOHsmGpL+K+aD3GOcHTCRCluo0w43z54PzCWskUAnp5hkn+0LALKkaLu7YNuU7R3VgOxicS
gWuX3iSICuUfqu2FIL0vDHAtvpS34LfsR4m0dpCw/7TUxFxl2X7CB0slMCPB1aa8Bp34GCk2bd00
LT0C1FPGV3Eh/gGkXrrM7wgtcNpsarOMPjIjBYdUk0EfKT+xb58FmmRFsLTSTaKytqXZ3Oe3CNeq
sd6iD31DjqUNCNXf55TAi624st8tp4q6ZMaLLcHVpTfibvrFr0nqrZvcvRWxdtQmCPvKvOoxaJAD
hhRIKhwoqWRlso35nyq5vwwc2i9FFsFEfuW90qTz7c73NBc68WjoX5CMl4nFoVJNB8uJBysR1HSz
fp6faRGMlUSOOSHy6eDJDPjDZtygXBdvw5k6/Pyxtu6Nz/JQDVWkj0axV8c6xj3DoFEv2WgrNKmc
w8LirtHcS6ytjo47MzTu6SOEQy0PR89v1TQDcP3StAC7r7aeDB9pbRXjMQXi5qTNqB+VFofZ7iAl
DP/4kmgki2/+57dxcA3wD2kpmhosWMMxSkAWJDnTNdXSdAwDpbe1deOc66WdLQYBVBGAJOmaq6rf
+kLsZJJNnIS60grk8nLXffJfUeqAVb6j9Ijq1iyw63mDfAKBFCNiIzWC3T31hKK6zru45I34UyOC
zjEmLA5Mrog1re6gCyiAzk9p+2cXXJtE1mJzd9D09eHGQc7U1eXCLYFd3uOHLyUZ8TkGkHbkg+E2
EJYzUAsB3Hsu8oHmuDDuLvT/JIUGtM2+nZDUZB64Mh0fGfIVNzpPlZHo212YlHsDhPUU8jSBjgwa
ywdX9Fj+CFG+uELQvRYcbyZl8SAJg4g7di3kwTokexqiSkg+0tRuS2lnWkgz0hKm8DYDzmdYXh/S
+UvOvqLFirfY2k+OJ+wA+hu1rLKCYBAkFzbenaAwG62002Vwv1Ce1tBaWEfrHZqghR6OEH875eNh
7Ifx9xNwYxLOYKHSXgLLHsAaTxZ7X1gMDvKHiA/eUZs/TpLIh/MD7fi6zUj+YY2Sp0qhmaC/BWtL
5IVr/RekRTerZJQqy2c+hWsJIpOoqFsAHBncdgZ76AhM8MJmeLFHZuTRkKBzrGPJ//JL+vZvfY68
lK66Ma6At50TQ12Vjdj7oPhM1shl4386Tuv5pn23FqphUGvZr/w/ZBi9mabkVIBIYd55qZN09WOO
2iAORE/v6uGmGui4tZuOTh4oMXJ9lSUHlsPYcrX8QoNrbj0TBlq175hV9T5SmESsogYuEzvp+hwV
NvqcN9OsOzfS+vqz8eJwh87JgFS/nUn1sv/CM+OghjR8FTuhbEHg84J+fKRzGUjePnBpp4Fp4O6O
A1218+aS+9MfkMYyN66FeB8yKrzyhgiBDpWKfxbIUpAPDAIDVDAN4IYd5sdyG2tjkCpzwL6CQrWc
4SwcThw5TbTKDgo6RkkdW5mIvFZ81gO5CpOAVUbCxefforfC72fidWjtJATfXFKLg6e7ArLgexf2
5X1GJarJqMaLiLb69mCG8j+HeS3g+tCFUfU6vemB1CIJ0ttqTHHKOPllcS+u0r2LNHkCBkngsA0v
HCZhXCruN8diru5v0gYFTVH4pueor4P9v652QZUh8luh1ct4aVIEBV8TOA9+alKmNlrRumhdygLN
pKm1oy7nmLyZ3dYbwvS9yxVabcqdw3mTm0oy/cjh4L886Cgwhhys3WY+zrK8muGX/uK638ibJXd4
ZErTjbF0cYvB7anYzmRvanrgGU9COlwchE5BDmzf+5y7KPKHmGiDVTP46KWvPBwmAEac+V9OnC0/
zq1NS0vwzD4A9KWAXEygH6M/Dfdq322w5iva6MfwCvxHXZrvSx70BCgq6QQZ9r1WHLtOWBkxX4U0
PLH2wjMy+qAOzTaYAkO1yaviykPc6rZPcHylNVrCpIs39GJgAH4QLPvRhIjekU1iiQvZHCdc3Jur
yGRDNWIB/ZwgJE60XL7POx27GT/xIMEAspSqVUJKO/adUs5QIQBZmMKU1BHBHxAOHoTtd73wnprJ
59bdbdh4/ghPX4b6SodgxUQmgdRVzv/nHwQtAHSROmE8dFm5edsNeKISvCYa8sdPf/V+YapczoQX
1Y+E91u154AUNBG7AGaPySMYIId70uiAYVmdKvuUZytb/l4gbEVuKOfuLCkpID6HaRIJj2cnoO2l
NYHWSh6P1hZN+w/2d7yAAPTC79bOXhmrIH85r0+efD4ABcnDTz5p81jJqw/NASV3Syldh2Z3ST78
QRLWSw6RcpE/qP1wf9zRbl+HoruiZcYO2qPWK3w48/rwGherH3kUutpslPggafnRmNRINmbt84fZ
PVvEJniB8rcEpfZoc2mvBemsTpj4upwvtEEGTA11ZhWEH/mXiO4QhFU+VEnURhAHc77sEeCptQh8
9lBEzlYjFtM4Jr8UmFhCX7I3HPPf3ihWf6yo8bBA0uDbrcv9j1CJRqiTpiS9H4NtMMUWuDFM37zG
9+XXHsANIjyWzR4VzUytbET5rQ6RB2nBWH451wJ6EAuQ+gJHtQW0uKE8TaUoAl3JvC6SddqHMRd8
zTm3yz37TKGIehhlMypQX6oW3QwvEy0sEgsAP2jim6Ihbr2Qwn0bon37rH+em/1BqC0ZFazDWUDW
AYMaJSFR+Y0E1mfX5C93JKswf133HtRMgDQNkyJrt4CAXPyA21CcxGXEAtn3GSsaehbWcJr6rup1
GXZuCU3LfIdcb36L4CsQm5azT4GKsFB1AD0uE6H26YxRnr9/lSoCi3SJEbY4mN/gEBoKp/jWMNdE
+iVs89vFyLxuLz8Ok7MxOyGZN63rr+YE0QR4+a5iCd1s4Vx89bC2OOt+ACAEDALIn4SdpsU+aF/2
0ul0CPwWNINGlmjsCNQ1mDix+R476vRqU7gcf8gDA288VbkjvCpaNHri3O/G9xnDaw1t7N7db36C
7oTocRoHIlija3pYMK+/xhFqENM39agbbm0+s8jh6WmRkepl7X24KSpR2pUGzwJP3RLr3a5iBGNl
XGwj4rF0SAiIyTiyfTrvLZGaAOEpYH5fBnuJlmxJ4xOYTc0adk8TCP+4a6E3gxZye5N7axR5X67T
jA0Js344sS+4aEJxGCbw83oC2yQOW5SiYxScks9vzxTVieFCn0sireP9ttD6RjLsdWirFipiMDHi
kXn5GsfZkV6+tTf99dHqs8Mc+YDhEXJuJPWv76YIEKnNghY4ieAaJzQDdvjQsp+PNtf0JqFYjhp1
Dgq12x2Gs8SXQ+yiLUcgT4U+Q24zxo/fMwtWWqf3/5AnUTtnU0n7YciCVYQAxd1fz8ZdzxZeJZwX
ARMX3kYI2zR8aJVotuvWSu5R2Wts1+AC9iBspdIQYF0jHEwI1IakpuJTMSyMR1b0AcUDQ1T2xMXn
3ZjsBo8gwSh8CsStPdQWbH6nwMOpafujw+wPTDvpZ/JFJBxdUJf+0f25brSxpbs6iZIBrqcfJB66
lHTz9vHMaR9uGYrF2IubfA/ZgbA9/JmytfxacO+dG6yt5GAsIzt2rgY/zFh+bonK9Gb+YwrdQYbW
oOxdXrhfW6E0oiZPoImaTYUlb3lvDxUWWZYHMT59daS5CBz6FY00YO5s+A1wFNuLOXwERZLz/XKZ
RvkSkZlSja2UkAM95h7vAKM9NoEr6H8TV8cDAmJ8M/OAfm3ISv62nHIKT5fX3gv8S7sYcNLySg2g
jjT3P1NHAVeME7HQ+PXjFDbEfZjvR7c0HzN2OU5ECV9rFTebXjuTj1WL+MitzMgAGyDzHQkmpP5G
7lj3yxujCvv8SNyoclBcAeW244qxYXx66z7rTh5T6yp7no1kSaynYmwuRluqUNFGeCCZrId3/+Ty
2zAk/MH2ZKgtyEvu1Okle8NGmmM3gTQTp3bdd1S8c20JMd88OFK/d8dCuYgdOg1zWHZt/USh31xz
JvpHH4xPM9UIckOlG9ZMmw8ixiJ5XFBuDNwi8uZZxCqmvOfvQeyV56hUZXv4R+cxIso5WM809nT3
Xw7pf7OSlDNHnaLxafygWZocFul00ryWh/zrsWYA+qTb9D3ctrjuJo5LdGaB234LZktZ8fq4T48b
EeqRaYMYfApG68Ezr9W/1fdddG/6JQ/fm/WIKYyJFF/53dNluLvOshZUu4+y9ts//TrOHD9p0iLv
rwwSJFpJ1SB+MlbpQBV3ZWHFGWo3rBQbfNrZ+lxdl7Q//KJuMoa9Sm7ySgq2/B6WBDdgTFKVjXpO
surKFmN8LkZ8kXPRQCj9SAK4b9A5nx4CAunhiahyyyZN9D30bC1AVAH2EmLb3ExntV1hMfo9e8Lz
9tMz+xjuy+UeD1xTXqT4/pCsPwCKUtomDR7s710vPwhjxQCSEtQZn4gun14H7FwjZHyCkPtndRm9
1givv+1j6fmEM46IAbllxiN0SqUl3Cnbp8YHj34gBHVTm4cHV3EljwhhvufMBZ1fMRiHVCV+uGXB
mH+ZV0wK8VD1pvga/mhpGPDxnV9prCyKtO8kQMZSLz+dHCVK97xZQp+dMYpa2+0dyyEgZQInl3kk
WaaZPSKwPOR6vNz+fimAqnOZQdvH67Oc/uh1hK6wwNP/oUoimm7J0Tt+DXkiHhu6nw1XAYeWtGTz
FUc/EC88u3iTdxmBV9Xbl//p2QuKIJ3zD7/u/V/Vyb/bkmdjhcWFqBZ5HxQ4gSVCY+wXTuDVvgOZ
PiWx82OTxPIdeau6SYlxLKGe7JJEZpz4Y+cCLvkVHEE2H0AIojlLvLJ+hsjMUTdmhIgsOGi/LiRL
17TFhls7HoGp0Y778/wOxxH+szsxvZoKUKhAe9rgGrWVZ97/SdOpBZ0Bw88BidfZkGDbybu93Odu
0Yb9UV2kKzobk4QoAT3FTCUhAK8WfdV5//CVgUOGqaBOUfFUzp1T9Lb6VeN2gIWO1IcCGAgyVmRe
pWW1Av94ZSqW500CVb2Kkfc4FLwVoRODw2th3lfvdT32AdVHZBFBVoyUu4oD/aYxewyyFbnDwPUm
GWmS2nL/cUWWrEwdcvPhriFsY/voaJQeFduLxbPa/m6dqobPejM+L62tOGmqGO7QosA6Bps+434e
6GJ9x5vV5yJElRhBzbFkSCIV20UeJBK75wiOzpurHH2SxqpW3Nc03pTijCckMTDJvhdN/EjebCBV
vacKm5j73xhZVfHBoskXSO/QCaNp4CoqknOAyZOkpBcGrLbGiaaVGdxmixuCtjVOXVyeVyaKicKk
MvWa7aVLz/NtWKfPPqLpUBFsLKYumJmbTu0qTSkEhiOCFXVZkdKth+G+L8IBMm6pl3HQf6Ahabi0
wUj5zOuyKFQgDYQdF3J1Gqptays0PFazsCn4jVq/c1xCs9zmJrHRQD0mZaONXLEV19cYlkDqZjgI
ZhiKRAZ2BAMLd2ibUvV1qEOoivQUG+pI25qb2jvnKSO42F5AlDJP7zJ/wqDnC/aiBm8aovGJV9Ri
3UYkNUUWNBX6nK/piBRF2UrlTID7RleRTw6OWz1rSA95BWA9KdEjPiNPsW20K6xdTeVVPlbK86fR
a35Gc+jgWfdmsf+PvGCQ263FcPARd2wL3yXYEA7IHv1h1KySdatNQtNvCbKHAAU4vopsGg8ArN7s
SyGpM+Qzx58fyVGqqbPfuB/XD/wxuSwNbk95A13Fw6RBDf1KFT5IlKvnCWdV68tu7U4u7+B6e6Aw
pJ2jsqYICFSQ2Pymjd4bF/dMHIV2cyy7FesIbzERbnO0dm/Wl4TexPnX54Gdk40r98SiQmHWgwQw
bgbK5zEvGLRr1CrwBed9Hg+3hKfYOKpnp+U70vBrVf6NY2sPD9syDj0/aziIzU8M1rZZ5JzhcKUP
gAtztUgM7Jldxf0O+vp7nJ+su3HQe48C2EAR2MwpZ72ICDOYSjbTc2Gp+ahl1EC1LsFpywzwV9BC
5WkXL7H+UCLLgVuLnmfAUlg6U9jB4MKMri3h6LwW52qlWL3B6DCg/oxpZf2SWalAKgIFC3IpU9x0
T1vlKZjXyY9F31dh3hU9gcGrMrZY/gLDtTlTHK+gjRNsKfnPnl74UdQkWBfIIxlinwAw66smx3FO
ZSVKCcOLmeYlUI130DWLZdfGvvJibjtwMMeHJ7kAiQpX6lE21WvZX7TAZKxuVPsqeLzRGjZujide
gwkbq/6UEHnH9RcUJCZcFJHA2jVUmfSS7nT6qV6M4lj7we5iEY7YuaN5vXY6uDQApSj6vNuyYKIe
vfLcp5qxRIhzQy7NqQIDdaUTiqm+qw42dmcTC/Aesi197DVjEyZQhhJgsWR+9JhUAXEcwNOQ2sch
dF1gxQT900WuHjnlmK/RGRmv6Hjg8XsjhpFMMcXLAq/dCERTFapyw/mS7bQTyovJ4D6wi1gNiAJ8
B0fioENgyppIJd5bBoUK/oGNkpVcTK9BUTZ69/Gk6TNAd0ox+tbeZWSboWmL9Ldz4K4t23e25Zp5
sqPXeZASX3kh+Si1ZnTVCXkUATWkEiAw+31xFdDm8wQW3oT4L26eUOTk+7jwji2lMAfrw4HY0+7K
nODihgliFxVhogCWb7pa/Er3JlqDRgdtbsDC0HwPPZ1JVTfiGZyb7LHauC1k3typU+gk+sqpBZSs
NACNgBmvSkkddq4JEhg9yimaLlyl2WYg5hLTfl0wWr8H9MEf8m+qe2VR1WyplBNVNhPjFxSe+VT3
iIF94C5CF4FoV4Rf9DbNnBn6at++UH0++0Gm+WfwPkK8F3DFVM9PrdqXKMpF665nrR688NLfPyNp
DQEICe1PxX+PxZBwCg9buqy4N8wJmG1FPqh5uuO6ngJim0U/oawYIehuTSvgqhmWrg8rbuTo3tvO
r4YCUI5CSSXC7wEGyjFFgx+lwYykzR0zyXQtJ9oWeyqeGy8hLSxnA7+qs7gLr7YmuqRRiHZl2OgY
pCHr2XxsJk+L68pvD+0zNE+XzJPRXH75sl9WdhF6qsvjs3LnRm6DrVlCmCdGcnSczrPh4BYRdQp0
Eka79tyTh3dwhjgEd1ydlWGoWiW2Utc2XFQTlcNb8zlAoSoqoNrXaTjX4ytbfbBVpZH11dXR4joB
agLyqRNb5rvTVC3tIlFXEL9Ou9a60CY2Psr4sLC9Au4b4RfKVX7zoWgF96OQuuuwMDZ7ZZD4NSa5
6BM+6cgILWzSLDrEDuObWZZVX5C82Q0NFwLOh1Vz72NiIlt7mhz7o8Hcc2RC4INbSZ/tGGSQV7HJ
ONOSRGa4OOXsnTmt7HcZ4opDPkLEEXJJ1ZavYbGO6nUK5Nv9TF7mmYxh8zgQCYs9CVKnwvLas1+8
TwAv/0+hYhSbytdIb6DmjeqzlG8JlO8ltFsm0tJ9ZyhtfFCIPQqIVuWWiyrFHF0WPY/PXSo8wQGK
EOI+dZhLFKGbJR0L9iTnf5OHzwU+SFdrAWBNJvUwVTaoq9fVeWhTGdNaSuxGjzoDvNbFr5jemLtN
G9r7yvZI0EcREkiCC+tVpkccUfansua8kQ0W7VcbKD2T52FLkof5ELoQQCwc8KcBe7OjVkDSqwIy
wSDxo2I6ockarUP8Ntj5NWXtMCqWOpo37f/vsML3RkmixwAw+vMPPCCxBDYogDOzJclwyc8e1y6T
lXkdirvFh8VTaNcul+9bAxc6EO20AKmcLVJMjC6lLT5cSUpbs8TVk7Gjpbrlb/dOqN9gCaMABS7R
B1TTuHWVrX+A6tsrLZTNbM+TCWbMkyUtD5hPA/w7aEvhreFOOz9yqQDRwb/lITJ64CTD8+lnCzQv
Yv5pt28AUP0Dvrec6AsbQSVwSfKeTPTYj10oqFpbRXe5X+Q66eEXkiZpd6kdU7yFmM+kzpq0dVuT
r2nXkhyKI88wMMMO1X8YCXoXMpR8ZLSOy8uXBbk7s8ssxu5s80eIrbt85ebDuY1pa75DC1pkp6QQ
KeY5eElvCyDZPGUQahCKNnjHKWYZDzgw1n/lv1izCcHZtPK+AaAUQVnajxmVL/N0IcUUn7//tHTw
tMofv9H9VTA8zE6XiEUb9bRyPnCfPijEuUs3MJbLLViPHYFJdEPCWnfh9Ktf9cVX7nAxg0KZnTvN
r+SS0ecB389utqbsHNwoW01IVASXIciFYxFn+zktyKE/TF+tW2L4bYXfMKv0VUVHXOvCtvcsJwrV
7HrXVKNbdc8SYPwm1zzOvuLUpsyrDsJxnhqHso+O6wOdVfogIVtluG50kbxoc9csgpnN8a/Ekw/B
3hhzFdgNJnHpWm9NgTTb7TzogNCjJvJgc1CS3BqR/YoxZ9LypEBazIiPCzTLgWOhQa/QSdap6AkQ
1UfJZDmBgw8W4ED+Nt3CPAJBGnJ7oJgcpop274gr9yu7Wt8i5fnCekUEoA0iKDDhohNWodAZkO5+
m/T/CPpMZfi8iIZmO6FCviMN50h7Y2dg/nbA8a1N5jxNzgD9EdRI74ymwPuRS6o4P6O/ENIMuGyd
2H5xNEvQNbeolUheWOzAkWDtCAozEI4lQFTU+4xzoajH3hRFIC+BFRVWYBzt4sI3Kbt1H/zCztD4
22XpyFojI2B63EZU2Rlkrggl472m3NLSbva9mylQ33kHjVK0Ihfeg7Qaix2qXGXCY0DbjXlT+DuM
FqLnGL7yAp1HRQtiMpNYoarg6HrdScj5L2YPPrwGdDdAJosIIuOUQV2fsgG8oS7udUO/MNiBnFTo
MbsqtDHN91WZMuwdi5D2oVNaO16pRL5mBzSa7p9FAfoRQHKdhUZOPj/NTrzYo1wRb+Rl3mtiMYRI
7X3wonNgkPljuxz9NxcaZfDMLXiq9sui5ZqP2dumywtdpEPgAnMwCNqY1f9XIh9aakbz44R+Vfq7
eyYjia05o+4If/uEZo7djlXYso0i20VIqKr7oZ9pBuDXQWW/K9/H3zx6WTCAC1syi4ClqvmBKTW2
oII7B8XtQAtThbcvhx+s2NwSiSOh3CixGUOL05tiWowCZ/PC0oVpkqe1gyURPHJhBgGzA+t6T4d4
f0/LAXxSYl2Sxfkc/JSEW5YRhTKZIXORhfyDl3MwPFvo4FhwGX1+RTV4DYxHX9JjWUYn0Av6yTmk
950PhA7RbCArDJFtjdF9ME2ZsyyUQSDq4xCCfAVcpHBjvxmUPVGnwa1z4nZ4SdEHz4EjKqDUyylx
bQOVt2UDVe7G89rlxGxv4WjPGAWTHk86rTEE0xG0Y8icvH9pFPJ9rnOBAlKSrVRCdV/WBWhbHCII
EftkEe2Dzd0tDuevyRYaAVWn2nXwyZ2gS6BJ8G1pK+vP5pFOmYoTvVAGoHitotHo/KXIY0XCV7qd
cJDuAW/poNiaHXu359LPHN32atSUyVjxm8RpiMSnj6UmERwDh7CRdO8B3nQel2soUZJR6MKhVjaZ
nwD/aC2+UhZAJclFB+JNEkYnJGbjJ/TBB3DyePIjMKoME2GA6RsHIuO/MjedwteYaOz6RA1dkDd6
cg2QQr9ZKXGtzPuKk/KUVZ3sWZp7BW1WLqvGFor8Pf6Ryexq2OxI7NkL95NDUpKssb7o4rGASN2D
+yEeb/RsYPYEtfRUONE8A0E+X6kE0V6qKclMRZo4+hPd3MpM4/JeWp0IOQbyvcdHBTjUyWr64ZqS
+J4AgPFPn0MaeBocdECW55KEfBkTZzBUwjd2GWG9Z8hDsRDUERg4yV+Gc3D7DdZgHNJy4vY9b1fQ
jX355HeCgmO71Jiy0h1Q6OD2rLfsjbpjtXEMImUPQRYWOFgjIlKKKpXq5pG6DFQNskadtftlH0T/
j8B3lrQuih+IW9TP68CkYajyDvSdke07dWllkU68GsSk+zjO4YWZaVmhR0tLnTh+BPhEieWYzm8h
eHMglwmOKMGYfYHZXkKu1FtQH/j7rkXsQzwBXI3eNF0EH56ZiGUH64mxS/mYghWBKE4rqZr/fzjQ
OVca724QB9hd4mey53Vjl8CKRu0rW9P3sOxRO70PjeSdqQ9eto3VDFIdFSATBEUQb2+7052XcH6K
NpxuVxiYAookyP/e5KtWJbFLV3uWC2S1l4N1FNsWxg8x9iVjubFklgwe1m2eg2TfsSwLhWwsjNja
hmQpqrTdHxLn5bzLdOvMm8OpbCplbAl0Q34YHdjYIfm3qSdrdit1YKQqB2Qaukq+kuFCdG+hdyAk
0aV/BNNwd/S+tksgcnJCgX1fe+O4veEvLBA3UXSEPnRSGj/giwnydvCWaOIh69InIHtr4BNzkdCw
8shm74PSB2bRJI9m7zf7PT+OFmlvwg8lqne2spBxHSJExoMsa6RUhO1Yk4ynyVX/ZHKEBs5zogaw
XzyPxVWGM0M60otKvvqEV9rf1BJ0zXBXri/mUaU73EFPqVVfVXarEJ1Z7gioj7rpwJg+NFCcY50n
xTjkLHrQBgq2DMfK9/VmU/Ghd9zQ8wWUQlF6i7Yh+WwtPHyWID6vDayM5kivULfGK67NwOfLH36f
kjQCQ0plE0/pTHCGIZNAA7LUDtk4wCNhqlyGbADPG+AX+tns/WZ3jerv4gKQZHGpw5dX1bWf5uo8
ChClRcpIz3FGu3/mO17MazJlLNSw47BonRRXNK+1iIfEU5lR3SiHJvOgImODKiUo7GKKZHcR48y6
LRFkju+QK4Sq9o6VLRPo6sRRMdkEfutDjLDLh+iCd525embXOCIe7/wTIWHfxPBppOujqeFI8hzS
7ezABmYuu4zb1gyY4tc7h0WcMwAwEvhnXq8l+EJnQaIdjzFKSahuawIpNOpk2qjfKokEFb1QqxrM
F7VbfImjBmwCZs5Cw9L7zIwf1fP9SbqZhaadaJcrGOZdp5pGoJR2L7SZhu0IdnxYqkMa/ahW31Ia
2hFE286AtUa5tv1ZbMcMSUGE06goPfhEnBrHv+6/VXdf9CYBAb1IoUg15R+xAR9eYidLq98cAEGM
5TQwL6uFvWIfOua9P3gmPV3Kn552p4mH1wvVQy9skcp2GLOLv2QsRuCKjTcm1e0xTY8oFNqI2ufy
7fTJFHdNeIHT/zTNtj4CjtjfUA4jwEbjEu5IP+gfM0mkJMR2W2uoH4opcF5hqTqKkOQj10EGfpcc
xG2eafbUVOfUNakMP/YIIvONHyHfKpIj0JQiXHQ3tv8BijgvVsNaHV/tAYWmNxIUiskdKE3L0m16
12MMOCiKu5/GBi07UK71p8MYrIRC9rIWoRyV9nf+/5BwIZgDpJ7/xVIInuAo5iQ3NLKbWNxd4U7F
ihy5tcmzGhKsYwsZA4IQ93msucOK6O7gKKItld5QUMplT2jv43TgK2+XV99GBqDCf8gK1h3D3r3r
BsipgG+6Wkq5r/Am780PSiMuuL75nhI55Xeldb3rIzHeVgOhCPCcLNxEJqs1x32EAFWd0xeWQMkC
gWlJ9IzXYWzrOeOB1H16HssWURcdkwSSdHPhFpA2lGtfXG0q7s4zfpmjrLUMGlR2ONSnRO5h0iDo
TxQ0IBGmj0LOSElpWiufRhSUAKfKS2gZFdWf8/1sJV76u7fH7az9p+cFs8NLokkt0lpr6JdsD/2U
H0t1+oyPoZXL/grxGkTiNN38fNxTMF/MnVWQcBAEBp7ccADuPAExTXezK4GlBwPmlzDOhA/olZLc
IEuy2h+cMtLodLZvFkrXk0DqIAWDoNljFbcimrNSiQk7hBTmXOjZcKZZAC2n9w0tRKr7frAcKsWN
+VzMz3DoD23pDmrRcNcoOv7tWVUrx47v0CqW+BHifKXYCT07Ma1/30FvAzGCEgfc6cbSxdBN43F5
KEmZlW7IAnmj3c7ugF0ogXytDO2HF+qzYydggF9v95hL/quvOwQCyPGOPbsD/RZzkslfDLOQd1Bg
SE0puezXQg/zNYst0TGYo2VGZGFpqaWEpSQ9SXkgoD8SVYD4HsjyICFEvWe7NHWjnmDvnXgX67lY
2fwqtdPw//745DFAlj6Jt8l4yRGsRl6Z4IxAyb1c5nwy9FNesp80b1CGkxaJyPmnaHwXU9gbyIck
mTGN6EU3bIkrj42+IOgfTo4xTWlJGwXt7XDT9SpJw6F1j9H1DkdVkPMzF20S4A4ek04xLEJ4D76D
Yg3uSKAj3PYOJzvc2lCf2TFdlDtWeiOCMjtvZ1ViTi7zq56QSJKJKufyokaKDssbk87kC32Gh6oa
4Xyeq1K+6KzVHCvRsb9g5LMIlQ3yLBaUqEcZQ1gddcv5ufTqr6LEPoV5MGq4webovjZ4shf0vKLR
X7yqRR37ERaQx9a8/7ROgwxT75yRxpUXaM6kvG8MFenIP2B/7mUOtp0rQOdqWQOwWeg9XhukuDG8
9W1eRgkjdlFsmV1KSlaG90alyVZ3vtStLxtotCq3y0TsLOh1CBHBIXhrBe5mpJ6ofPClaXmhkHMv
GQRNncI5H2wuZol5rhkNl0/dMnTftFYoDY8v+AGuDR2A/xSWcGlubeB5mJc4PZRaR0Ib/kYgTSNO
WAc/ApfbipXUVuM6aQ+1HhwlDDtBCuyVjLMwixnjw8bZLX/1yfq7B9ajl9Ojo2jGnKQapsMS3uUQ
x2RCuj+Z78emgAKP8m1t/50xQAQ8RqU5rsJ4DfxFT0J8Legi/U0JExGXH+ME991/4l9MpwkXLCSZ
UGpZCZBM7q6p/IsK8hJ+rdEWUekVZMUFCpeM10HDA+HHOKItSeOD3b3v/Cvn68x6tyLJbKzwo8Z3
X4ykvIIz9sLtJ9uzM+xqJwHz9wuMriOJPx7CATPFqJYtpEBBE6x7Z90yBZczKvidKCZ924Jyffm+
rTD+eOXVoTveOdCh+x0I4cU2ETjKimkDRRGoQF1btXrrwfiILmdVG5Qr83DLqsD9TLAn1aCFsGZW
0EmlRCl3p1B++aU+u+NWGJgUQXAM+N1fyaEcfMrzk84QulsOYPWmwiu8/mdOKcf8juxd1BK49KB3
cj1rXutLLodzUFwZSxMEYM5MxGsbCim/vLwUIYkx7+WATyWHs4GFjvI6nUdYWAqdq8mNFvBy2DEj
BX9vh/kB/wnsoOIajNOJE4RPxXk2FAc/qAX8cNJn27WN43lKy5dgRkdXijmBIKY8M3Mjrv+Qi6Wy
lShCpaiRMkS/gX6uAtuY6e9xvZ7v3kuqy3PPor6x9sAEyAPErzypyZljXyW6xHC+aQvn79uTaWy0
OlkmnfD9Ipsx7ZqnFs24r1aBmqPehDWiuxXhgGTWDel90Sgx3FVXzgS5gWfnggkMYT9fn0Zq6uWW
stldB650wiX5DYLJKpHEPSExz5Jzwy9Ju5Yz/9zU+VYjX1r/U84+GkRj7TDveiurITqsxWFpgOjh
Yt2Sjy1XRCGLsnL/OglPbencnDBdhUO+VpNIzm6B2bCH4WWzGkVDUqC2/qjv40d0megWVqyLDZYy
6r19d6CN8CfVD5aM2e4vFDhR4A8q0fjsLNJG0nIYJWsRy3HNtWgFwbiI8nSokaGyybI/rpkkFJK5
uEI/67O6yyrfj4voHfnAsF5DxJwcEX/GionR+Vdzdv7aTpDXGG83ITfdAW56vfO65hDggHc7JHj/
ZFV9duT7b0PiOBbi/2yJK0JlKiEMe8NRqI/Wiu76Wk9IUNVmT6EqTyZh6BOjHu/jNYbDPDCv8bs3
8LqrGNMw81119kq93xgoEcgLg0dwCU10ZPWsYl37ORnYwzqrQublR9NtPcJ9mamUNdV54glKG2Zh
3h/kYNRg4Kfqp+zeSld6SZ1nqLyXowY5qR/Rk7Yq+JkGX0UjmdGK37u4wxPsQ4Uiur1tIl9yF4qs
R2l/yGjGzkvujT6jpDMRaa5+TpSzY1gxoqyttAYpHAfCVFkmmYC3ieJWa/ATjiEmWlpTOGBGBEkG
UggDeRrWq4zGPbLUPo4pes1kexQnJoAMb4s6LDu1Z0glU4XzKxXh9hLMmvf9ywkIyTrBiEKyfFun
JRRRVOuoJZRghbgxjJ7k2Ub8e67kXTJKuIC264g3K5kE1dy7cyRFT2hOvpqzWOPuBM458ts/dQUa
AH4/lQkR4iT8B0KkvqwjxpMyzLLeOGV8UmczaJw6viKLJM0c+hnTk5jjG7lJUATgTbqxN+9hn31y
CtjWcR/poo3v9wvXtECujXZhkpZt0EdT8GZetrJj9VCF5N8+jtKSf43zGhmf5xbTKCkw3PE1ccJq
AHY3azGi7OEnZp3NmkFO6pOuKv2pTHDE7xLBGPy2ABL9D/jrVxL65KRKrMPPVHEEe7w22PEcr+JB
vlV9fJ22NRbectjTvJ9ssmGIoRFRxzSxtzZ1sL3G1fevYJZmiB6ZEOWnTaxI4NYxowrl9X1fdVrE
qRs8bsg2g40gzSCYKzADFM8WkB2XIQNTz+aEErabrL4mSgMc51AMuIXBwEUE/hYc/mZhbJlVsjoI
nObPtKjPZtN2o7RSv4R5cu/jM88pMtD0pwrhW4lnUEEnR46PuRydUZo/mBYx6FGc68fdQLAiObwA
usxXoQOGYCsm4sg11LVgzRGo20C1y7hR5HMD8ap499s2OD8HLPUUDMdiFqGZAm60yBNBdon09yMB
ozY94is7asoh8u/EN7/B3ub4GJpamARRrL1dk5+bBWh2M3pEDOt5HpeJUJVXUBGxhiOFBO9+u64p
0KkE1Kivs+mWUwjVd/0a2xWTP0ETPQx+OjeBNF1P21Og6IauyuKPzZbniGqdEVPJssqw6sfgteek
ochj1gYvhQOrmeokhl+fuDLx4kQaxhNW2sjygia2iELjXGwq8s7R7myvUa1bV51jZ4k5bkLoBC6O
ozSL+utdZGYmWqb59EOn9LeCoNnYqe1+59rxsgb5qg5aoo/swO8dC2qWOde1Ql0LmBog9qHzaj5b
yYudsKLdFKn3KzruntmJBrpaCJ+Xs1KVjezm7alznrz+GfD6XtwAXbF+y1ZcKrE7OiWdO21hTB1N
8Oy4/wdByaDCsQso2tFpGZ2R75a1rYS7WcCQbimasmJ1s0aHkT1LjHTd/ErjmZUl4H5VEzWOtTJY
gNupbznyMkJxXJ/nM3D33TRvclWvYZV6WBFBY04E9MPCcaEIEl2w2IwdY/FH1Vug61yYBw8CpuZs
R1O+1yDFpx68/JPYxD38ZUjcWXXUEYhlEi6hZ47wqKlbEdZT+OJwOeKj50mgNzDMrNGh5sQ6iI6l
3LjJJK6znQ7dTm4Pill+Y50nURyOSNqWNc9a5rGtciP24dknA96Aq8SnCe1fCcDbLxGfosLIUan7
E3BrPLdvJelAswz5QogbD47esIwpgtGqyNsYYJN4Md62qsXFHejRKR2ryX4XVMTSaYJ5L9N+Wemb
gDTYSw0NPy3ooHKLPAQgMioFk70khAT9FeGo8V3P6En90DHUOKSQcbcYGt/PArVcaQbSDr0iOdwJ
gfwPcSIG6NYtA0IynBxWhKRYW+atT3FvzVM3dCL+Jk/iUr1wLyqbyS5/pHcTVp3FO1Fp3rWOrVd9
NwV6VipH8CjPIuhaILsFhQbXbHwskPRcB4ecMTsc9g7tc7tRiWay+UNO4bLVFQ4yXP3A8Dlveywz
QfLJr/iGmt/e7SGOvaEa42NzI29+e7jtq/IYDycyHHFGDVYN96H694+uyHOLNNt4WaMrU1brRgWN
9YL0HmcHwN1SUMAqBQizaj4m6RCDkoTi6zjGBhjWM3q4KrP9NzfwfLYYg/3+5wFjEpM53nolSJ5n
51jG/lAKYsBI2dvOKZZl7WPnmnEDvGz8/XnyFNZh0K3LDVA8wOpqsPNigMrlYDD6H4bHcPyHhOxv
jKqiHhvS31JDbO887+bqMYQaQx1fcEe00eID19Z1DS8T478MqHWkNfZo+K1IEY+0+g1M1A5+SkAw
j8rtrKtpyTtFGI3nJZZ+MmNwAdTCPDL1jsN4Q8W8cl0LQmizGa+BYynIIgSOab8FvZ80Ly/zdSj0
Kyv2p43U7C/az9Cv1sQX2NOWzOQABafblixp+ms8VpfuTVoaVT9cWmVMqHka/jLlwaPjgNy/PbqQ
VfoIp2wFNfJsVJcWxAbWmaAK51rw0gc+yYNLsJ+tdy1AIEBloZi7dMAX9GiX4s9bygctb2dKialc
ztCT289sUtL3vPsvEEntr3uIo37t374ZLtAE9RNCjRgKrke0J5rORE2LUWTUy8sMadbREwu9c/d0
UDfa1AcUVp7JnntjLzICca869eTZ267gNfwaJRlG6bpheuuN6Ai9XwDyFZXkDas8dAlhq/lwdwJy
x26ggX6mNihkPwcHGqFz4x8LBCeKUcVyzDjb3/6Yj9I9RGsu5+7yth2Za4V2mjZu2rRDoSUe70Pu
DzfVds+wK0WziVWWCZzuLZWwdwMAsPwyAb76Wy0F2d852ZcHO+O9hNUkXexmeeAOek9GPPLrKPJQ
MOlVCCmq/f02AhY4Qqd54UileEQJ6OKCWMqBG6eeO+A3MqgZY6qpXNam6NaeuKLyhWNZXmoFX1X7
r25x4V4UOxuIiBQH4yETytxXFMTw+QlUvndLxP4l0fCrDEofS2jiC7PoyrMzJrjWN27mxyT9ua6X
t1O/uJ4MUVuWckAz6r9y2ZPmcdD4CfShS2EFwsyWbb5ki3sniWnwnY3cVn+kdtvYm7sjxWCdjj8p
Xe2QHZyB3l3grQrEw9Afa+MikEHmo+JDv+JQ8nYcQIUYR7U0IbO8wJSdD0BaasLyaBQUXvYH+yAn
GQ6Q7tOEB7n3igedzNoiacJHPVpeZBgit8+UWlYo1eHkQlzBJb/ZE3jdpwXvNejFlNFkVTcuOElN
vmoK8/P60VA7Pqtely+Q+Jgmc5itFbPVLMA37CLjRKCGSQwUEGnpbYMZlg+CRryEHP2cwChjeOKw
VF0CVIhR3oq++hR5ev1/2Vtxmph4PI8U0vR7u+bsI9iPW4Q8nCYWSI3dcG34vo3XctTf9Ow8AlCU
Je17C4XQgoI5EiRrGRxnMJtxIjLRF18wbMzMPCOGwDYVmG73yEzKBI4BTENMYx386/Mzs5cY7VAO
cxLGVEJT4jd7gY4S0t4+xmTcWclFTA3Ic/RzwupJ6NBat3RiBwuZT+wua+STJt4ejQVQoaH/coQ/
2xNWEjNLiCs2BSJAf0UgSTVULiVREgEYkry7RBSZ3AiQBvdw7UN5DQH63KFN7UBJxBSmapb8el2o
y4lcUxwYTL4VBH/Jtv5sbpZ4wwIebDh5b+tImMv9lttf6TWKXbEbccrgJ8iS1CF9QltpOaHKsDP8
JF000+1CvbvHwrzqKTCEu/oURous6XFVp0mqumvVGo+gTO/UMqHw8scvrCveWcKotoOyk7IoKcrP
ggZ/6/7/bKZcscVfrMGzdG6wEHPn+19WtSgKuXnqbDxEWeTSXmKPlAonc3BvZ+ke3QztCuPUwZpp
mOMUZKW+OGkax9+9+Dp/5k8i2q6dFKLnOxrYPcRrDD4hFaAWETG0ISQzjCLwEOdUcpSdM/Wx9Pfz
2OU9MkF34LTPD2ZqzcticBa4yAnAeaXTV7dCjReQf1FdORgdg75Pxm6+2ciS3kQd/4ExAb0Z6KPd
ybimo0pMzgVYPxxDZNYpK6pc6TNFxEDen5utk5GlQqx/gqfVzlCQnA/k1F4CcFDKWO7jbByNqt1C
1ahCUThAhArusuFeItO8KutwZNw62IvJ7x3mFbMYi3I78tNrux+HoskN917Y2nw11WQ3K1UaRcHN
18CQbjXRpagQ4OI4kixtWiSHSJ6sj/KDAE3yTwnJFLTzZBireBFs7BpDYE8HT0DdV+0Fn01dbZtb
IV+u8m1wphqcuhgVQdDM8yxp4OGHuMsbMLCvMMpi07ohNUlvNZDo6n8cgpK8td96bPe16X3s0m2V
c9X5b7B5UexiQfiml/BSP+sozYMZEH2g6w9bOO2sPlq+2prn3yZa3XlV6yS5DEirMU/fhgkG7wbj
DotBQJplTXZtiKwwJXaPtBb8Kx+5I7eV/9WWVs2xTiK679FLsMB7oOxC28ZNgdZZ5hTZ2AEoHpx2
fe47MMecEK3VLqNyZlmgqGqrml3LvvahevTxo4uZo2Yf4v9bPeiYDiXVuMZ1nsgLCyZQRgjSM9LT
Ow62OP0h4/cRCvG3HbrISQUnoZrGOdQiPEACQoWw9C20y+T7p4gYl+FMHxYyI3r0WmiU/BNcHCZj
jxFjAWLCOj35en+rUK6mnhBYdILe4mXq483gEISp4ZYZjtZRFBEip/BfQUEN8vxzVnOfiSd/2H1S
TEQxBvzaz2+HH5z5WcmZBUSlN006KWTqYozLvzO4XxoPSt3Ko2B8OllHbLCznnH+3c2i1lI+owPW
fjloNJaM2PrHeQ/Q0EtRiGcBcQhWQGtrTvz9BVkXhNzwZCpS69Zv3m+y92qMKhFAzspx5KwTbMEE
QDT2+80rVUkGyY73VnVfJsydmUV31sfXxfKJGb0tH25sIOhedIMfOJQ+Ln0Peh6qxnaolmBJFYDo
XgJP0mFqU/HoVTIGD0yP76PUMQN1zHI3RM8yepl4s0wwGrUayJiE5I8In9SZ5twumK7w1FzUIuCc
4IzY7R+T4RpvKUyCMkxrvBVt9ygiNJnTgdiN359hsiVJIYkyZ3YNO4a3YbOkLoDtSHDugimS6Cra
ZBt6UrIalHpd8Go6GLQ2seK98FlHIjDOmosAPjnPpfRISkwMBsILF1Ck2u0UqCqmNdkWoEG+btsf
qlWicNEHkPT83a8ZaV1oNczDvENgOvQONjDTwnkoNeUh2yCP0L8dBni8fK9+RXsZlBhg6Htcurta
gfTOp3WaNiP1THHFtPPMjQgi0QxHmUdX2CKZBg7+tw+8kNAWKy8DqDD7p9alFjzdR6QvJU9EsWNl
ATnCM3wCmrOQmO9iVPOJJrZZwlvZabRT/B95U/hKjJQbowWtK3xDtwPWQuswlpOE/nZTJpTPQbE6
LrXR+d8+gtfoCO3AM1vZeyYugAmUCF2kS1xQUDEd8ZZvxYeR6aSmwKWvYHrwTv4hIDWB0kDj7TXX
A1LG90alEoEO1ICTYOGTXA/vobbE6N7GtGcvq3uDogKojWFVryP3lQ2/lJWGc0T1KXL85dEs3+Y6
yvq3emi5HySpYySIKpZZG6Ko2k5mpDvR8BLMW6ki1/8BpIwRzaz2+k+2dRCjaF2rSIgJZAPktKfn
1AF7TBjgcWK3+6eQsbC7Iqdgxz5+jVGQwsgkudRzABDMMIUSRRAHM03ScthoTe6S6tZX+VZHZ9BR
xxLoOaj8hdoQPOc1w94CI5Pjfm9ZFox5miDCtZc0LE3ntDqUR/J3Ih0j4YYNTi7YalI5UBVt9BBW
3z1S5uGoTeE6/gdQdhwsBUboIce3RdswzCURmibmh6DxNbzPuV9CEIi8+q9lzv9TLaFmzAgVt1mk
xL8B+Zyh1L6QHex2TRJBjLtvMs0jKly/flOpKh6PZlg8O3/eNKQim9nPftVWV/SKEhEdg2C/1K6n
BrSgHA3KjJcLNQXRGvvNShQbP8DGPamw9+IKJD8eGB3Y2UlsktvRFc5I4xXWGVDBrJhemUOoWpGJ
YLxX5NzkOAIoXEYD0xT+dEFbWqOjuT7HbCgiDlsLUcrci5lR7qW1tLrA4YdUoIQC31hg2l6N4HKQ
KqcRy3kpG1Lb1bh/3OPxUr57jrkR2EQNxHWSKn+fcJ4ad+4XM3iW3erSfxGYbPpXQyrFKReoo3Bb
w6+tHuYVSMHRETatOZihv+09+xm5A4sYRffEVfdL/VUMUYFOV+SPlFfW5H7avPBuJIlYx92vNuF6
x3Athig3hKrh2TUBxdwnYiqyBGopYNqqdw8jI1cdl4hsXOIK8L7794r1XgJZS9e/7EypppoJN46U
yUzTP7Koy/RyxuOurxvXTZsADKO7GsGHbTEsv4rbyNJDsK4uTW8/ZbAR/49IxfUH7eG2Z7NMMWAT
jDIthY7N4Xve3S73R0aXH3keKSmO61MxOLxf5nQNlYVqW7+ww/FxEFsKwSL9d4E1bn+FLb5DIJwE
meH76nlN1oklodaPyheY77KPlxZ5gIexdXtyebRWvOZyCRrgavhHVP9/DfVyM3flPDiJTpdLTxzN
tnbWSEbLh8TqBYh0msk8YFPlSYjze8Wrpj/BU8YyWvJOCtkT0So7XKwC5Hxz9jX1upmDE5uUdcvI
Ns32Dtfn/NQxDGpxcDTowXJrpRFfWpCnf+Qohp7gF8YO1dcxEjcYWYz4dUK92pnnnF2Q47N1xKuM
yoObPlsVUImQi4bzRDUleqpFLu9n/I3U3FJiQxBEEI87Tv/hfivvO1lQOO2fcqTLTRIrdYJBG5CT
cVA9DDNbwuCBbZcvReTiNXvsk+zbhPS0qgqIzua9e4r32uJK8Hlh0BRQHckHKeiIUVUvyPd+mtTd
E8tPzQBpvuAcP/4H51wvNsWfwWvG1Wy5gBxdlLiynE06zvLU7+HFxF+dJzTOOQ2OZwkX85tOjSn/
oGzMipZWTV/VTCB/zWBbR7xjTt8nUpq/3yYrQTTM9bjE9iVxAQTOXgljIrxsQjNMOKgmEh6u0TSr
Gw+xATZUjP8wEhyY1xll7vUW7plJdqBKKCmPpKEoDPcePCw/AYdu3poqa43ImHv4thLo5vDMCctO
VfWejoFqWhT7RRqNHpiUjbjyPhN+HnOOdC3m9CwSU47OSqrA4D9vXtrjdOfFMsao1ov/AI7X36b5
UgCKYoehqbgneh3fffFY7D+bY4b/BGq/ho1w2Ocv1+1BUWKD+xYCPxP0EMpfIRLGaJ8mXfOGKoxS
NJdtXSJ7q/vA0lB0Z9QjnUYnfeocRNbajK7ia2vp5cUue8A27/l45Z2LJHbkFTTQ/DLeKorzgQBD
8lJklhcbzlo6ap8LHwmeSXbxjFIx/sOAd+JMAOxokrJAIbI3aSvBmsWJNvgkiWRoMf8p6uwDdOTx
/l0x9VgbJ+BmkXlfgDkqLbgvhnz44d1FLoOJ2uX+vmg0nwtKADPf26ZRy/STFjtHcYQOsmSCwRi9
SSxwb8lGMD7iEkdNC7GePLkINbs+N+iSXjNNwEhRJq1bx8VpQxO+Asv1/+MwdhvGC/R8LaJ3x9S2
rT5oHgVUJHH9sY6c+DV+Yt+mCynBYqZ87TyKwqAtr7MVKKFllg77TCZmQzW+MtBOwsS5ctfEaEjj
rl2hh0e4s/e3SFUZhON2KvAoIkB4yo9zF2olZ+gn1XiChXGzB8abEpEAqxrO0t2odl927bIqed1c
DiuZRzDdhcrwZsMEoVhA4IdIrNwXgdDRRobNDYFeaufDeZNsZsCuarDgK+TNGYVfVUwW0nvcKWZe
bimPRux9uQI1eCAv2+rO0ClvzTYI3U7kbDvzBrGO1LG7CIuozWTkPks/OTVK34+YKD422go7VdTi
r9D/aEQ0foFk8z6EBXkTcLJWsiF66yTUgvR7LYpLmmx/SQjj62ZVi6IrQzO3KrhZU1seuZdw8U+Y
YRyWnQuMK6VYeXjWhz9EM1HzsvoxhW+7H7jM76xettItYAMKxDs09vfQCodIlPy9GvOUEbO708jB
tgZAhaBnhH3xm9DueF2D7Gs+7focnsNBmCwmY8Xi7PJouYHIurkJSYZ+EAOD4e+K2JGCbrKVfS/B
ehuC72hksh2wbeTBhAx+XYr9w+qhsc53pq8Tp9CAROgNGmVN5YZTlmZDh6xXi0LPC6E80xnC3pUL
H9A1wc3duTg6w8iFOgikPrylwVfipc8zXt4mZBYefR7nS86q/wABL2xX2/h4A8VYXv3b2NR1PHcW
b3UZPQ1O+2uB00fV2ZJxuI4C9i21plkklaK8q3RF6YftXXxN7GKDdkGYrUeWm9Zb+dx1qOBQcJUM
FKLL6VQe4Y+XTJPJnwVpr2pJ9dpV72TKaBlActOErN0LYUo2DxCWbC4iDF682EBsbg3t4CRLXQoq
Uej1wTQw+UwOY0dWh95zQKraVzdNOnbPaoQSZnnunnUqlLvn/Gy4F4wi1phmr2bB6+qjRPUfnvT2
2fUK7QAmoZoL+vzLRCtoKIVms8ExnpzxbfHgL+JXDIHDaMIr93jIJDFCFfKOtafYmrLQGnYJGLZa
Q7mbLFDNbaSPTvl3znJq4SVkCFstsCic2508XWvHlZ7wwt0V/Ga2YwXgC2T8hf0MqqVb4RiI6Ul0
0+jfbmdieVL7bBaFzOtZRqQ+/jPHfbocfGGVLxbwd/YcU1iCmVs2Uq/6/0EJHONKZNcIZ99CJUb7
M8X4tw1qjsUywBPIuUEgrqgZIul4svvbYAhaNH/EAWKv64ZPqPaHU2bsQDG0iSEO23JYOmnakFwp
iREIfFYBaF6jYkcX6aMjQcEogHywsWnSpFaC1A2zyboIJMVr1b4RrXOvGWT674nWfr3s2SY9m3A8
22RFviU3ZoPx50vTjafGsBri0edZaFATYYlx795BFiMTyS7roPyYm6YO41mdKHQtR6stx7Y+P9nJ
1d1sEsiQXj8wE7vemEc3LqLWE+ZD18v/G9YaIJ/JQ7BDgs6w2he7skla0D94hvOxSyFzMKQz+bSO
sPJu4aiY+HPqXbBWSQAzPDLAHyu+xaG6PdJeDDFEW2YI+6pRW34FbhSmIHC2AsQMisOppR6ZKHMl
swULFAQUaPnJRAnDZNDianIsX6ovr71By79VwDcit36BHsUMEVbQtexA/fKGL5nM2faXA9lDHzcN
5V3urT0lyOaRARYZ3xdbEjNMM/ReDe95iUjYkbU2HHL5R5aMjAQ7bLqlxc7Odee7PJZsdTWarLu0
MEl6LKW+8p1bOuM9rIi0IqGPDch1qN6FbFdc1O5Fmzk8Tkw9ALbhqmfbiZR4Pc0H77pGVEN7cuUU
/ZrZYOABpXwjm9AJz+XAWx0CsYLYEhsCOwizJ4RQc8AXsHo6tE+4vtdkisZaZDg+3i5h5W/dcDfb
h8VC1d50Wuiw1/75AKHz3sZeND9bZhJLnzRi8UslCnM369M38EdDNp9IsQU55RKSBdVWF2R76Iqe
PHmAvTSr8nBxPnWZWCDOGtVlsq0BPfkiDSxre7k1nghQ+C0Vd2AQY8iqkBBbc31IWTyZqAZaWMGx
XoDwCrk6KfMdS/cgaolZOg9wf/RAACXRV7mwQMev4Ikk53y2eSASqgZkst9/tcTYxmqHGs515xoW
OXU1gErWJBOt8UrK8zxVL9t6cvyiZZQjdReBcZPLnFLqZNDThMr/5lIyeu4CybJ1bhSFCLvWquwJ
ndax8Hnnb7Jt0rJoKCoTyJLXumS0/pIdLdByLuD/JMd42p0Lf52mWk6dJyskAnCmZ/pJMo8og8DC
yEWyokSZV5LTeow/were1WEzEs7I7k5k59Hh3+TtsqyekXaVOGf6yInWqh3U84+Pvg1phYhggBCa
ei9klcFE+M22AA6FwuKrWwWSFOxV+AWAXviU8KXR6rzWlS5HHCROpfZMb7lhSzQqLSmd+6tLyZq8
x0/dsxS13HbVx+jSaRjboIEWgYm8Yy98NUz6yqo4F7w79QPdncAYfjcYU+32202WqwYUsRJCh4g0
FszEszyugrcH/h6rP5G6tJ4zw9S+PkiBK4G5nf1tlnjnNl0RPN35BD1xYtCA71fPv4VmWm9g6krp
h99APx5t9cAeRANdPq4s32G8nCJzpu/zpdjD01k40LVP10sLF2gBDOszI8+Q8FwPXpANh08cA6So
gHufsbgV/CSOHnSEHljSgq0RRUgbL1iof3U4/Qc4p2QZ6WkBI/6hbvECktmFRV/6Bm+zNmLQiMvz
5baecNEn08hCNZJ/1ovbD8sq/StT1kaHLaVspxSuP64X3d5bXuCPpTViklG2Gra58+3H/KrTjoMj
qYd/zv1r5Lrg4TIebQIWCBG9fuu2jdG3I0QAgD6bCgRFacWbFfc2stkb+uQILb+DGXMPSVpNSJ/f
Xz48/t/VTHWvmGB9Agtg3njOGbv+JaDAf2wYS4RlG4aZkOMF2BIbwHDRCZ4S/K2zC3vg0ZevN+pR
UKQdH+i3eZjOS9XbDW/s2k7XxXOn/q8ceGuoaXvXBhHqX0jgO8HAuTMFC9rn92y6bkTyjVM3fo1x
+8xiY1lECpWcwli1YHzeRcJgJrYWJd8Xv7uYhr2qtZUNANvi72xDnRG91AyL9SQvHt/TRCoGMhIR
xJx6CqlWYT+KkUSPHe50ZcqJarExQQTviMIu/GuvCEYfezkSftifIKXdXxr8QzTCyczbG0wXhSgu
D/GGSxjZZvo2Csa1Y3eXjqJWjUxrUzQE9aIAtHaafvrTMEB55N6OsikJ6AoefMq1UhlAERYmbzbF
Z98esm6DcQba9gESM8l/TQK8Fh+kWyk7ihUxtsGgmFjJMyva/RUNmNA6BkV+R3q4nLFrsCOKCyiq
wbD8Mh2BjOsTrXeq9mtgtphzgSxeZisr038+bfQwcO+YKve28xyqTGW6jCUPpG9yPEXevxv4CXUZ
2L8K50KyGIYFw6c8BleWsjRy3JITUJFA2MF5B8kQLkBLjFnboxzsH7tcUFYfP3x2nnoup6TS0CAu
P8MTi/0qFSa5Ji2rtXBE4sVNmPM1ldqbfKF4+H07S+y0+T/cnNWh78PK/UY+Y0kc0FqGgWUf7Key
rQWs5muNgjIyOjOSCwPGZJJwc4yTtXsSlmsfUNJfwvH4eUIXLGEb5u11mk5HsOM3X+2XYU4JUWN+
9w9+ztnrnm1sh6GNL+kTDFiFgw0Rgh6TWkl8eaH3RU4eRBcqDu9mwclo2CnAbEi++XkCkt4M6M7z
bW+X+gt1178q39p2cCwduxZM4uB/Sp3OjefTKTYLYAffZvTQFTdxDVTag4kkUTHj3bG8O2uqiFUx
RLSFzuWIxweodeO+dIU1O/gNGBuK3DFwYfg7+2Thq01Obz6m8chM/srOXow8omXqAYq6ewgJce0T
iijUNlowx5Yefl4BlK2WHrIHCWI4n9Y9N7V1JknOI6uZEOXnDb52cjyOR/F4Jtxj7UnaH9VQD0va
jHD1nk++HCLG2MDFhof+OwMoBbVuLXellAu7DnsLNDHJS1Sj2cxwheARJIyBgeebW+qgR7VdScpp
DLp9d036KtXjJkrMrXIqZETi44moB5F0O9Pw/0Ims/5usaOClAkvfOZWATLfxMwNKBrEWWa+d/V2
l/tiT9Ygi2mA/CvcNYtrv8axDYybKfou5R/qmExTEk/BukHk+rOD/Jruucp/8hbrzyOF20sl3eeD
MxoXc0D5S/8D7PRN/hnrxvYPx+2qS8N0km44UtjV5eMHiWBclnCBZSJliWnSzXqcBW/j9wLWC8sN
eN+OYe9rJgRy2hv7IcCnV7kggiHANV4RQ7gFH5r6/W9o5iNwqx6+sSanoJnGRJQshztj5Wx1Qi2o
sAaBbxysfSm1x19T8ETdhtYasdHlpyj1k75+s7sjhGhYjexyAmgvHd4MsdihP8flvJnXetyTHQI1
/s23tbADO9EDF7uD0BcW0m5lORe3K3TOC64o3dOWSpdCYznIzdToUeGyMKL9DBB6oeQJyF0ymluM
RyBJv/WtYY+7MsdK1twBHJVkErUGRsBgP0yx6ndDEFURxVF1WofAPgAa5xJrOl99uiu7PfBHQJGg
pa2KRRWYmWQBDagwF8SSg0q7DLr2HtaH0rRW+GG2b6K9RRCq/Vyp7p9DrqpXy2m8EVMZ1PTFZJDY
xp+ej43BsWgtmor6aGT+M5duueooxD8YRRX8fy4/OztSckQwkuED1C/HMs3OIcD6GWMGGGI3lHKD
qnu0vfTHuOWpMp8N5vqZ8IJt5M0QFR2wdXAZ5rw1X3BLD98xsEMTqykDlYkLr0qq9qk/D7sqgGvq
PNx/xrZ/8i23kuO4MR0qG8Oa0l4Uv9wXBvqWj6xjhrJ57xcTf5OSC3VQqAiujDxWee4iNPjXJKwC
SO2lFP3TtFUMmrrxEdzNg1vm5nOR9CRiKIRRrKvkg164q6yveMD8um861XB5mmJ1sGqw1Eg4tvM9
U7w65fGrcO30IXTZc4scpJEQzMz0G8QAnXtaA4RQRtYE67764lgo+/raBZLd7buCuUlGPpXcrtPw
C9xRkJQWzGQCA7a7M74DRxzlgh2ECPGEFD3VCkWNJFwbPCEDvoE8PADgwGMr78ips0c2HeeHjji0
CHDZbm2q07KgWgGhhjGwnFpDsF585wjcQM/dKO2Kf6+HnU6ltgCH8kJzRHV5CPfVJ4fZ9F5ct6aM
3UwyVfeNzC0mfb/5gIZmJgOirC7EKp4MFAfAHr89wOKIIaxNR+WB5Jyka3lFT19SfYFtzSmsYBrm
ANTjFvJ25iWrnJseSgmzcS7fmJuXs3pxK+hZgJhfmcGgtBtFCwjYK6cmYRcI4Xhn+jonrzgdzNqa
Aiyztfw1Ykn5Hbb3+tIlKVPzM5dD6JVMa/9WDZwvTAbax04nJzLXqHR6Q9GoBWhYyLaiK+h7weWf
w3wwvc+BoKJwS9zOdVlrooFaONDQYXH+lrI+L+9qWI4ZmpYH/o072zhul8nW9VY6cOiRSsbdOyh+
xhpW1lxP2B31VYV6n4dvHaIymvVM7GPEypsZabRHEQ9Iz/ZB/f88I30yNmVyInaX5An0AWOfy1iG
KnxZkUu4a3KOCbVVPYduqVfKROcTd2nZsD4g5fYfMBdQzbbhJhSliZrECe3og3b9CM2yv0dwyUCP
7uAbD9CWaACrcq1Bv4JBt12c552bGAw3S5sxCq3zuhS5w/Xh5p1XHF6nZYLtz+DXs8ximfVAd674
gDMShwH49t6PEyh5Tl6XBkRa/OwjcDCwOLUw6k51Wl1hQrck+RynZzIuItY53pbrHrkBa0AE5fDz
4jZ98DYGOX5w+ayX9SQlwAVH2CRZF/IzMuMCga20GNJJVgITnEQ1Y63o/Tm3m1+KIGJoSNxdMUI4
aZ7MSJpBKeTguKaBEPkJN0mH3BR8iFjS6jStuGa6DQvF/pvsmOo+eGriPQCoKsTUEEHphXPN0MOG
dLJgbw2uo/s9ZfgRsjLvzxrRj8JIkmhIzJ+KvQhvwWkyW9s5Z8Gfq36WSBBV6RjgejLVcUCI8nqO
i91BALQXUtSFn8Nad72XquV44dzKV/AfXi60fkMHZiE9xEY01eqj/SjGgM1ql1x0QUsNR0m2HLFk
NzqMgoAhOJzU8jKt5zi5HGBnzS/HbE6t0RGyfpYYJ2bJBM31Vun38/I9go0v1ljY2XnI00KAT2w1
bhXAfDTbdONRcd+WrRTVPfdXli5eQt3U9RcgUQjrBSERHeGbFA6JryOh83R/DMk3if1NKoy5PbeP
w6cRAnJoGYYZy7wibUtECX+HpSPjqj+Mgoz1+8QECvfmBv+bq6Q4qcPNb4jRru1fPftW2rnObxUe
qZTeZ71CzHSzGTejlo40LGrG6PoPWQev7tvdjWIQerL7uJYv2uYcHhMdxVzJTTCK0Ca/u70e4hSH
1P5mjmGhacKTLpmQ5UAyv1UIF2I8Usw3QqiIfdqC7WhoUWkzxGIFJu83Imypf3QitVLfl7nxRXrJ
Rs6UCbeFP/O59LdstcqSsxx8GZBN9Azd2lHSKOVGz1fmA5p1o9mXunNoNMeutYJUbN3KGF00CM9E
5qdDB93qUa3CeaYl85M1L58hdarvWADNchhZe1mXZA439ngQPpV9wNMMW83YLGbZTw+LpXUZanCR
uidkc7ziH9IXtT5hQS3tkK4cz7ENxai2fMtP9Fl6ibuWWB//w2Ay07VGB3tXx927UMWNsqtJrjRQ
8Pdpe80P6kersR3svOnueVvlFK8akK4hu/sdrQVKrE/OdaUn2qOpvRelDF90s3eptvAXKnQMg13v
PgD0tz5KTaEYEFjhPs/cvktIDbnpvb4O40+/alE+wWrcGMXfXau+7gyil95c81JyoI7DXwihor5N
P6IezsRPerqsH4gWJQJJ+f7ehDik5vJ0y63M5DWP6BZHEJnCT03eBgTRwKPqDd+K97ijw9mAdw8a
K233ptBvQnqZ2NFL+NB7yiGILrbW/Z4isQg6ss4YDPHjJmX7agtN4a1EjqEhvud2KD2NX8atBD/y
n56Tdiemen52+V2YFwDjz7IDUm0dQRT1PykU9OCMkhFWIUgec+AMEn3RunujY+M3Gi7vrBdDWy1d
WHUuwtqDvfrekXwFjoVHhiV531YqoncvbYgOWAACoAhBs9645nguI9IFdLdGBOB6rfG5ceeJksij
w6SB0JJTsrbU1wyeNetTuZyEGs8Lub4FaYeGSXkml57RhXQVWK5EFYMvlDmQFd8OnXo4rkCXTmVI
HOR7GTG9+ca3HYWoZuyhONWwSHdw3x3ewbZF4XNo3pOEJtotC0ew11tGX9Wcd5oKw/8gKTYCursL
XaX5R5cvqU9uXTsod9MqKeaETV3LUhOY8hv1Lirvf+p6tAjuxXRpCwyJOkK10/IzTOwLVf78GeBo
+MGJIbPxBgSRyI+wLSNZ9H0eA3jgJwpN/AHJ4CkBJHnBotSPKnPQ6VjcKpXSuGFSHGfifBHJX+tg
sd4rRqoYZpjXxCXdhdfM200qT/9qr3lpxprCkZm/e0dHKUUO69OH9ueOkg6h/uZExxqrNvqZtRdA
uJx/U4YO8CGdMudS751zb6l5ii1M4n/q3ubAE07PMUvq4ujcfrvBHvxPuV5zdMRtMiKPh5BfPwus
HUH7Iv674WzddEI4WZPSm5rGZp0qmjRNojrp5uvPJa80FghN9EotZm7yJpevU5e827VrNVUCJXOy
z6T8/poTKGXc6wrcRxXNFwUoZcp0iwdr9be3xKEXw9Nu/nr4n1oLHo9UkTtRhCAUgtuWjfAweEOA
1wAGQ10GU7p5y1YTyK62dPhRTaMiE3Oi5WYXogtcf+0ISLwcoFaVeDEIm5nWDmVbNgW9P20705gK
aot0dCn0L8TXZyho2oYgy8FB5LNGZ0XUeseGbyjidv/gnaf4dcN1sKim1iLKrDKUQSQoHq4U4efo
6xJ6HjDP/eGK1uWcRrzKzcyNWyioUN8XQDcONnv9hukVWEVrWVeghdc/WvVKw2Jw5ZotiKKwvEe8
XqdTZSL3GaSJDgrBFFCnXqw9/hhmBYp1g8200ucPf9Qk+OfTnHyTvWZrcvk1xu5Av0kdy5pWz5f0
KxVcyiJm41WIIXrrMgxtUhJXLhM0dlRYA6GASEUmz4EBi4kR9LtSCLP3WFqFxYrN/7nlwu7GfSfg
kP7Xj5ll6BhUpLSVXzFWl1rESEpjfUlDwNbHrTMxwtJJX8i2pnrqO0XnQWHbvFD3XOpU06ikLc7r
QSKuZHGq8mNDTSf0xs21CY/ADKTKBdPpwq3o9l54qUVusJJHngjN877vnhj1VIn6G5zLgq551f9e
g7TBfnBA27cBELXvniv6bB/QVU6J+x8KJZLUUvjprdkjpsl645PPN8vr4Zi4HZ1PA0PN/HwzR71A
2K3GavgQ3pD6jL/2ibcLYYm1+0xc/o6iadHW94eywnmLguzIqgo7y2y+y/u39cMWk1QDAc+Nwwur
i5ZiUAd4UobHseOm/gRY1u3rJ5E9Tmfhr3Xvnk3Tz3dLaLAg/cZ9xcAE/sbcCgMoK9uyBSJKItI2
GJaVlNu6z57mNln8czAm6GsNlHcjtE1cDJZ1ZhNy02Fn9OPczBIH+Cfmp30T/ImJRb7JTqZm8vU+
PyGoFUrdfTSYDnZERs3qKPUxhMHMCb54U9cIV1RhmoI3O/QgomseAAk2tTJRuYF28kzUVRkLrPgW
SMunLiKgFrTdz2JYET45L6pCW5RnrQltNS87eLeddc4AlIru0iMMM72qcHieVBUi6LwbU6i/aAOQ
XMDp1djCTS3Mae7ON+oLpYqXrXQXcvl3QPRfBrJAkR/mkV3dfaGXEh3/vH5c92y/9JbFP1XlUeG2
sgkyuLEVqA4Sne5pV1hyJAXMDqNRRlfiZOF7NZK2DrjWl9erqWDTcXqbkkyfy4sDUDlE3PDrEswk
cxXVruGFuhJuLiPtZaMarcXOX9hvfYUzKaOZqJkWkiWILN+Qnu4awZ/jRd1B+c4Foftvh8pwZbGC
nvnnTwJ0l8W0L9ps6ycGTTLsLYGIU0KZUpNGJUrYZnr2afL6tbAPXNDE91r/dJqwKrFKGDXTcxZO
VIv67WH+DGd7JIm25VdpDnxGSaPjHdrfi+P2/Zg/iVBkdktwxHAq06nIQjTz0WcUYGiacZmBeMvm
rvMLgeUHe9jJ6jcCTiMylmuUv2tmZmW7YZyCMEj1/UqGonR5j55lT+IXG/v7XToD1+lutWAlkWFy
eVXYduzTso7jrQz0WnXsb1ZRZWQ/S3ZRZte2rbkE1hypuDVY0Scfs0UsVcXZ/cjuamxTZ3ifcoLz
F5n0d5xoi84nW2hEh8Dw+Ye2RshT6aor4dDAGrOB4YqY190zUeyYJiOj6SLiTrPaUCPp7SQQ9YN8
xCgxdmLRKEduHv3mouKLqODmhBo/7khZqhGtRdCANSLyIb354qVpLRWvwJzLHtZilNEkFSqvB9XP
uCj36i3uvYqHBxspeaUwhn1BXnPdJVaBTE3YNELM+RTfu/GzD7jAFvs5HCt+SnKVQfD3pN70w3Dy
RAsJfamdBpEbLINz2B2q4Y+O83bMNK7mqg+F7H5y30VoPYngGx+JZk/jvH3kAR4B4NUfHswb3Vsc
VmT+SbzgWtvn+CKLGccEdf5ahTku7Ix9UTctCyHQdB9RsXqBASpxMsi4Qz0QCW879oSIvgaI5Jdw
PIrw9yB/mLjObn+V+J+xr3ue1H0XKNLI/7Wo5BbTyCmBlsisLI04nWddXK5fe5aQHScqSQY2+JaG
RsaVYpzy6MmarG76ZBG9fHgmUL1OyPzvefGOvGpxgyDh/Lp7Fu20RfHhjc4fjN2nV/Xzo0o0CgwB
g8p0Q1Kt+3SzwxG0iq9nkq3xJkKOghEQ3ZRcm5OjgonfqvNrONxn45TFUV9LxeRCVCsA1ed3fR8U
XtahKEuZ7gwAstlKhCheK2m9LbAZww0moI19Hwzbx3zxHP3TVgZ2GKvn22TO/ENmY1ELj5mZa1X0
3Tsim5Qzb6wYS1Z2KewT9c8fHELop3reZg7njrHPBT3Qp5u5Qlb35WHIsnZ0I8uOer8IC9GUdB4f
eJzFv0F5G0pNlRRBXz3hmkLlgnyFamMFEPobRB59sm3hBQiaYdUSP31r5RcPOzl0UkURAIUrQNVa
PGd/nxezVh0158wnGIQkuxJSa43SLpPfcBruo/Uf6+1nGO565q04jB+xyLBbW4ulARCtoGUfpeFa
6obqBF2d7xm3A5t+2L6ByBZUXMSBlZTi3yNdzgPbyA7zOSm8wwOKjmHIkKPUBDYUkGZrheuVk0wn
Jp4gJcMzg28OKzbRrpMfiFD6AcnRyMk8yZipTkaTBKjAP7tbjpzXY11aVLBLiIO/GTqVUDkTFuky
ghpY4og9jLPKCP3sIkjr/VpoSNtBQDEqGpk1xrGTz6UmDkd5Y7Ut8YUPA78XL3fGi16WzfcC6mne
zQFRzKBqJqsqIlPljWv/EGRfjXczI7D1ivTEbG4MZ+pldY7wMe2n0+YpVPRA5k3sH0Y9TP8HnjYs
t4cBNSgOm6sDnhVSz/eN5wCaI84CPjclhLZFcMH/3Kcjc6Xf4iWiR9hLhO5YzcuMmpBRypy8feax
lzb/BJxiXKOByiUZEuD6fCyGag4eycrl3lZHLt7GaEbB4LZofc9wWbvy4X6ntJI34YjIq6c3wJGW
nw8WbGlffmI8j80XBN6M0ReE9s360UX6U1xsEULl7kNgkPgnKqMkfOREzSdQO5JVdXreJiW+Z1en
rXHSRzYG+3zOKVSJ81iPJ0lFMpqj+aDYyZIcDczprUWsyLGn833OBwxpI0fXy5i4OjUTLpuG60ma
h/q70eymqXF5kajdkdDpqgU+I41b9gQkrTRIndzA4yQ2Sxn1WIRpwWAzqZHT7aDP6sMCVdkA4FC3
TsGCC42mevCbktUk4orI2du/Xu4kJVw8kW5X1pJlomNZrrrTbQZS/+Un/V1q/nBhaJH05hQ4QIpU
el91fdvPai9c4VaFWFPVHPUjqi9tPl/JWquitgc08itiEHjI3ZeMNEYYF7RHZFzrqc1lOz6ImL/V
SpDPqFK5wzvzQn2UpuDCK1FXnyOxc/kt8YBCHQxIhP8VJAFp8bTTZ8xX0ewD1HkWThMGWAJy6ZIA
/PMqS15BqWxuhq7f/wbevd+kdDSNWl0xbHqH8aUck7m0O56ssfo71qYuR9rOQYF/ZjQMoxP0KpVV
h6bf1PY4JleSfeYVcquPXa8trcx0VxOyf/NLpUtGGbLv07Ijf/nSSbEG3wBmq6modqelhvLOaFKv
AVaJ6eYkKCb3QGzAde/1Z25sRwsQAx9XC6wtYqjQkeCPWPwH8UQn9MfHl0lC6YCM6D8Jq6LprTRn
jKL3PiwHdUVTRnFOYShS7pGjaTw54btcxGDN9KmLPEiG1zWjTmRWbSE0ZTyjGeMdmywWoew8GfG2
bAUQyV76mn08GlnaW7752tIGZktJmho495QIT/hDO+nJYHnbU4W2zf/aGdmnxGYi7t3oT2T5Xm0S
svymqZw3rw7mSNWDA1PusculZ7y4FvPwShlkfckiNMIQZbp7Px6jjurZDlMd8bWIu5zEgY3DWbln
++FxWg4/coSCqIJp0ua2DKgRPpGRKgwFQ8wpKzPpn0bt0aPYi0iNJ563PKYXa4u/8yRip9Kmdpoi
vjeIZCnlMgIWGOmODL9dTwqyCNq9Rm54qOLIsdj8mheJCFqQ+HUlv2i4F2bBxawf6Tk8HaJ6AQKm
rBAGkpWZWd2QWoQ79KZ6luRsSsTA1UxZYc0C8f7jLC28lgYKTUM2K/w/lv/E4jvdA4y8ZT8ENhSl
o6NrXWnVsloieVVvWtYeToSfyQ7xNmvd2i64aUZP8YpG8iQLU7P6jcHTAfQdamjmU2PLjlLhB9Vm
+QXBbsZ6k4a1jPvBiIwz5ba0Axjj5NK9d1SEGs9zNoLsQ4jjKJUZjplZNjPEtmj7eQ6KSQk7IbSR
XyeE3WToc+cm3TXGQAnMKJvUtHOmj21dTDMnO0w/f/C08ifZ0xnry+JosdgBFhxtpO4hMCi8/rWX
xdA2+bEZaZo81QK25Q81fiWfAZJBTiLJKpnfKJnNfFXPKB6XFpa1tb+ZXE+mV7V/70cLiPB253zD
EUWc6SErLsDbEWsL0CPRUf0gO9QYPwYwgdukIC9xPKbpVUTlkekJ+lXDzxRtjCsIBGl6V2mS6rY2
n6jfKIv1dxDr9jS68AUchk5FWBKm2BAehMWP+MgY0E1oiMz9zk+siKkjt3PQAPgjiGH84O0fRXnQ
dsmjQ2d+8mao9j8FjCeswHPNKqkZIhxYFD3xx5jwQV9dd+6I4UHw8lNKIVMlavf8V4pwej2NhC4B
nNdb+L2V6w06Bx51oj3IWwhdL40+YbjMy2rCNt5tWidrLP560Y3B0vUliq5rrtyb62oelycTYoLr
8O84r6+qDSBu+c87eEe13eGLCEYBUbHar431UjZnUusmK2OHFZmh+vVnFnDubBoj+zc2qfTu8gCx
HmgGAU3SikOXqnl28yVqkJ5lL7SnWj2rBZoB0lJP4pIwZrrhrxad20otuQ5QR2Jox/Z6evRBM67h
BvfXuKc/CC37uqKdaa4N8Oc7KmWyjtNYheekCi5STansZcKq3oCXyuKFUIwOQyBf3CLE1iea04wr
VlrRUL+ymfCAmVL9ZJD86znXkhENbvn4BcmeCpyO6E1Vd0NUxOOadvUZ9A7/5KlNWrGjQ9XHMu3y
nOLN1Ty+8jsg9FablMfsEExO3941IXKDj2jmfxeomDVT4NstMQDLQmZTpstCbRB2RFEea0TTkXpD
Bbz1DmmVgi47ZKPLmnLlLJYK6nkfFNzms0nGp9nDshgu39MI5dg1WLQL9u3ElitB19He6Ows2y+v
5igJVm47VQqvqnfQBz3XvLBBXgnBsmqfd6L9ur5quvJdq14qDia74EY9WyR44YfFtVTSx7xILtga
q1oXz88Bj1bTDf1VWj6V+gYzDV2qxSwI/p+o2QrKV2oNHCkpBPoVrV70iN1eHc+dBQc1qze3RIE8
9A5Pb+9QFKgp3Iikv/ZgzaM34pc3cebEdM4b6014/vfiS+R8KFik4S/lynAbBRqCGn8GuBo/RDam
rC1STN/DFNdpptqrrjcDMr5ZlSd7oYXVEj81AoVMO5uMOGR/G3oURFa9la/HarQoP1xw7k+veJRZ
xjtKK+wgAU9Ou2iggmmp1YeLDXS+fJNbhDKSSlNsB+iSEtnVfL1wU1y/Odl0xg5ycN4XZc2NI42e
6PyWzWhKDvt3ZAfAZgIJOMy0jRcDy4sjZQMxA6020oimTZk1tTvNfeClB3MRsFGj5KRbFJE9uVST
/5ZtTuGPi559oAIh02Ns35NFJhZ3oY3LQZOZS4QGlrEvik0BvFCzFQ8S5B/+gI/LhtkKnaKseoQt
a00WZb5amGcB9FmUouxFgTXqN8Z3jop1dwDZUKafBD6h4sKzrjg3FWruXWbTmBF2A16tE5LK4K/K
+YH2MOkdyAMGS+dkLGFi+0r9nHBQl14hifkmypzHdPrPnW3bEbgqaDppJEYsBtMu4Gkmyhqhkmeu
WcoBEbwD25NyB0bpr0eXtrdDj+orEzRtC3u0UCzHA3f53X8SBHDbLjbXQnQ8IgZ0XZ/TinXzXuuP
kq/nMn+WgNw6Shd6zJgsrCg8u6XzMtz7Clm2kjVbE52wq1XzADhoPMy/r7czj4ZGPNT2jvf347O6
l07dJ/koCy0xcgAm/26Ul9BtWOkagIVTZFxqTrRsasCjyFOwinSxoixVDeJX1hKczPDrdEjd6L2X
B2TJ8cyvuAz0aojCOiiskmQqKKaZlx+hfYCAzn6HpPAP2hWM1HD4hr9o1oj8B70B8uVNTXgwxxZr
nMQLSUldIJasx2GOasohejthERNaFMfpIM7sjy4CSgSy1bTaQdnhcDTumMzbHdDPHYFSOniCy6PN
CX38Krfp3IaSgQCqNIr0rL3GCPED5iZJtYrprhI5PlEbm1/Es2HZfzt00y7P/Ox/KXUSHWf5oWRX
Ia30/LXPGp+W21E9wVX+9r4dA0PPg4dn/ArcTUsEvMDJKOI4P6IlAIXYhNWdx3KbTgT/Q+uoMAme
QLVF66hpL4e2Glnc/bTDcdxRIGA/232HFpsif4VBuHRnyG5YHizcdSdG+Z0XnPaD/VzhCjxhQ6Ee
/DKqslWHNkkKOe22XMAjOrVHN44U7+deAwO/GzsBvWwT07atiN+gAhwxZN8XxddniUPLsPOE7uI+
eAZ9sluJZ0TSs+E0A+18jiwdNlGOoK0gu+gVzji3f0R7aT9eV1UrfMlrXJILKYdLaQ+gfFhaQIzM
deYS+QlFa5GMVblmPIL1VjytnVJ2aw+33A72/a6VR4ww5IbO2QgnFz5GZ163JhAV6zvNhxPSJgvN
MxJ2Y84o2GUoeDhdhX2kIEl7HlIJNB5WPoeE7813ael5qvhQ+vC6ZD10fy6Klh0X9RzHn2pJjFcB
sKWCEHf1GkAz6/TA8FsQCrwVlMxvS25FIFoRDOD8nw0XuYMXRCDJ2aydFJIXNcozGgkQELtxyKIV
CaR/xJTe2q0Lm8neEN0jwkHwDoubBRE0Mh849b/lmdDiqdm7tY3W0CmfG2YtagZ35V4iT3TO/NYr
0vXcHqdEH7Uni5qe4G3q/UgdCbLX/rUoDTcZmcz0oXq46uTazyBRxRXDKu8J1Du4E/+NxNmR18tj
1a7/YdgTKIeTnZmjEVKfHEWJ3yp5GXQnXtfUgK/4AmB/jubF1Ec3YIGBf9KyMZFrPhBd3dN5DnpQ
vnpsnKue1uFhpt2ojkKKHNB5APBa583A28N7yLnk7mHHuqHP7P3R2bPVB/92TBa2jHJgJRe721xh
2ghiGKk0fXCwua0SesfyrZijlWLVgagh19Ss26YzQEgpFUUimutBCs9u/7tvu3zSJowloTje6Xo8
Qlbm/iySDIfY90xvOP5TQpIDqO5uqwa2RYo9+kl86I9HtfvCGwn/9Pc43qcd4jLw1Boo/ZXBwsyw
BCJhsuc55ikYLGLqF+4nDTJZiDqj5uIjMsVvnSxaFpPgYgXDLA/KTpd6qyGMuVkAB1Bu/1wuubXb
42KRrAFF8EvrKChDdr9tersic8yIq4BK/cN5km5qbnNobS638GhyVH6dn6d344utHGqCatL1CLSs
gGOFqCj53COvqUCegKQlQrdsXw20Bjbnka1h/JkMJO5FlfadeUiswLa18CJDjyEYQ4AgC9xU7VTx
6S4WhpaktRhjrOIK9BLV2nxGEQkTxu0bFdaVcqDXDgx6cPtueH7lXzGpVNcCOk2qDNOA+lprbuQC
o6RN0kMTDitF+4XECre7nzbGiR9/WumLjj+Q91WlZePpkqX7cDXWfmiNVH/wqjU+9vyeW07zY3q7
QkqM+AmCJbiN9opCHfqOPPGH+a7Zjav7K2ObIRWRanBWXF0827yX2p9SyTSwwwx5O7s6YVSK/F8k
m7t4bX+IwosafNj5rBVLvqvEp2vVhWmrfiNYSPLiAyY1SeP1XC8a5nwxGoXPxy2+ZgHuq3wJZHvg
p5O3aGZfPJgFtWdc2RyFJrXvxr/iYM8A0mSiNZgZs5X1LIcOXoXQJelo8xhJv4e3PBQxC6ycwmda
ZBt6oGjBESipwI+jSgnHWYZywbKg7Nx1CRcdQ6v4SIRNDqR4iqtqKdQwgh2uoaofIDaHAbKByf4s
pPoTEf7AhogjT+bIzAa/EGHGvFpMr09vgCLRD5DZkilZy0bT67bi2kdT4UfJC0ca2kPMtUGjoGXT
EfVw4bRYKfKH2Hb9mgQazK75gfO6Hzo0AWuoESjr5v06u52R/SJeazWOisr+mLIG2eLTaaosrhGE
Jx0YHpj5q0gi5N48vD2//upeG/xQqiVZRXV/DyOHc8OkIFAlf+frnv0HkhMXiwNWKJtFInn+3lZT
L0XImas60d5AVCQxBLA2HPPp5s9yr1MwUpgPy+sYiTYJxSsvQtQ376S2lrFumtXhD/ToGil9KB/u
+r1fAHjxTlsuPoL7WBTYu/mCfsOHm8YEZfBO72FukXAZFaVX9iPsHZ0tEPClJwa933Tv3+TwE3Uf
2gkEInKVcwrpNVxYK2AjgNq8TkA9YJ20kobebbpMVx7dBweVcoK2tH5F+Qg795miW7m3WZwk9LMX
tXlVFr7gkXWZ0iMCw2k7s8o6C6Q6YBDm7200uWt8W+rsLQp503DeM6wVZ2a5KlhEPpOifdVFNVDH
d7kJQye9vn0PyZ7v/yr6jXys/eAnaXrMvCNuqHfTREqJ3Nke/CjfV5Az64Ci8R8NkJEd6A7agXWM
8ozZogIXHwgcDVJBB+3Q2oMXd+miB7K2/HEuqZjWV098K41B9pSFbCTl79tQGpIRLGsT0zORaTgN
rVcyLdRPqdJfE68i2DM0wLdjnpYryJQ3f6SdsuymJMRdEkUsN0ZNx0ndWDZn58sdnJJty6lLZNP2
+n43kW+iJHkNhIV/2tJYNBfsDWihUynt9z6vZ6FeDs617OOk5biIBKHq7dp2FAWP1MNXvCYZZTXe
en9+E+OSZVvEivO56Gn5M7J98Cmw+1DQlROfzEbpvc7pPXZP7HQvPhLHfACy7C45Bp7V83OlwRwR
HHQzdcdZwiUZSBWqSog/elcV2oHq/AtXI5uXqH2IZB+n1dR21WSvjQy/MiI4ayeKvcfWeGDUn3h+
B0l8DGMX7TwYcBQosKAZjMRFkMMtswA7jkfafbr3wN2QdaaioQbvDFyVbC5fFRl8ShG8kL7ggqZ+
Vyor8nyoPc9EXDH+UZrCW9Tb8wVmngfUSzl8T0kEjuZ4lMSWYrnbNNamnQ6YB0+zslto3f28aPzD
WyQfNnZfIe3Z21D9tvQzSQ7YXDy9GfWGKHTDkUylPOhK4QX8RV9gUAfXcln9eW4H5UhLbJtOos1P
ajpjqTnc3D1VsHsW59GAQUx1frr+oN9MyX9gm/V/7sBQgVaGiQuVZT7lgmjbAIEM8t3nzKN2yBf1
G5WPJs+4hQ2Os9XyB/tmE1jV1khp4YkGjDTSqq4/HImDzA/w7oScBnWZBOzJfl+TcY7h4N4C3m2p
NZS4Hcp0ISBHwX9K/rrypxf7+3IyZ6HAtf1bqvPy8vL8IzJv32BJ82OhE59s0THdrcmr7kacZPAN
cJRwkaESthjCOQexBGmjHRLE0HlpKthd7c6zjI5XoCh7R7AoiPjjGe5ssoNM/uIGz20nu6gaw8qE
w/DqVulW4KK2r3uKe0Gt05ZkN9mLg0GTFxoRKghslE/EOdMhIOKd85xTTkzbXU1mYbCQqe4OUI8b
0uoCxztTUSt4kz/J+pIRBDh1olFlrluyoBtLqmt6G/QBl8UweG/iirTqHW7HxlXg4nL5KlwLwluP
XmasFoku7528ZUCCtNY2E4T5wcjs6Q7tfVM+SunNXXkl7ENv4kTooZcJZhw27R7R62nWAaWHUsrf
8ftae5KVc1U/l3KN6b3OGofVhhFQXNdOhVFBTTtR161CfqduKLLtGVl2WUuRQ+BUaTz35HIV39DP
kbrjyPC20p6U+OQxiCRxjJthZgJ5fAcqnVH72PcdjQ3M2pULI8FVfM4Vl8i5B/aEMj5UzSt+3bP2
RCB5MkTvkHfpD/60MNnGxaBUhayehOZBu6goG94ePVtDsAm576lj7PhDryik2+fUv8wBp+CTWuHb
CkYcR1CWJ98i3y37wZ7COvdLrJ/INRwewl21j8d1gEBSPcMafkg70enkL51fqmAKdcdDW3blHu55
26oyf47FFjP+3QdKDCKrHcsVLuOiHhnODQlp8JBiOJauoUQRjZIdMEcujMn11eRHldLid2H4kBU6
MsoyZyrVqcV5cRMwk63+fwY1yjacXVoDuouy9H/Ypze0DFr+C6wKYpHvXmwouGgNFUDNUamD3pLn
9ZM9JXInJH0BlNu4LNArgAT7dxekwTUMSg4mqFQ+ufZCuffWf2L9RpLfQTRGzsRdNgHQRvy7Dazk
Sb8qfbUCrfEfo/vOA0A6+inFieocpuk/L3wUWCVgJ+UMyCm3/8ye0Ol9e7/uFIJKmR+O7wNMndvj
BCkQ4XI19nxKQnpgfjeVZVSfBaoUOm04L9lp6VBtkMVCCN7GfBYYFKq7jsZU5f8GFZ57unlIOEHg
ePSit9MS0ZwkEzMc2TraH0Uqc/z16gRPBTdmYioh0LQR71BIy74ySPEtyCFdnCXCrGmQgV6l7RqX
+GBiLMvLe0ngRoCtzuotzA5/zZJvAJzPObsze2d9iP4KoSCHGKFjyPxZJqCc/ZQwpEYJJDYVvmnX
0uSGG1HoFXbquGQQjUga2y5wTT7IxUgJBF/Nwhx+zlgc5BXk2V28Na0xRouAlLqKrr1GA2vZ91np
6XPIso+ulCSSR9HPuk1oQ4ANQof9QbSKejq1nNg3AdHrPDlE8JU+zBE5bmVgflGMh87pTl4wdway
taX6hfCtDdgWiGoYnmdPDYdOcOzAF2GqnyzwYqDR6n7lNPLbZkQZnWaMjRPoiV/IZTGxHbKWRoPw
1W074s9iPMHUQCyFEgqRTaNeE3bNesRblcyY1af7uKl2UWG6cZ96/WWVkEGSeIkCs1QfNoZTY83g
Wg6CqmEnyibs0OOnJ1MYoI2Gd7zpDiewP0+0TXmbTLeL6IFuXcf9DaLqw4FmNw0tt5zsytgfQwZd
GRYr0Cumk2no9HftkH2IsI+MIYWnkqPCWoAGb+66unq+L4uXjgQN+9h0dy3mkvL0aprS4rNFRtrC
28jU8RKYukKXZB65Vv55Wuc6ZeyJ9jz54LVw7LsxgYFwnVA4Bn5vTaXNwWHDF08reH9M6jax4BPy
X7hyRvy7Pg5dbzgqf6qiVdH5jRc9LNMctQDESMCNbN1dNxiWVKFECkvN8NSuoI+jauN4i8MykDbH
OI4ROa1BXgVhesd44MseLg0bpITxDM7Cgjvy+kp+MUM1NxQg4vFNIy9zr8wgFBGi9h8ILzV5P+1A
+kGCvklqnJlSyHxQy2GI6upiJ8tDpdW8QttW+Zq/TcktrQjFV4PEbSPYN1Tv3tBqyXgisUnLbYeh
4SpFVZ12MzZ8qudkr96sJm3Jd0qNxKcYRBXccybK3yVMUXujwQoXwr7XNy0gKjMdHxHfLrR5kiOd
1CL9rdvFXj84W64/Os2Zs1P7SQc7L3t3n2NH6loMvYbfJy2alc2T7oYPrzsFIMGZuuRPCZ/01pxr
3uOGy/JBNAlAKXDjuWL5+TdSZJe+T+e30yqjUxeI7bLQp6IKAVdJVUfm4EgT0SkF72qSeYp9NfPy
kzhABVT7OwadHCDNuA4mUvUGunWfwuEg14T13zqF/m1VCKjnLLAYrSBoG1swlqrAW3MnFxrcKoG6
1ueBYMWTgT+I0MUqFu1Up7KuQTH0qg2SH41QlRlupH+rFn7BtQMemFaHSD63AsfHdlhLCubrjU94
ADgMsW34Z8R9LN1HPy6IhQIM0qawvsvPKVIz/ARRVDWsnCMXU8R5Z1XriNqpXxYbcxgSBG41AspH
rRYoYCKRGvjDNjv+j+N5sUC+UDJRkIkTXuqSqKWXZ4rshEuLN264tKwNS9EGELapVHleiUEqWIWQ
CVKCofOmrJXT6odeUsA9jk7P6bDMqoHCX/uyRf/zBngDHQ7rh3925gZ0g1I8EUbbvPssZVFslKtP
uKR1MlhHH3FEsCTSyjue9zFBAKOUTjN4h6NbuMdO63CluIz5lomiUCHbz8zTzApASNMk4hYXGwN5
qO7lsQabrqLb1GPQ5vPj+KqzamnNDuaQagGsUqq0t7wQhPVvGw0aGJ6XjlnakNxwFi9F9b9dnqZa
ncoh0RuyQtPEdCgVNcwtKsWXK3znlb0xxhwOT3DLk7cb2KWTAeqWGNlPuUjORF0nzvld7q+h2g7H
CnrAOlE5ewrK3Rv6qWhFm4VCtiN702DV6C1ob6Hr0aozCNRvw7SDGvxOVVu5ENElUx6dUQQ72thx
weJScLK+PbhpPUDKW+cWHW2xhfQOWekFTU4xP7WzlDv5GQwMTeDhWAlWSezYYq4KQMFoy8jYPOXZ
12gYT7WY0oW0AC+UhYGYhg7Ntz35xFsqorqDA04gg7rCXvpAx+QvtywdXDimjBqJ9GIi3wKO3UjU
hGMcLrMHfQphiWwmk+0fin0a4922jUMk4TzZEsomd62HKegTxbo9FVf6YRzHpexw6Y2XwxRzMJ9c
FcBKlGsSeiXXvCPGmFEKkuOWRPhVfzrgpMHChp2vU/IB9L+mf3Fjlj0N2Jj5ikY99WSa56iHwfy/
r3zd0HgQwoIqqxk+k55NGDWE/Gnfjkz8kufjnLhyrvvc6IX3nb51+Ay1PbMzqhlJ4uExJZDCStLn
CUdFw55PUTlcacLaMQoH1jWk2V/qqBInUIVDY+t3WpcHmB4UcIVIzwTEEB0rNR7GZjT+4DMDAXGk
4701yHGHeFYk2PyEAiramToLVIOs5ZDRcf51Yk5Yjbts0tTqE7u5E2yLRPzsr8nu2GV9Sp0Jrqg8
j6UysJwpJb/1ZRA2k5Z1c5afcdNuPK73NwQrhtbcAhXiMW0cDcJ7FvgGDVetck/vimbmnRU6nyRl
TqRK+OvmgWkL93wnIB7LCvz54wkATJTNXjs8HsCx2nIUPbOd1DU5If2os3yzt5meA7N4wK9AKZ4j
+HRUuHPA1Fk92Mgv49Oow/JVMg9ytaOJhFSJLuiXSAov5EJy3dFx51Aem5dPKbDTmGGv9ZDR2Xe3
9TI8G2A0z+NjhsLdDg8XUuklj1Wcajv45qwo7soVE4+gDzjjzLqqmtk2d4MmPKPQ95mNr1VY+QWe
RaN3Q0wZ4STveCHgsf1cqixoxmhycrZ07AwZH5bNOlUHa2Ima44WF430KveclH4UwkBE9j806L6M
1jb/B6CdwW3+UOlhbUKLQ2NBzv2J7RAU/SYPnrUT5lWdD/JMea/9qEhttZrvctvp/EVqQ7qdLH++
x25UzN9HN8F2ytgg47qoQB5OI40StvkXnT4yCEMa2EcKfNSEmhPZMbgR4UTc6A9H+oqpZEa4Vna4
wJph+/8VX/xlRjFWR0M4D7UZtq6+irnQmJeIQt0gxmRlAEt06TkPj8f+hmvb+Q2kDrEP5ufshp0+
KrYgwsWgl9GPUfek5g+Mxonb8H6Q4D34lL5S/8T+GIhNPYsNGHdzFho89uTRtZOcQL/mHyOAA4cE
z+e+HBLSKZNJeEb0eUrcv2/ITGv7OgVwWgMyTNqDOOMv6qgbi0DcLrbKGLtAD3EdgcNMSbtG3Kvu
hbD7LFbFJ49hxNNHHo0GzVtNk0X9TYHUbU08cipsD3xn6UIQgVKpQXgmQXaXJlmhUdyAwx9flCqu
8uk2iuih+66Gl5JtJOcBpy3OFoAFZWBYLBF6gO8bkQjVJaP0eeTCJigB5MmDX7EIb2NOW4F3K1oG
GUmYPyvkHHc2/3FIb+zyPJWO6tw+f+IzTnA9cB9OesLu9ja+OQOS7xdYsLnzr9Cz+upNbzIkH68U
xDFw9zpM9HmlaXOTNOg7CMeexwx2r1X/cBQB6VS3He1o6RzB/oPvHchis1Ogca2hlLgpPjm2nacz
Z0Vsw8DQxao4vZgzxmLJWdDebsM5pjOS2u2NGN4jXdEW8Sxz/1ViIR8Gp0PjgDUSIB7W497KzlAB
QIANqzMv6l5RZnHdGyfFihp6Tg6WvfkEEhTYfMdqLwltHdlqw67amQOz2O0gLfO32pvJIHF1AqXB
w8T7xBIewAbgIbQQ6J1o/soiNLF3BuvY1y9WzSEY9mC5somvfQxCMpVzUaPLnDwqDKNwnEGEYPB+
E96gezeXzLoyKKvFlT7h89B4HWMDP0SIZjXWiniONP7CjpayYcMAdENt5RJqA7omn2cz7PWwPCVe
mPguVsCIGs9wJ9Q9xEpKzwXtgG1DRF958kzFHpl0r6hWQHQewpI14d+8J/LT5wa1ADKIIwIWju32
c43C8/aI1L/Ngo7mVRHAzLAwEzkpLz1K0BM7ACQPSoaJLxzs36Ij6s709td7Af3UZTUzaT29l8kP
qDkFie0AntB0LQmV219q6YVvbzmhVxWUIZyQ/pUjRAAQ+VR/+8D1/HuRULJaUYwZsUqpFbwZkYGN
IalJ3j33/lRTTKN8kbFCO/thmbdytjaDZEEBeUWoVHMMpRc0nxLHN+D5eC6HetERXrrR10JcFkKx
C0pSku/WuAaXg43D7ZP0a9kJaplOJNyLoCK0RUNJusno4L8d2z76fOzJ3JykfaOX/tIVp6pG3jdo
x2m/nVjj1DhgEeCP+qCxjGvjIA8ExYusw5N2EqqQnrUtll/wdrR9Pr4MYFvfAHNXp8owg1Mf/QsY
Th8JE+M0CxWSdcsCOIQerMH8ChfpHXvaYh593pxk0LVZSiDVaQnCbossbqWP7KPf1JwMXWRnxiqo
OoFdNSfW/GA3gpPi7Tiv7jzhb/q7+zwRECDkAQfwEI+cS+g05gIw1DzPuUD6HgRdPkAbawGnEuIV
ZAZPd0rA7oqNPAKd/u0UgYm3P6f5AmRryEF1suZp/HW3SOfAO08qGYVlSlmguwJy57y6Ay6BSSbm
DVhO403Ls5fCuSOLVDGEUpy3d1Oz8PZQ/A0OIAWLbqc9erfRk28dl9voFMRmcwWESOkPs3LrxcxD
y6wm5hnzo/n2pnwdGZhukeDJ8n/FKA43R89QxcipOoKuI0/ZMDeTvap0WYYYdcp7ottIh/mts2+l
KPEvNJzyEkTV5uXgWjum05eCjrlFCuxUCTKQFjdFUmE1F8Vy133zUGCnQyZmot65lXX1OBOBJVDY
O8QCtjU3m03dZkKgpt7qLqU9Qc/ZlTfaobHN/szh+cAE045Mx5c809ouAEdAugyO+dPhWyg4jsyI
okTvjspvYChuJMkomfM7ETH5xdk1x8O55eaddVYln+VcZno2m/oqaDi6W2MUUYrf3JdC8yoIy5Ds
JvIr6QSU9VK5lPwR4jakeNIFGTz9V89qRdTD2onhkPpfXBBuyLvkcDiUnl+zQarw4A5ZJZKW1+dA
laylcdBaK5KlMsrlSMNclmq/lcsPlXVC3bM86RSF21D3HVlD/QBpq24ThOJBFP1u9WvgRLCOWKx5
voZQVmYFBp5hLVd6V2/CCr2QHHWvi2tSSJmjoLfTiQDZ+xusbIl26b5KYfFapngwcMKGInzllz4w
NQY7SM1GoyGuDaRcyGYyVRahqbdk4q1Gf2MuHn7jG5G/a0P1BZ6cORcmx4haX89pfkfj2ZsetJ5O
AA2o5CxqgFF6S8IcBUMhj36mzv+so2zEgWYGvsqxnkICJAmdeo7g3dwWf55KGFsKcmQsRsYYcPRG
k+zz3rC2WtTkDSCyiRK1m1h4GXfJGkxg32bDzRNNVQ8ucXWwKz2pjybyvNzchr4TdebPXFFhYe9I
0Ja2cOrVGGedLQn0BwkNLX8/Z50athvThsv4BrZy3hvBM/0JZFy2PAwfeMlJ7erqmsiWP6KKxjn7
fKsG2aW5UGCoAliDn+cMENqfnu/ng3Q3SQB43Dw0Wn+8y5Wv8E8mAcRUM7CNUIN+WA48rrOEf+yG
J15RN4vr/dwCZ34UEciGn6sAVEbI+aTNh2oID309WMNo0qf2QIJI50VMvP85TCNTBoTybGtgKmCJ
wbrYZqkvC6vLLGcGr//Hj4vbrkzRDifZclHnsjsYokoz8zz1lWUJwEt5PqAzrEgg4qmxieNsEazs
9EWaVzP4i5M9HZnjErbeRCA3PWcRRINrX7ebGkP+D7f4oGlB6DcOEV3pS7WFlT5Hnhp0NoSNiUlh
wRSVxMua0cXUicb4BwWx4bZnCZz4MoBrfLzPoc0GLcCSYA2evEVcgRRGe8nrFTobrYwd97UEtGfm
50ZEA86mz2WWqCTr6T5xCtX2KwSSXGcM360iAATc6+WfQe7Wu40qo+XDkbPRFhVDVfC3dpcGMqj8
VyqB2mBhKX2J3d25mSh4qgCiZ3hk5AEUCYFN3lnCGmaldcOHnW3e8Msak6MYMw9L7No24l30iCrT
Z40km5WeTLzLFHr0VgUAn6lTdY5bI4z6hw8dp0glpp6pI4+N8/Vr2pL38JPRMmUf+HoVVg3j3hEA
eaCL0olJGf5QQf4xeUSzSR2/uJBZ1hlfOvyElA4lEc8wb8pwJAWrHXSGnAzO9jtDlgTnGKrQuoSH
Mp5WXcTXGXr3VZoj4Q2ucL0c59wPIr1O5dlYs2s+8VISjWmCGRDv5yckcCXjG21mX50uv4xV7iEd
5GY2y88keO0iEuxBSl8bGdjWcIdFHq3aakYPYB/FmZgxdxEHG8bKP2aTywpcgH+9IzIe07Yf3mle
T4OcDwPwudFqXvl86fKMU+4pwdgeiNDQl/OwLRjs8KjLj4RIc38Dkw5mP9C2k2g1anKxYLLKeIkv
5mCb3I4F483kPge4jkinWAT/2XxYoBEpFzdPqVz1t/qyDeqdnLJBuelukXVqRrm3IhO6XlY7ABzR
8kaMgwtiybjerZtHIFyJNQLbx6w8eI41u8+mVFYdzhZc8zO/L8jV/Q02w3cPJtfno+o4U8Xr3mD1
9l/Q5zlkRuqtM891ghExM4tUmtd1fI/QzPf5zDLC5b8SrXWHPD48Mh3Xyb7Jnu7t7BPmieYc3WQK
c2J5j4BxK+oxuRs6V5XtLILkRxH4dkv/2PidIkQZAyV79G8ZJwIRSRgDdigomw5gRtjwIjfExQqX
8a8yGMU3jyHij3leuSu9fuwm36oOM/1r1tzd69ECirlLIa2CHSj1JVDjqK72bKz7hceXmpA308O9
Nvu+6CQ9xg7lieXMJ8tcHxfnbwNeXHXz3rxsqcbxoDLY7FIZQnhEvHKGAyWM7NG3DF6zOISn56f5
ItwZVQ29D/4P2p52UP3fMWzJQmDXT9ZyRbbzfINWmwmgnjkglOy8TvGiHPN0/lR4rQfR6aZP4kx4
hs3qCzhZemjR0FrC6GGP7eup70t/TEtsFbD4kqaMaWKQuXpUCqTo77M1HoWsBImdhAxfANXpBI7d
PKbennH9OCCuINKDgr9BSQhac2IO86k0hp7wWVqmEHxK3gHubRPlnN1UrMHyyfkjdbthe5dhl1hm
mFR2C3ACIksk/xRn78c9nz65057FlKs7SdV0OkQ9sQftqz6IOYQtdZ87acdL5N7Zd/e4m3MdTmDH
e20af2MGp3DkQtqv5hf9XqhtiMzdiFHx1SR3Mj7IaUt7D4KNyqvS77jPm8vkjEZJXW2tUHjiBUNs
PMwgcog0VLvynA8PNlRh8s5DzvSf4PmDDWm//DfiJgJGXhlgdC9Ur7hFKkyYJ+7WgcTHQNomZINV
6b3uRE47SgqrfcCDaL4EG4HcKrNoEXvLA9tukrlZYX5feQle22810bIvcP4Nk6zQ0wIfU6vVtjQ8
9KFbKlPIVAnxijHoHEp9cX9S4yVrmbyJVOKoRCOi/79dKM2OLVlIMzGmQjgYLiAkJ2b+yLheJumH
7QHXcMEaGVorrKUb0p66Z8jcE/kSLr4Zkb6siuLynkM5A7xEl7UjU2qL44ZWJm11QCWAUU7eOF2K
wfu5B4emdmv7OueTYmBQbjhp07yKmFWeYJ9w3sUpKhAYcrXgjD+8tk9CR9GKf+CeBrEFflFOcdbF
r+8SZNLZewft/Dsg8wvV8byqzVUQAvU1NfKE0gOKb0mehkiBFCde2SfuRpFPWuqGz2WOzVncDJXi
2dIuoLSEYYqQ+KsFs0mXMU1Y+5THp88MKuV0W4McnS5iIPqVtkPVkeFCjUdHttvaxoGEAShWRWTl
3DaFB8PonBHDpmc8Uec4BDLf0sxjQtXOr7oHsRrzngVhXKYeUGnvZo5AvfXIXwku6Eykm0gbg7Mg
RXL/ivrLryJeVNH9G5QOpiUJiIlXKz6IJs8ezChiausNq22rCX79RVoZ1R+Tf5idgjmEUCoSOEH+
Pp6Y3k0v+Vd8wGQa92UDD2pw8T+ZUGTZNJ1ofhdJtzJKZ+h1Vk9FCzy4xTP+tSPDdpxEQXg9uSm0
A8dQGrDGR9+7dy3aPI3M7qLgbMN0alMqjO3nCZ09YalrAwRXP4QDdjn2rx8sTmyVUacwE9vpc8tB
YLKTAqB9/W8otoTPiu+Ra9Gl2IaL4uu+lzY3GMvaAvS80j5KurjP8kt3jR1QtvH3FoL51pZN1tYR
RfqJOTCJydQNz2kgFlbqWhsbwBTLAhX3FN5Um+AWx2QdhRu4Rxptct8YLnYOWWIy/h0+d5uzr3kt
imnEZs7wGILs9LGbsL3JOaADZDht4N/VUKqzHf//XpashfP9a7Stw+LNbcCdEc6VcdggC/1NT/W8
pf5T9mOTb9bHXNrF9bE1C9sDPgNKIQcEphy8Ghfjuq+oYt2AliiC80e/XPwUvxiLLF6KQ1xee6ax
Aj2izbgu3OW5xfCZNeXPH75a7iT3gCW1i5G9otDMk7pTBp0yEcELcP4qsYDU0/jnqgdGPJnlH00G
bk5l4d25Lv3+oeEylSanUOAWDnUcQ0broVIoCwRbyqNhIMG9NZSaTwqeYIUmHtTaeJket8qRuax6
W6vbOMpHORVwse1ohPIb+8iuqfIHGNgNYxA1MkDqk0WmcEja7doV8HPIeqcZ0M7HTcW3VEPx+sza
PZ4e/bMUQ50lcQOhw17XRvyifycS7hqwh6m1l0Tv97wzzU1/UTVdY89+FdKe5Qi+hqfH33tXGcJC
2wOez6uN917A6T/+hA1KGaf4dw0ZDnTw0taizezI9G9Jri1X3IWnIwW9N+MSdXb+stpyuHS3MvaK
e8aUMJUNvo2Y4csBSYQNIJPfCArI+9sN0J0XVBmV5UX4U5RwOnTgJz16GaFVGQnRTbun9VrBV+Kj
J2t0LwLd4vTk/MJCDukf1Y/0HoAPYryCFqR4kqyAtbfvdwEYRc0C4wuCh79tkIe0QMtcC/ZA95X6
ud530JlVrJbofE2fzWOe3juF/ecMbPbIgfC8a1zpHBMgMiODkwJFiHsRind7CO6pfsMvFbcn3DPP
F3TkR9oE8TqjF3jZ8o8ijy4zB1ptoEV9QwYeJLjY0kV0TSikDz3dPGktl8nZXFSOMydlHN9GdQok
op/kb8L9EBeZnBVHylNZ6+CW2iqVVvfEz63t94OXBD+O6mo/XN4vfBhoYD15njdSrfJKn1hw1PxC
ortUnc4HBfpWbdeafRWpndYHR9TxS2imLmvU6oPMgvNT9Gxtur/f3kMxS3VcUyvAel+cGXR2coca
2aprGl+xTnl2neaBwIhzM3kYUPFrdV6/gLKBJJEyKRKAxmbIOUJe7I188r+3EXLxj2OUv1JmZce7
CTkDTJVNKXY9NgYvW8wV036hAhQaI7FuJLlOWBPYuR+wQmGeVvuz9WxuiXk2t3ZWdmR7D46ResOe
A94qoP4wJ1Spz8SfFE5wUuRwhyuzlzTRMAnuFagB2Z2MJ47svJw57m3NvFeH/bhyvajVYIZWU/go
6bBA4knlNCg46h2lpRut5lPq2k+2xCSdxBS3Se2J6xNYod1cpmRJbqga9NPYXC1i4AxVnelnWxf/
PUvOB6wF7uxDlnpNbaBEWys9UdjPXiImPdRCu56yyi6S7hg2wBwuiJcr7XXdygNrF69Wnl2TMfhZ
SrSzSVpPW4GCFwDQY9yE1sZkXew9r6ODWKzWMahjE4MhW2yPKIJyp8wRySFISBt13aYZYhJM1igO
Fx3jU2kNtfpzV6QK6mOyun9UavACFhpko2Jw4q86aoxU78cYMlwC2SvDRN8rW0c3+YoNFKL10Rcr
Qa2IDfRIHHwiKR8oLcUyLawWcqm6kSx15kJsocz9XATRv2OhLm8qBdc37kauoBJq2wMaMkcOBq93
ucy9UP1Y8gYnIIJZLrNroFD7Rx3LEBoMel8PEJvA+Z7sDZ0WoYKtrQoJPCav3XY6bUIXoiYE7FkV
IouwYlDrINaXvObU6Wb3MkLlJV1Lpf25lP1JLPDeMv8+m5gly3F++TIkyROdK4cAdUhCMdY9Urn7
kuXmU9aOfuxQk3nygBORCZvL0RXt1DQlLAYEKegK57uyr8HfUWg7fH2tNnkUj30VRE2OMNHlPVn3
1zkYdxHT9YwJj8GV7gMCBnTDEtEqKgfZP8Ica/x1uKqgE5eI0sb01VtAvqJSraz4xHW9BcoVd8zH
yq+z1tAk0HcXnDwoBZzLkiXmuoYI6EzXiLGSKNGzHuMJfEUUtI2tu/tMMcfXTIfMr9pAbxQ9rS2m
78TUM8+BnYct3zuSTv/E/4sqMo0aODDdhURoN+yj98hODqig9AXGSeBN76LOYU48N9WMqSEU8al+
vgCn/8+6k20PeZYJOxpOL1U+QemfI/6nacC0g3WHDmjZvGhF0ZsIr/Uv1w75QYInr3m2OM2V+x1s
fBtX9RZTTZBX2BqsmP/ljgxXv/ntxGjZAKYFJYIDdNsto+yMsqWVna8OmBVkLpHCY6gu7/RZebRe
FgXc73zszNCdb8Cjzq/Ax+l0aSa07gDElQU6JyMoj26HQk7dNT12LIhzh9Z3kHAyrjeQNQaaR0iH
WforhmDKyR4sljqD1MzNiWhvda2QP7ORugpQbwBXPD36AcTidLe4ACwvnvALEQck9CbFC9s5v2eK
BbpLZ52J5vcKAHb7ixk1Sm0inLf4f7LLHBbknoaJKNP6eTZUbkZrcLbZrCd5j0eAjJTjtMTHhIgq
QraZ8TQYLKOvDGEGJU1urUsKAJOfexx/p7H1SsVZOMZ/vOnovz3fSVZz0s9sCLMi2nBPmcIMPwLg
fnFAbS2+llPYw49dkdNihQnlUYTv9Sc3mDaVoj+q89kiQOvD+Q9bocb+uaz+VbDx3xT+qbYBIkKt
vmC2aoR6PCF+fw5DukwO1QKcssvCn34o4rL45ow6KxmXncFX12UnA87LvcFMoTZK19PBp2Ps0CF+
jrh0bgntJ8pw68Ej9zrLMzu8/rfDO0ZsbBRel7Koz5GEoVjixj4P3NzPIuBo1chdU2RDLi+CzdWi
niQlZOhkzA1JoszcsgNaJrRl/TxCY+h7YAtkN5FJydHbPz+551wCAEzHUvEOnsmR6E7uWomVglDl
T/cHUTXgdxUcfLODDGR6wlhkFwsMIOzlWHHdSGUEMXCmLr10qUlVXW6IuoFWajTroFFVVfjvd1ts
Xg2GpNmX2trPMJZE8xE5IoXJ9YR254aaIyIkYDx8A7wqGPoAOORqSpqAWv6hMezZf4giBzjUNZKe
7V2gztrTxcCVLHj7TBYA3PwnSISnn1hAKLLvn0K3Glgn+SNFLD0yezp3xiVTh9ike2dKXoscfOug
kJ0htECl1PMCHX5/nvGJT42plgDTIzY04mxmmyvfsWaVvj7Ntg64HOQtmB8zMbnA1KQJ6BbxLd8p
yJIqQWRhELG9QttnjxmBQB36lcw0Lo+F1W75jfWL86yV+X+FffI5/RAnlMLdk+fR+HGd1BU9rynN
Riv4mWLys8eRMqiHcUwCsYwGTfHyXN61dgDkd+5JzQHVAhLl5whBhZZQwXX4tCB3NJOqgqJONt4Q
rOBdyab0GCRbHuLJlS/Do+qaOL34Bk8C8H1ZL69eEEmYxW6saLd5ZAOKXqCNiQ17LhV1JBEETBqs
0O9pilJWktna0WR9Af/DeSBWAuNzCRjTVRwrGHSIHvgdF7OATWydzZDDsMihTIpMLZ83B6uR5As/
lW6Dj2RxuDuufj2LfxJ8er/7I6Jn4dc9z5zaKTCYvWcpCF8CRdfkFB7fRp40IqiO330Dherse0YD
tIEVtV+VcApMsET6mYi3HPI3s57UcOeaOo9ACNVsY3AKtP2lrnJWQCwakP7a4tl8xYjQLP771Fs/
zp7aW65ToHFrHznuLToI6+zUtL5WycMFOwz1j3jluztvrflnfKgFl0jKb0vD+mUjTV90VGfYVuFL
dOitqSgicc9lseG6KeuPTxEetTZpraGkFfRKk6L8OGqBJjRjpNUF5FAoQuGZgbK5T8z3xxK2C0Be
7iW+AUHkEdmt2YWmaGdNnugJ1o7rdu9QnUdlwu4iquOh/eKrjXhO/SSEsEXYLYsv4HoOgqhGJu0n
IthaIUjJ2tspruqGBGyMQwD9LjR7/JhGR69feZeFTxjoPi7taq8my9gxhSZwJob1tDKWd+ChqdVL
7+DwSOcr9+eTUKVFJCpEl0afcUkYg/VoQmpqUKSy0d3LKTEqQsQgjg1gHNuCsZEcwXrDVh+z/8/O
/r03pdW9RyHXtTxplNm3N0umyx+mCgd5KXqY7I+6vkz4hqlp5mWWd0vHZWsrEymMnJt/IJnXklJe
dUvnTPWn7pe2EOh+u59JaiscFrfo3dxSf1Qp9fZvmfWiwAAqAnHisEoER2yhms1SbHDMNYF0Um2c
JvTuMQFrAiHOSXuhZEjbRkgOnB9dWrA+oUs6Wr+h/mGGe8Wjxz2b4HCzPTL7Sq2Eud/sr1SBYTyk
L2A20KAZ6e0FMZgt+2hsl9jKs7rGTiBUZQcuGTr4aP08vB2lP8xdQZDMbCIiqb/O1zT4KkRQ0m9n
zGLLcc2GUUjF7UuDa8UWIoqDvsCBAZDpn1fvRtbuyxD2nQOR5GrUwZmaCywjfT4NvY8kqTXKBR/X
srPsEnAjmAAUEI84PKH628ikIw7m+6PKU9ROkdITwKLmAhxbuCgD2n+xjuPPVI0PBmOcrZoKPLKF
OdZ1TWdZd1aLMMSqWGZbYVS5CB2dJquYXT27lxklz7JUX1fXiIxbtqPkhaHYdT2Zb9SSPn8HtxZR
01/TYfPPrnVKQZYUB704B/EiHckiVhKhtHuZj62wOryYeddWI7H+VPoDcEfofyaWCcUNLmUmX1yy
1AKhwGxqLii9PLtrTGleYrrSv85K6VKZAuDLQB2lGq9uzIC8o04XOZezrCLbmm+pbt4D4JSbwC3M
sFqOyj2G0iRkmOtn5NmmTpshvum90PiXzz9jMFy59QxHJYrisWbWYQPVF3SbLAl8IvlBjOs0g54g
YUZNrj1MekDiRIKxEq7ERF4bi/ZoP1pLq0ebvL80lQ/XjLDST8C6MOO9WCQT/LD2cd1hPQN0RlNj
F6eKbrt5KwkP36q1yZR/0mHIjlxym+Cm51oVBXemKgvORI4T20ImlQdf4c69IPknGoWBpN8C2/E+
3Rjd+tLb7nZ96+nA795/YwN37+zACRPL0utE4tNJJDewUYY/3TkkUUk+NmcQCm57RqyMHtW25cX1
+B/akWjwH9X59w/OOOMCcBOKBK7GXK1xN3kePi8V4j7z+DJNgXMMY3lFQO3GrH81qIDbv3RqScUP
zXmd3RDggFboomMzVhIl1bXPHEAm/i4rLfV+HYuzhjPnTw9oqg8zlSdG4+d3+Xk764HhjnUxCcOR
aEqUFRHfC1IR7Ny2z3eEUF6UX7KyI6ceXiOp7jj6s65FgwXaPv4MMUvFe/MslvKW6t6qXN+Oy9/Y
AXSRGp/BZPCZ9I4vxjdsmVF2/sZEoxxDJZvRB4stJkfF5zmaGEbTE+Rq54jNyMbfI/PB6ceay6Vk
8H9TWj9BBoR9QQMHHIeW9vfkoCwum63yjnOVCMeuJC2XXfWj95QSFayFRB94IC7oYbiczxOodPqh
UOXRUWJIxpLrhAJsQVipbcmgazJXbRi2mokqk24UMPZDbDQKQuYFTfhH5PnZEXjagyNrgpj9Ck1V
8ptkUAWPwCG0yS6nSY3tj4yAg8RMUmGvFQv/rGpdemNmtOmewtyQyGmk2ukdsZaJp5ktDyrIcJ4/
82JO2LcX+UXJYNfM9tJgUtxMSid9+NVCW6oG+c5ZVET+e+PxKvnO5ecrh49NDQPQGShbr9V0B7EM
du0arY/Gux9L8M3ffdVVR6RMcJyMoMnbIOZBbQvEJQOuxYYylQ6KOLGGtubtarwp0sUSB9Tbj4T1
8A8Q0xQK5MQ6NRJlcclIsyvJ/aFk4znXf9HR3kA0pCaujfEBo/R0nYszOvJ8EmVLJFSrp8+E5kKJ
yz+Vhh4t6GL0vwWuh1C8SB73qYzoWoPo6Mp5EhvHAoU+NcLvih0uKwxv7Q2kvSBQPUmK8QXXUH16
fs3ZAUq2DSh9hbnZwfPgR6TLyNeCgpJve3paYlKZD2DzRfh0DKBz/rOZrccSchtplB7aek+K8rXz
h9Y0YnsIvdmkYgvdjUuN7NP5Ua0eYisaXmJ/tj3JWjZMau7v8tLT+ubS/VHGagrFrIVQblwQP4Y0
e645XJRmImCNx4kEsJ0mNncjCROFS4Vs83P3ok/i2m+Esilw3Aew6N1HDZSRHnjcdgrOv+uCrMUO
Gsr3y3dGWW23slwkvOz94Ksg4RnLKiT7cCFd7vCRbu3xI+TVYhMRX0Rc9R9U1RicbFpeSq9P5wEM
AtBWV0SAEhsYgtYVUq6heFl8BE76NwXOj9LGKLlCU6K96V988SBve19GOxbPkTPKsjhwPDNklHs1
Ou/ESALrDHpbVyRO23mTQ4YaWcs9HVyv4qE3P81xK+dX0QSyfxtGy9iDvW7zFvEVh2VCJgx3qVio
9LQe3FXsj6bXZdaq27KK0wIRenkjbxWVdGPpQpuJmM1DMiqVmjEChNa8k4utWN6I/FvJe+K53MGQ
/wOaUxflqkmYQ2uu58XM2j1vloRaHwDbVq+SdwCpCLlFm0uqV/FxpyMRnvD7pcsfiNmXgh4cnM3n
pzdSshB6SyJVZuMq+Z0DPjDE6Ei+cDKJrGcM/YhCKHiu1OyYIP1EMuxwtgdVKUCObf9Zm96aFQLX
JbKnUyayZq+BnLyc6jvg5gVty+IGaoj0a9AbQqS5u+FwEOkNSoGeCOpZCVVDKefAiJXqhPmU3/N2
4dMctbXaMc9KmmCOPW6ybW/YxpaXYP+UQ2/gv4XGp1O7r0O7pIc0Y7qmTamVKv/jg+lRNBs7txJf
KfhkVb5z6VQvD/HrB/cH8AX/0FHjEzhKnl2XcF6z1Hupec2S+PcHj16vOS5EQgls2FVpCdiXbfer
C/4Jlgk6GgZwL+/uzfFjl1B1PjSLFMCoWwSU2irW9T4yB/fiDQT0mCp1NhFk/40s02LU7lR/d5zK
bc3TcwCxX/0p4zQJg+04rR5jhQwsXmZIuZREyRGJe7rtLI1z2fqx1X8pAVW0uK3IJSIVD+cruG6O
zbGfTdPH157Km016QteSwas7tzjGAIHcb6jsHWDaPKy5pLYgh4jW3IQNjLXgFRw81D1l1mKa2vBg
AwjDOqu+TzFybMqZnnJIGFbl2MXy/Q+8Ed24Wdq/zZbEUz4mEOqj9ecMMwfdugcv5dPuXP5Y7q49
FOR7Wc68guYYNagaF0kT9eP+XYvvnwOIeplHcE/DguibtNSCS6CyF7A7I1WIE7IdJy/zL94TX6WP
T7PnIufHeK9dIiJy7c95GO47uVFv2Exk+gckRKsSddeyl4ouH2Qz6GWfE4uM+OKyJgQs2cNugzGN
JEciQFYmvZusFaW3AE5R8gtePRD6nKuIo4IzXoL0COl4XXplyAj4kjR/eTm8n1IQIuj+5t+s5xH4
O+vSdbM6FX1EuebPfTJk9AYQO9BMhSIUjsHUMdIAM+X/ryHZTNCcAi5MTMjvBS+4zDRUa3uAmw9X
3NB5G8gaJ9B5PWWypZMHCFOSLHWqtr1ADYu9CyXV+NRQGffxCeUBdr01dM0OJRxVC+XjNU4VKeyZ
bY4CoXe7V/rX1Hx6Gfif1wLthKjASnnNrbA2x3V7wMHSiUIRCNNGvgGbnaQWxX3K5VYCwgXIcQUs
Kfbg2Y+39dOmF4xNfh8Id1z3u78CqMK6E2Cgoggkcw42nf1DOmgoysFFLiRYB11MswWBkXekwMF2
H6EjpyT/IJ4tFDiRyyL83uA34yuCgnqiU7q04jyLN5YGOD0YDImPJ+peLXfDQxB0+aKT2pywnSJZ
tEIP6AxUjuk1Jr8esAUWKO3fg/RrZYBEpFj5WpxWWYuxGhFBJ7EC2v4uOPaAMFUPRD2q28TZRR/h
GNQBol/j/vuLbXwVOi+An+D832GickEB4FxDXqOu9h8iiSmMf+ZlDe4qRUFZMSMm1QRpXsFydmuf
p7RFGTj3RYCc5Jj0yU/4aGTI4opIc1U2zPM4Sz6WRqA4skrySNP/Ux4DGQIFWIbSR3WrCOpELvv5
bC9MOseaKbFkdMtFMPRScSqMdrzhJlANFz4Zo2ytjtXdLqeZVi42ehbT0uUYHBHKX8PS0SNWMwlX
mbnSyfaQeHWk9nasolRKy8keLStf5dnICeQBepLp3xDnpoobi6qK1U/PszfN2NA5xMGL3Jr6a79F
TVrDrYSVm9IeYuhZZXzHBkx5P/WgvTn3ifUCRJoHXnxKU0NnO42U6Yco5w5JOvY4TgCj0niGxFwm
vdwbkyXXtPaQ60vV8jdWb+ZqoTrLxBvFPxDpzydeCxq92IEnT0txbc+RstHbpGqDSVNJtWezXlOQ
3TvpZknz7iPN/Bl5Dw6g2wHgmc0e+e+RaEllYxvzZdGN15nMxiuQT+SK76tj5kK3Fd8iepuJvyDq
Ivz+5sXNWAzXtH/3aafd5KtcUXtiMLwIvv2jWTMn1xVaYEzeYSUkfeRipXKB3lCMAbe7yegmEtfy
ocyd/YKNeTcELraP7LntyGdLvF0YWweXJLpUuyDC5/u7eqM/qAtRBVARu8puc4i3UzT62UM0vaxQ
tFo7iSXV7jl+EwQvXw3ZKyVLgpgC45WMnw45aXolGOI6YyELjXW9mqbztxqZqgWMej6UkOAZO19E
VhNfqmEcUDVUfH3cSPbl59RcZ43JdclflBgzUxNHJUn1yEbK7vyDuMsGyBt+9Ko4ZHO7Tq0JEEq6
K0Cv7vz7rIYVAUpWlBLb/HtgweeEaPqPtZXUY0aW3gG8NAdIsgFYYgHbr7RIUL5M8suvykN/DLXi
tZQv/mt+tpc66gq0yOVyKUSgzfXI7/x43KomAxChHChQ0EX/7BQxA9V30r19v7Mv9oD6Os/SrCT5
S13bjFAmANBuTAYmzcu8IWiuTGqlipCBUntmNvNFanC3NYUGYrLIiouHmgQfFube6zTQ4vz1apON
QXA78jnE2hOiaRUuOCnRbZiohfhDJjx4VDpk4YVF6uU5nff3gBb3FD8izaWHefv8rLXAdCNRBLvq
Hvt6WP/KSOs0jsJxlXlY6ORtKEuJ65mWb/5u/oZbfl4YrtD0ruVQj9j+yL0esJfjNgIgzh4/WUo3
MLMdqyc3WzCWGU2gFLL32OK1QyDOdNlhBlJMFuaWbMTSY04alWL0QPsxqINCdLUl8/dD843a8lz9
7o1XnZgzP7g7s6iT2Y6fgtLZSCk01jWY4wYvhPz4rkimTuEKy/Aj5vUhH1xBgzJxmQHesQOSS2HB
4ZfThwDFtDXr6uiA6dGrqFEcKtWTJ2SmU2j4fMPkz8S7krnxrr60ZlyCbjybtGStzEIeDtqVbL2g
XK28LyRD0FeddB8toysW9MR1w/hozAmpv+ssP4gd22HYAO3T75h/JNjTigQ6reK8scQ63DlZ7hii
5Zk8CvDGWe+pQS3ML51+ha/g0FEmB0IwFEzEQOwpMG3njtF7o7Xu6GqNMXFh9xDr3YVziStEXx4x
LJIDJYNwJtZQErMOsuHE4zWmPULE6lqWD2a+gINLS21PKWZr0qcsleMQKA8qkO60w2MhKJoqnP/a
rjnOdqXCZvzhNheujvV81qZYSVzH0n9Qt6UaLUeDtwjy6wAR0sP8YFo4M8kuENnMiYBETjCWNuOM
hcLzNF1pyEpDL9HTDn912txJC7xQIUJ/sxKUx8hOtfyIRZSHfVpdOa+dsCTY4NZn4rBpCIPlaJJY
zjQ+PKdqv3dO3pOQi/srwNNrdcJmsLZIrJUAsZ+TYapag8VwdOhN9JPBXOL7k9q9EmO94zEigR53
8GTMgz646y0Nwkl6EntCb3d2o2IC+Gp0YaDhVb20tHiCBIylvQjKxlY5F+3mIL7/wj+YXmD27mSM
Hxwz9fELFRYmcAxLAzzRdDe3sdtIpsvEEQEPEadGWFCFZK31qrGCu9IcKesT4jPl4iDBGyKNb0Ik
aseabraSOZE7D+ErioQzoGfhbQOWORmcazGx9lLKyWn6RsULfcEXgwTM7PYnKi+0nIY0Dv9Av79K
wGHSzk6QPWxsEHk1Fy+taXjhXvGz7VzHlW8mI+fjr5i5tfUrC9BSjcvC86VEQn8R2DTCSSH9AFWh
WKOQ0iW1qg9m9jjOpQ+E6e6H9crdshQj5aLWAdh5PA1Gqsa860VOdIDvaRXDSTs3s/YHP9OIGnjy
oGVLF7KEuIpQscEwXFvzTASbm8Is33edv6X/lKppsNN3jcAlO9P1qKCy0g0m04/yInB2+GXhI9Md
UwTJu8HSbXCQ3DsNaP9Gjz8HntuGNZtl+umRgdEIcx+ZgSOg2ZYM23rD5AmrOHiLH8IemK44TiXN
rdXDM0EVq4NANFfYCumAsm72uevIA7wllX2Kv8kqe00PSctsVc5EyFFCZ/x4r7/iqizY1tiBw4TA
gT51ZmYZJH5MHJgIJtXmtfvs0bq1sp7WMNtTI2yS1fOl8dqEbROnVR/ALEicvpDhodnO0z8fZGsR
JLdkiFXYbFDXoZrOjI64zjM6vYTb/HyWCv+hDrOjv5YlJ9HROPqtbl+UAV2WZyq46i0quo0FOj13
Qz0nflmkCwChYWd7ltt6xcFt4Ac15GC+DSQNnQd7y5ce7LT1JXo+beV4QEZpkbQacOG+jd/9gRE0
LMH2spcjYMQhehqP62tp34qAd8enPogXDxDwgg/osxRfxHPvnS5rX5afgerSYVhIsxjKhG1Jyxjv
+P80SYPAhNgLPatB3szYNYAhHmUhWEFuXty0iYxf54gVc9Y3lV8b+1DEU7vzOJQT0MxtX0nHdykJ
wIsN0gf8gRdhprJXDrO/Bmvpf7jKv4+ttvdr6ye6/cnJWZIWHtz2f4O4IvKo+XJnaxn4mXGdML8e
oz8j98r/7uFTUb1Ui0+J/NJZnJ/6mXQItKbygVSc43GqXLUwV8yBPbNFJiKpky+RPVPtRayqezYV
HJwaL1vUq/Co8eGKpKFh3I61kYbiBKzf1aKNcsywVMAqP0mHK7aML8tvRi8a5pJbuX5rbkPzYSVJ
qqtYbqhRbmIFFCDdKQCRg+vOjCMUKP1q52zKQhzVcffvyucKxA6A3kvZdzjAnuPSoCxUfKoLC2vF
hXSaeCpsXbNLCv5Nw/OTOSGiI+QVL5DnUgDIQZePKihbRgnresGIC4KQXLQzdkK7fHq2APs6AaYg
Ytpsq9UBGJtl0I8gxlGrPQlVc+8zoNOHk8nfuEznttZahHXWr7lirAAmFYsDdvuGDeq3esIPJ4f6
E2d3HWXcNj1/hBUntXgG1sZtGWruVg130u4c/5lTIenCPG7n3f4zcZZXCjEJ99/zPRGC5j1q50jR
pAq1k0vWJQCiWGqqvZL1tI9JBkMaOC0MldIVMbF3JBjyOg+uktmKfetTcSskd7dFfDiBIjsJYD39
Rh+Y6KeMskv/Gm771QlnAXFJByQfAuQhtBv+SGHxm0lNI1Q19AkBu7aAOpxAgjqUX+vWRsH7aTqs
6+6a2FrWoFtrjZ0P2LRZS/s5yUAqInHffWnSTqrzUk9YJFiM71CUaAtwD/v4u7F6ZNJCYOs8OQEM
gny8VRw78sfxTk7DxHxiOPNAGXr8oDMbNjeq0EuGJUdgTiBbhhbFmBfh5GBPHOQjzV0aUOcVHiJH
1+7S70ZIim6QTXrjaUh7YWkeo0CfyaWARh260mtcIMHQrZvrHZ2B2kTSr93NEN1MU+QU+C00se+3
fSgBjkAeKAPh+qKdjxD/6c72bhCfSFwHybwzDMz3oCNg8GpEIgEbiHfzshv5Qug4qJRmbXDNSg0t
ftiigLol6K8vqcuFJKCYGF+uj2e+HhyYuxwgYfCRdua51kyhCht0JcGUUfsVgQih8BRuY4zMH7jM
rCauhpwrNtZWcSrqhXPNfoms0UEpgfCuwF8zIKnTx790R03nR+UBLacdmnootyA+vHxQeWGBmiI4
vnnodK9JfHNhddKMZqdnI/y3AzVbmPR7LBxEHpGYHly1QVcoeTq0by68IUMuuwLrB5tlY0fPmZkV
gK1+3xSSIFsN9nfwNGLdROLFaOYk0OwFQWg+tDY6lwomSUfPtGHFW/EQf7f4y6Csjelz5LzsrodP
n2cqz6o2KRJiJC94crM5stqCPaDjXuk461BbNh1EIsNEqv1duu3hDhfZ25jq44ovOmEfMlzbnjes
8aOhQbr1foPeKmQ7Nvz+0VxlAmFyLTAPyZb57k7erLOQ+BB2rrbkvg3aF8mpovWWg3yZPhuD5HcP
bmuF9S9XjkEVViudcsdG1TJ/WJBZ1bILZ5lFOSsQheDu+O4J6eZDYWqZgVLwJBrxvyLBh7WfPoYu
5giJW0RusuVdpBDsHV7hKTMuhVAbRqvqJx6XeSL09KteRIzuz8JfPeBn7Z91H6AIT9aqhoUsVMGK
i9lJss+zhADwwT4bE4liFjTZ4kQVvuV+PxuNKwQ2aKpCcxunuhSHBv5eKe0RaBAm//TydM4wMrcb
qM1mQoPN5L2BADH+FQO2MymZHIZLq2+sGrI8qvq/XZ6qvGaHj512DHlF2PtbzjliVxSjG//qhCqw
NDOYH1zrlKceLSGHM7RLycbKq3a8A3St07O8vBEA11tlRFpclUQMpW6aUIRdcEyWg7E57yAV/R92
wEDhoe2+KHnk/GhxRePScDeXY2h4tEmHc24VBZPTuQ5mFletPbAL155i9EH3mZ357W+BEYLW0n34
5ZTf7oWDAngDlXhLTRK+KjLLTfKKfkpCth2TpmbJ82jSGVXcSKvGMMMRprAui31v59uV+BXhkEVx
ntT1+GbLtq7DJmy8APHo3vnIYDSLWhTZeOlJ+RxXGe06H2uMexmGMB/yzZEz5bvpCkUsvEoaC91p
mxqqsILZ9T2TYM+P6WYQT2nET7Gs+cs9TTIhZM4vnmnu6rXKXErazb0MYayRhvHM5Giq8yRtEavr
9E2xS2Ys/lR8rNxFDjb33v+RscJq1tz2lRB6re1v2v+FJ8F+Qj0oG3K2+8zSyvkL7CM0jCJvRSGl
df1EZDs/Ej7h69B0PLZ4imhTrFXoypue9I0sRpNzrUgtidIC1+msc/6+KM0gffikdfFvpsocA6A7
W9BmNGxLKMrlU2LNxgdBqpQ3nT8asKPQWkJAXPLZZzj65ST/J7Ton2YOA8z2w14STvYgiEnxi0Xs
FkCZnX0BBFAYUQkvReU/xaVXO31j/ma+Ye7z/lGM2Nm5ipYdQMy891BrH6RrO2BTVdldxsdD0Kj/
QXA7IntRXNi8MEfaC9Vuqjqi1Jr+5wulNW2rC5sS+2hYfJIR2RTQY9PmjpZgI+NiKAioulOLTAOB
Z2MtX2LDzisgx3B8XC3KQ7VdJ2Qw9gygAdC15IJpR/qTy0mYyfBMaFv0VvZKrm4TaVzZ/iAJMbEG
LqAf9bgSM/BLUK/dS7SApn5MN7LG4XmfJgguUwkBM6/vAA57J5EdN0EvpSdONK7bv4Sw/qXwwwqR
fQkg+3Jft3nyUa6lBswsvqT6XBCOZxQIP01Rq4teo9jJDI5g80Vrj3pAU3E2DYwL2vtT9F84aLPU
IJEkhrh4ePke1jz7STsnNmr0pzwzGxAP7YPDrYvJ95oLPZiEynqtYgJ/aou/RlClhqWPJyP31WsF
5hsK2mCaSUWlTLxdj4VA9mmJbxC+OoQq1QXPwn1wBN0Vp92ZTx8/tQeFpIx6Zk0C2WOkvxYJ25DD
O0Uhxq9rrknCbGhbdkZJRuGh2lI07mIdAjsIqGu+tq953fX/8Rj/agPzyxgLhUM77RU4vz0GQ8fZ
KKBaiGL0lZn/WP1seOjGWGiCtv8Ysbwf9REF8Kph8bo8fKpFvM3WgLuJm/fUC2ihCn3bGv6jgy3t
0sKwvblHgoBvCZlPPpzFnK2DCqjuuNBsqV34asmePMnb7JOA/f10x8JvHRXad2hhZd+GdWROKp1r
pZBmGz+M0CYKuqoqb+H2fthDbhFEADoTsj/MESxW2C6u2Ogp1hzJdTCCdsJLxu9JL0sLG3VFPX9g
886Wba0LgjI5TH0YM7qfJ5/Dxkf2xYA4k489r4EIOdcEBv8llMwlTlwKh0BvT6kEw9rDDTG3Ikoo
oPeHbdcJS/UALXTBrCMrIuIVc7mDV2nY0bwdG2v5N3QpbvDdl1VcXiCYg2sgRnpjqzKO+szIlQ48
mGzRULxCo9P3c3ale9iYKi2aKfMCahBkM25OuirTnY9mRSQfzbZXK7d4jjmXJnneyUXZNGBcDu15
5sQDpWkc2eREbdnrANTS2m30ENeNVEiXRBxne1VSSgxbppNPhaWT4v10NvIYpwvXZWw+ZzPV1mTV
SUQY76O34Ve5/HjjIHzYdLXUFRIaiFpBQPv/IL0DkfaEo6QM7vfn096bf+sD19avyeys3I2reXBb
M3rxndzxmHj70rrBh4Bdp1CnpQXyE/DXNqAn78fTAkgFq05jYQ47U6MqHVZOZgQ3F2iRtCiEUEHX
i2uS7ENy5avUSJ0WQlCiHKRY8VN/2ZhmoNWXsaua4jbF+LX5piw1tktKGaNHKiH0DxzQEG5eXmkA
B088AGIpBn5PWeCF+L/m169pHsZ0BrNlYBVccRdRIgRnwhUqMlNW4D0HzqBjtmgtHek++m5W9lMb
BiIWikgjRhhA1eho48CE0gurDOZEuLV09OXNgk6pAoJNEotgroaB6G5TgyeyqnxuDtINbWP/f+1O
o6RLDUNvtxxXaxhIle7lJ77BWS9atWi4+VQTq6TAbOeDoRrk47bIDM9SrnEBMkBJP+I3WrpvAUMK
5NxelqPys7AbUnfEpHNtym5YrePdl3d6+7PmpffiLX8UnMKWHcF6KztFwjDoXdfZLwU13g2HviNT
Zc9+VwA3XYyUTKLNDQLNI+Ijlf3DfrVLekps/ZAs0Ah2fle/Lvj5UKMtsL+TtFbGGmgReeSZ9JKZ
9g7KdnV++pvH0mHaqMwgMAsYoBoh0djbHh64iJs/Rp4uOT7ZgXpNbq/WSYTT+1NppJqHKBI56wGF
Nn69bI60oqnaPLqAalwR40GpzVfs+kRgzIystMecIMUy/WYJyBqn+IxCIyazVbT4lHzbwrTnNaF2
B9pQwyAWGV2rflCRxif5SLz3iLuK9DU9gCdqJ84UHCa0baGIdnXAF+OGZCZ3NHvY4bdaL7jphJ7t
xbYW9L/bHSoF1Fpcd8k0GlTqYbEDolCqjYRL5cDt1HqmsyYzOkklnC+hA+F4XXVxGyXphTQD6Cwp
Zl8nGvzGSCnIh++rK471K8qaMcujzRWb7zYg/in8NIrpAxoYXrhrnFDQaDqSE1XTjSRpnV4dxexs
4i7FRVjb8JTKkW8KFEmpUopEnRX94Tr+nlyYE+1MypmGxY+MEcpjIXpK812b3R01GTHb+9bj0ROo
Qj1UXCE7sp2rZi+MSZrC3x9PS+FqnxBt/4ojv6NryCOFmghFFs6MBmfpSpH/teUjJxt2WsH2iNkw
yOSnAIix8B2EVdLGWxCiMdzCtkjOsEIWGKv530WVATauWBwWsa7VwZZnKa/L0hbvjHNejYgrmAvb
tSINyd05ZPgBiEy2geCkS2m12KE9vr3oEN8xrl1z9ta77GcpvrHEAvBA/sucxVBqNnmg/jJ9m8vx
n9undvX/ubL7Mb2huVLHYMZ7bhchzjQSTtwKXk4tce2iBadrA+OuUk9zZZc0xzPSKJaiJ+XV9t5e
YvPUR3zqVqoOMURqJzi6oqZlDanUc1q6XJ96Oz7DuaNHcsYgWW7MjUJ1SMvJxhGIchPlj/rf2fyy
qhlU0k6oD052yJVWyiiO65g+iRDP9HU7EXffJ1VTd8et1eGmnuq0sb7B9zj6e82oCLyFifypqDOM
PZG2ffnKze3p5NjseBkqMaqm70SXPRH+iAhE1k/mdK0T5UVbgJ5PsQ1wtH1zKwb9Qfva2qy5/O97
DZhkg92iHwPGuhp8PvpXOqeSHMasiccuylbojsiAr+WNlSJWuMcSnmlIQt7Sch7fBDjjxNI5AH2/
Ae0RmbiJURobFGuhySoSbIUr+91qQCzpe3rMono40FxzngprLEkuk1VguffzM7hCAypfc37Jd97s
VrHFnSdQgaTAz6V+c4WJA++fLJaXjWcqM9GODLRwMuTm3HYe8n2tERO6lHcaPl8kwAWYloyaWGG6
l9feBNDZ1xDG3Z/U5sVb4mfWHMdWfs0rRkZK44z+3/oYrAQ/FNqCbDHKj2lRzBwfyVYYTITSQTir
wO4wr0s73ulI7ksmBFQ/HEhNk7YwMFdjuXff72aTMWd3JALq6X/b00LLP6juwZzuG9iomrDia0Ek
kAWU6cR4DdO/nQDcFQ3Rulj13fR9zWkiWiYnGIp0vNisy9fkjV64Q+GrhOk+1mH4XwfWQAC6oH3p
cdR7qsGeFVuIxHRCoBew5ZdpJMhj11Sx7I/mEv1crxZXCkS/oWVS2LG1nrCF3JokehSBdszxtIqu
JCL6f5IrWuN18YBVeI0mEDgyxbFVVFIBtoUbxdQYcs79+Om8VOJDZZ7Fui7S/eIWYZo6TJJcv/db
IZDKKGWyCj48hUSc7WyfBgvgw3QsLZD/MZt/ukqPYW3VTcR6a1Wo++1OLkdW+a4SKnlma/xnOkUu
W4oWD+hCJXN4I5oInHLu2p2blv4wwj+0kbOAuBDVZBwOZ/MO4YUnwgy9Wez6LpOezKGgZZ0BoWcO
3GYQdBKxGbDsteQdFRA9VMsYI0Fy0htVThdrlCWv4LI6jyutq78rLdLLLZoWkuWceM88a+UEB9Pj
1Sp4H6CJNdwmkjFT3v92Zt1JJYdrdJYJztrnVhd1+Se7Iz7liQFm2RSJ8hv4WxHkLuNeRWU2FRn1
fLsh8EKmFZXA+AMkNaNC++q2X5TfgyLjsDh3pgPnozaAYN7qSTREx8ffX9zUK7r050sU8O0cE51J
iYwVsVKDVcqN2zycB7eBwDUuVZNYdlG993xULATXOI02ekWcIjm1p/K0mGH8eN1H2K/107HaTGaN
6u6+1CH4ivwRIyomuNOFYFLyFva56XlPxscyNhvRkNztUVPMEZ83t/enb1AM0RVvtPLQR+ry8Cod
fu4bIv4DQHHbLrjFCE0XmVjq8OOUqhuixgzq589yjGFc2ABD2+hJhPS0zw8ca3bMlR3CYZIdEkw1
dNCkw3HXcF0+U0D3ntaJbZUm+SSVPepXNAtG/w8xUHK6NHd6/d6hjBaj1sRKq6dviWzT6Iz58TWf
YG62aIcYyyGSM4DgQY9F0Syen6rj6FtXGz4dV0tiKv4abtchfleOY7q4CU0QCPVBvVIhqKWL//RP
UaZwroL+jV6QLQKQgNIVe2gTQVM9Sm3gzcUyMcEyArX4xDNXxed3L/iksqvwRwn6z8epUgI2LJGv
Yx2nGVhBxDy7HW0R3Ipn0E314D/i8pUtCb8GuY1PohIB9uU5Iq9aC+cdZ9lHzysuAimpnYYwhVb8
FLXAdXaXzPOcK6+mh77SMYYEqoqPJsmb49zdLI4BgegiBG/LV9QknZaqra+vHIPWJqOTiCeZfKri
94iW+qT7wL1NJSLBEKjfohkirztsm3QwMlHDycsdr5wj3ynBmMy82FVS+GrhIwntg0EhmKkqYZoK
COBdSmcaEb0iwYs5C45ct8NTXwLPJ38eXu75UtqkDUuYE/bI7mcJJ1m+W6zVSHXCRK64ba9kvZaZ
KUAJFWPyru3/6DUEwI1atRCiapG0VcIbk4au1lHSi/kJYb7aH5MoNYCBgph10fmhQd4IaiNw0SNj
CrT4OteZgBZK3jr8KRs/LbKLjF8tCB7oOZ+h4MVEBd1izclainj3L+/ROEyCzVMwjqS/PyRrDcXD
wbjJ+M1zCikPdm8CTnMZFhomas056BoG2j3OGRErKCbVfNSczhUSRXP86ztCXmFTSnuCr9DktwCz
GPtEE/zP3IGJCkCYtvobM/0tC0exjauozxcTqRibW0dEG4AyGgPqj31xtelvPdnILMqy94fzs3T2
V+CWTEORsxyefv9HPD+ubnnuFbglPZ2ca6A1fa5cvt4+eBwM1U16uAiRGt4xUbThVc1SRFmhewiz
i71DZxtciX7qas0aco8AQFpjchUraYq7chkS78ZUhSgKDXl46fgPNU253eiT/USQcKKFFZDGvYXM
GPRNx4Hy6IqDPcE0XFvkDfBhYOTJgZy2ia7RAmDNI/ddUsAmb6EaAr4kqjGqmyqZITa0Cc33JEpq
vOJn5eygpEyyNgeMBUlIgD04YiTA3YA/d5ZIf7aRPmXSWUgY37DZifWRC5yGRmmEdzGrpHjNeDpo
FkWv5G5+pIkHup24RSgqg1mGWNUtkv+oxRUdm2PVo/ptRDeRS4CTSOhT3h6TvziUYNFkRCDoGx1e
ANkc4Yr95DP39Fs6EZmfhVkEi6wr7CvVSKoIlQrMze705BjHhxeKHpgDO3bQ+fo1PTrWvSAWR8zs
s/VmC/q0u2CM79HwB7htal3ndRNzLU3zWeN5nD+fUu3mmvCdJop8WMLi/UqW4CjYVe0C59hi+Jgn
CAtMDXyIK8jjRYDsZxvEj68bYSDX73/B7LIO19CLdQ0YB+R5qCGEQOmo7CXwG1Ec/jLoBzgTCFvn
vYqHBm1jfGbK4rEGFu89Eu/Z2A0KqZkw1PYuTw1ozH9bdlF5QPAr7c39gTDLRBjgWwwiLTieLB2n
X2t7ckSNm43orgdSr+BasLGfHy+K9vCmS/I2OaEnMlXW7eNOAjV3BM61vof/bl+stNCAVzymES6S
Os3UlpJEXQ3M8RJhOWoon9icip7hrffMNhmDaqDRKYnZJRnziWOJlSd9Pl+ExGcLLuIiWULc4Mvu
U06oPiGs0nWMr9cFu/IEqCYORYALn417Ci5XafZMB29AtobG+aVmhSWHoN+LGDG+TUXwkO4UZdbS
7OqI87x5UR95/sJ5Zsf28noCduXi4qyC3ngq4aZjGMYW8oPAi23BmzkSDw4F8gm0ReTRnkfxeWEy
hLCFDHI+DJ33BGo/z2dOnhgK+mLJVpJof1i1UOzu1anmJjh8J/coh2WoO3IVFdryISjPp7gmC428
nsVjRjpFR5lSkt7r7DU2GBQRBbQJy8AoTyXygBQz/6qgcgIS2QDzh3sglFPTlhNYWlzP5BowMxsC
6PzodAJoBeAxrqIs9WYh1P6GrAnmY6e2qyeTJtgss8nHjnD9ERlXjOXIZjZQ7Y1jjSavRhTWFF6A
qmli+jAPwWXlt1GOG+W5yzFHNVX6t7M+1jRZKjWlPx21DKnWH9eEplHOryAO5NQ7vKingPoSz9fq
3Q12Ken9dxG8UbQkyDnN1/hJmtemNfnrZuiN+rpphVSm/oyeV3kP9hpC1vGOFJrzaYnIM+7eTYPK
YIFv93qOLy1OVMsjeX5OEWUsmTdsSK9SfuTxriTSeozNcVa6MpsC7Dka78re6AWZfgErokOgtmwo
1ROP07DBRFMbgEzrM7vzadt1D3DFG/iTh5ODzg3MQXeVg1NZ/Q4MWPGSKA4UhCzusKTeKfvHlAzU
PDgisgiL6xBB4Lkw13r1u9ERmrXH+HaDK7NYZO2V02U0dMBNpgq0ASp14ss28v4P6N454RPNChU1
mG5IXqoQwsNUY4mBPeQbcvdE+32IkxELVFczAD1O1dpsCyfOHLtM1zB45G6gKIyX8zbfTmPd+bMk
NrKSLE9pKlXoUwNJi9DPCQJGBaBpl4rr7tDzd1KOl3YcQdofyJ8GdQr4R4lQV3uI6fFeOzpIj+tR
D1KYTScPrx7qIyi/yJU5Mi6jnkBlOeqgX+dswOzObKXXnbC2UrSTl7nx5NQjrl6yaHNrE5Fq6x0d
aJSTUVcSnK92YkO6zqC2mRezfoE5czirAxDfU0YtV6mc1Jv0w3Um0REZP3DGYX3CZf6A9MexZUdF
OrWKFA+U0R6OQAepGxSV/eaKuY2pOr/0JrL81p8ExbJ91xPs63dodnT0sGdV9zOhUtgwF12YVk7b
QcmSDwMnJ+a4lzu05vuMK1+RUGyi4mCrJ4oLALSXkEO/BeGnzLEC7GzmeTeRCRRPUFHRQ4f8dhas
gU5vSh+mpDe1rk0lCyU46SHpaPPVMyQA06UosMPMBx7rbG+z0UJLPrGynuP0SRudJMU9QvnfLZLd
Byp36/j5zw2w4TrRuGtum7g/m461gF+nEi9D56lJt8a3P4sUoc9xCPOfpkR3giBD2q+xkf2E3FZl
0tLeQHVSEO4tnWc881kB4EKd9H1OGiaPKg1c2IJuWNmP2CzlITnd0PKdTTN4NrVJjFl9MRRr/FEA
1pxpQwqOgwC+HN/bPWqO9TdIqgwXKS+22JtC3Mcb/uMMRX0sm6PRaGdcdNoa+fUVBXmQrGpALJ9p
kW234Isf0MNahV0+PDZRU1e+lcIPoF5zYf/S7Pt4zFhogaxSl3cTcZ5EUvkJKBOqY3emCyrZ8qFh
RUGc/p2q9hoJ3ShkmBV+itedj0FBCLh/AJalfaowu1rmHyUFJr6nX7V0epchYhF+2OrEpASBdxJP
v5bEOoN9uQRipcV4k6cqj3wlo1AuSXVzZOEa4kSsBXtN4syUzEKPm/G6Gk1Dhiq2QwOF4Xru9nbb
RP3B3JZNwefeQiQ9//nxtI0/kUt1vigy2dyNMqXIjvnPOUQth7/p3hfy63rqL4OWa7JBcnUTs76G
ftH2rtftSL4bfDs1Tp7aNjMor0II7Yctbsd2uho08RD7FMEkZ/STVnNYTCtBWPo8m4ZsSdyfbWr5
6bjuAamAIXzNnixRzr7maD4dfD2zleHTxDHHZMKKM0bGSt4O1rRYJuap8Q/98YL+s2B7UIBkIjMX
FGa/AX25zRnhPWQlPiOReKUoLMkOwePkyfZBpvnAoX/Z5g5cf2afdhoRpht8XWXlYxUpgC3h4GW7
nZalyzKs0KDl1l9zkbzd0B9UvMGuiKC87ZakDlB5QjxY3NFFPfyAGZIX1+UR71udIrzXAssFgSl6
Qb8JAszplDtyeA5qGmQdx+JVKAPHPd36R9HcVTdgareK+dtuUYdjZDCSo+qOf65vRhkyCKomRiAr
LbFIKbtU01cDN11GOPqv4bAFQ/9SkzTc72XzSIU82IRCxK3vNzDKH0WgRx9wpt8psoIUbrjdwbDe
4nUlRRKl5MocFK97j+AAl/BagaptbjrDGGOAfXbIN+fYcHQEOVzibhJXkonNeeMgxRG+tNkLQ1k4
DYWIN7PzPIEBNU/whWuTrlB4PnkIyhUBe6xCjjIGxrWyB4UBlWonVZwqXlsvcbUB6+zI8N8e/Yc0
l2qJ0NYErV3pc/9gtxgY1+Vyz4j214nOhF2cHl3aqyQNkzl+K/AaKxyDj/N4VV4/GuAHISBnG515
JvyldjEqG58ozbdt/9NZFcb75FTiHEuIy56bVdFZ4GEc8h9l/Z6heE4V/OzZBVBilLWwrF47YVsa
vWdx6IaCqcAmgX/L7B+n1s3mJFAQBHOm9wTbYBs9YUQfPuW/Tn/RZMeHA4i4bapGvX++D/Od0pTA
qs4xwLwR9KikH7oK5OORt+dYV3W2cAYYkW25abcStUQnxVf5GhZvPXKX1LV5R0EefN4xuIYHhj/1
pq/BugUwqM6hS6vu3TwIeXvDmUf69gBB3BT10ChTteUpEE5tc8cUupxAA1/RqQcwb9rlmnZFV3J7
VznlSXvsJbP3sNuOVqj7J/c0A+gATzQEhENBfdmznR0aXNrFOs2ibab+jmdsVoyGe5daQe6RWtyJ
VMNYY+4wOeUNywMQFU6U1hgNkInyb2Ux4SGTLqHAMeshn1qVN61lFYUZMrQrVn8Y6m28ATgmDdhL
Aqa3dl/GeP5TF8qyfTJfTlPdCl6dMdJEFYxjqPNX7iZg57vl7eXDx4l7wcwuG7E2UxwHB9VMa7KI
eWk6+RmdpeyMHEuWOTiaEYlFzSclsQ6o2lV31Fs+eswFGprduBY9Br6zW/0UvJjJ8petza9NnncN
80ouWvZ1Yfz5rhVKU4hAbWFzIqvq4wiirULPZRxTQHHOqvSQ+7uEZAK5Szz6ccCFZ0l2GTYY4TrK
F+O9/eFnXYnkP9S1nPYnwgA7b9LbYo8Fxtka5Up21q61ILC67Z/ISHkQrmwO6M4OAKwl03rHM/Sg
SAK8r/Fe/AKOFPUETgbliM3diNGADpc58O5m9B4HPVHOE+GmA5NzYZFueysY+qqNw/yuUZE5AZKM
PmjOXEnAUWo9BhKhnz87/rx6pz6gFOLRc62I2MFBxKiV4kaZiiMx+MDP/CoDl8TlUfe73ncgOqb2
yNdFrWOIzziliQoGtex0hhC4juGAa/1V/zhepI7OaqrbCBJaMH+3mNTxF/bWNisN6BHXME92vaZd
ggLoEj2J6DtRJ5sSyyHC4F0ay2hPqTdxiYSzaRpBaHGu3EGRNtZ1+KPR1V7L10JnvpaKLHYGC0l0
WPEZwsLwG/O1T9eP+lMuhyUx/E8rxlpLbidCSBpbbbmFoMaUPFuUE8BU1z9vpfMnLJxhaTB5XMlq
W/ELFpVWQF3emHYxZ3azifwAB1UCLvLE+b1csx4yjDEkx55TjonFJPhdptPCq/TB/ZuMRoLnqmv6
k39OnVX8CkvOD1vUq1aa601DWHhdvjkEdxUhAu3UZrpDA4avlaXJ6Gp+e2ZDhupgHWBEYCBg7L9W
9ZFTuTC82dRjungoGbnDqsI0p2rrKRRGxqEe0QRSPS7lypZ+rubfyLyENJlJx5DOB35H65eHrkTo
+3bnvYs1zLjJaQetzs8tupdDc5j/qt11YdPW+v/1yKoOl3uube+xG595LWAZyQkoqJjdSTeHJHzH
bPa6za+W8KLgQ1rZ10YhjcEUaq5Edx81gOxUFlflfqNubBMi3vHUFi8JsM5xunVw3l9HFoYAlxAU
QvhoeqCv8XX4IEwzlAOP92VhYvZIZxvpdyAEmL/aPPfs88uBlr4C9/jHIUO0prO9/2mIcmWYbOFQ
I/rkb5Tg6Rnwoc46Ue9SKElLW8KYw0mYNe2TzG7ZaB3l9gKJn4R4MNTzZcQdXBK7BL/0jBblt2Y6
O6/anf0SJapsGEVN/0J1QSmHLf6ot5OoF1uzdh2ohkxAflxGd7MvyofEEy5hgL5gh2i9rwXN019J
BdHSA6l+AFk063cuasRo3UkSu4zohe1I622eNDrXDVumcboUeivdi/N1VBvXdU5DR7VrBkUr+qnj
GsZxzeSc1qEZ80ZhvnEocnvqZbZxhY4J12fjvwU/gMw8Ax8Q47gat0o5yH50M8z+g16lvuOjvEwd
WP+oMZ1PGx2Vem/DE9vhDnlhNo69AX5uu4lh1JqdC3AhlGDgiTPms1eu3f01YuFQQgfyIjutdBli
EFEKdBnjjxgnn9VOAORwEbrvJDgRVNqLaI/f7udcO2WXtzlwfEsbAY6FBcM8Jz3LjMDpwLyU67Hp
QHeHgf8jO33zGddkVOQJImCt+lyA69eGeyDOeYO4Sw2cERaWtdVoEQWpVNu++yQPK3wS3lHTZJyC
d1goiI2so7IgfOWBMNK8MOVfPn5vKxfWpg1eQHTP9/F+rJlAKjt4jL+9tgvAmMLC9DTiBVxUIchJ
2YrsYc0O4EQ8NLPfuKOtm9bZYTs00kNDDjgNRu7xO0GSjbiIdzjESr5MND/KvRNs+AHVB0hClQ3B
ESQ/VHRG5l/SmbmeoiGZMZ4D5YKk9y4VSXS8WvCa3F4Ls/h+kdllfQFGSjSQ/qJZHr+23AhZuV4k
t4D69xI5DVzD88OOj6vs1a4JCq9n//WeaYg2D3xXf3A2AUnvXTgsaz+BS+x1HKJBjxIJNKR8ROuo
bLaE0d2fw7B6f5GDRXtVNRuf2bpqBIS7EhxxNdrl4MmG+8FU8J9ObzPfKQH+8g1eR7TZKmnSl5xs
+70kJ+bfl5ajpD8s3mu0gU2S5RhiNrGCplBt2vz1nxmyUFyRpZKAdgLyXErxCxNyJmY8Q00WLkGs
4elwaKQOsIF1GlGbb5hHVQy0vXIlXsC1rA8j7eCObegxu7VqXxFE4KdUC5vrfwutLJusUj3b+2NY
6rHT7dreJYcIhNGu9mBydyE4mzYOUsJLutjK/pGjbAFCL0ZnEbAR48StnJDYxrXihSVkslYy9eXy
Mw/KzbUgxSUxxFDI/1f4aJbPNYk0HZz2EqjmkfSOZsf9V9BY76m8NS/Jshf1yFFHipHCZpZkzX/s
ACwuzGcBxtchc7Shbr6VtHbbOggwZOFKzSG2DMHeXZepfSh5xldA9OkzHMLD7CX2Y4Sm5lzZDBLi
lcfdi/G5oqmNfxLAI7R0ySayDTuETBou+mr3bWUbMPNJomjtE+RNcR8hpQL/P667HlO+qBXnC8+B
ZCvW8T3XcCV3LEl5L+uQ9Ju+BmtWayjivybbIdWWALUDE2Z0ojZxFbMWasiKbAebV2DzzND19O8x
cUN3FLQRP5wpQbtMVk0U3S15bEjk28yvucsGX+dvdVHFGSV7oT9rq6GRncw/+p8rvwuy6MqXCLCF
F88LUgDrP0tA6SX+LXMFaS5hWlxst9khJYzr4jP7f9icYTjqJ8vnXp8UpKViz5wTorfqFq/Xt0ZT
X/6z2mwc2ca0ejx/9c0TjZsGryfjqosg1VIsEZF3IeoEmLp9b8HbKdUTKUJ1dYJCMmERAQdyXjdq
Y/QsHC+xG+SsnyaYqJDG0cnz2yNBcw6r4+B1W6vB8S3idIWSURM3U0UE+fiB/rlznEaJaU29vpn8
blUr+eY6MLAQPaJg4DEKKmsJthIMKWMVAzqDpizboP446nOBkdVOV/DJE4F56TnTqY+Mh2bxF3Zv
6RCuGouMsmgrsFCJNtUxC+8/iZFoHILNs6C9ixb8+IRD2WfVwR7HFJ+CTFds4ZpgTeGHsNNUftYs
Mt27zA0SEaFk/b3ryTOyVC5DSm8HuvRnYaXeuug+QtBEEU602zYH4ckpO4+8sSKfVwffJIrxC7Gm
Q+HcbHDOf0vYfaR1hfH193tWqWeBrXdo4+cJB9dMig7DWfIefglgocIZtt6aB5cdd3SgiNnBj5yP
UPmNJGxFWNB7xSVmk176bCC1gbtpO+p8nh04LBZ4PE8p3BC4NNECdlmC3qKUAFnhF96GLbapFnx/
sbF4igunV+zAjxre3M+DeI4eviCBDw6ObgroK5hqLCzS4YBPAjJblD5BmlOSUQG2d37afPDH8Hzg
U30Tq236gSpGgmTBGZE4fqlWtkNO1Bc58+CQEOdea6H5FP06hdvkNrqHOcbOKonnuliavGmYKAF1
xoqHWgrEqZeceC0BuBmGVUipcf5nOEr7t0SDBSe38HNQAkLCdwAKJJedtQ5d0ZWS+SKshu56dteq
3/uYJ+bizsS/cmLJS2bbW0ZAt10PH4Diyo3v9oTTJquxMH8VKM3do6mq4PLWlscwVvvldB8ONL0k
2KWlFB40SSzMH1plA3FwpxKXmug4QanrHd6+hiUrn2WxWnDWPntynssY97K2JlaHUQhosqutdIk4
nOg7q0gH54QDWTMlpmRWX7kWN+LURZxEO08blFIYOUIgrQr4vTQ7Fb0C+sL9OdtFLtZypFZhknUQ
DQQ//yocYjeeaG5h62BgM/Vf+5FRrP+RasQyZ5oAp5UoF+o4mttdWTsBTeco0A0hstLBproFx+L2
QxnIoFhOoX86gv9LAkvLUtV7kWPo4Iwh7lDp1xIo9zPehSi3EKEvSTMkG4R3ue3p+Wv9TZx9Nuc8
zZWPaQ2e8CsgmPDNAQv9ToeGSIrf/hjFXrrlUDh0z6VmlXVNFI1CTUKgpnRek6kWWxtjRCxNm3eO
O8g5t2xtlUbcQd+ELc6kMvKqftRQobS4BH4nyAgGOxwQGTRAOa+O3xHwZWO1CKZQ4+GLfODZAMXm
t9o0ZUPh4ItjrIuWge4Jio932zOF47V+KW+Gx3N3HkDZgfMoUj+NId5BkOu6Zp7eTrXwJ0c+yu/G
xpS/PGO7In7aWbSWUGDgzTa8EQPSgRe5ja8nFnwbxKupkVXaN624LFXCAv+X3iLGXMNwxX5FkBqY
nSUXRnM7SiYlNBfvcIIaC4oyeMikRB7b9SXVJuJxRZHFmyiAeaiHeYaREiyflUeLzB024TwxgesH
7hRbejZjicLkqG6ET7hHsMcBNXe1+Ic7/619iYp13O+DzSCE394zXGyqWpweCvIIFjr+XH032WeQ
OKruTQJjiBPJjXYxP87+9tBA0n0EApmZ6QJmH6xlHz+y5q9ZCsyGKK9hpGRVj0/3h2Nx6lPnL04/
BBp4+2WvClCkOBkcAeHhfUXUnm+gQ+fOi9H134fGmIX1vKfPAA6F2w18sSHKH/LP+Mc8Dy64k1R8
yWVxtlrMzimtObW6d1MV6pIQljakkXggWH92mYukKOX+cyT3euSeEfVWyGHPDjSpzywnBA5zrP8h
7ehm4I5XctjsW2mwTJdNTqIIFEtICWX9JLN5payhRe6+Oi6jUUOf4dYaJholyajtwSY2887fCTxb
GwJbTxjfYR785O5I2VyZ/6TDujMVFVUFgex272V/W0z2XV867ntWCvSFEoS9dsXRkqbbdxT1pE+r
Kx0YLOL38DiZmcDX43KyQP7ANJBWP8awQUiM03kR+pjdPpG38+5B1E2da19CX4MeEQ2ZNN5ItM3F
ejIPGYJj5BRg58H10EWExK5AF/b0/HS0rhzftur9sFqtawlnIHfqgZmzvup8KWxTnLEw3LaGGeKO
VU7dbWsYoBlAzaRt1W6BWE48zrIG7Rd/dlbuITKo/Os8Oa0X2YqmLuCSm87CIGl73QUq6k9RtgNn
fRn57/V4x/6N0qAI5vXnIsZJZ8P7YQt9D094tvYMLlurmGQy2pphylU3MtH7QQe7KlJdfmPb+aDi
NKKG5Bag2IevTEtvjwL/Zs8+KjpDLZLVDUwQOcSmJicRRXOpgblhidbdedRlTWhwM8C2bvMTBDh3
a5Kdj2CXl8SN0i9+pn5XdEFTyNG+j0nlMr5T9oWj8plULJly9dTLPq+bVPdyonS4a7n9Onh6s3R7
rn/m/0mJ8H1ElAD3iLf8FDEztpSfsoXbq1HJVLO35AoFw1Ty9D4O73y1+EF03Xqtipxm7eyErAUZ
hB8+pLCdXNa9r7N8jO0djdo5pP2dIEhTZV+WRVu3U+58ySr7oTndWhVh3/hIwxTtueZZJ7wJiuCG
unlx1sJfrs7DS40eWal47mY0CNQuns1+0UJ8QGWGgelIsepcFDZqGSs9VyJiTw9qxh2C/BmD3e6e
saN8LZHkaIuPjPvn2vcgNebBZvAeoC2Nj20Z2XgkOEfO8uJ0DVK85lmelNsMMFwzQH0k5qpC1Cwt
Zf+qDnKaSA54YQWfwkYKLfXm3dQlj/RFePFBAYfGykqSMlUz3j7tapC4YCrcIK4AGJ+2+vO1g1aS
DR9H58S8qew9UFWMPnEu4xnIiuhL7fLKEdM1xbVEb8+1qh4Aa0WPgriXeATCDBTG/hSirSkS8UfA
65ls6ieJBnCBhvF6qaxyeRZ63fvOSvK+dYcnGyg2KcqGLxNirsYmi/VTAmzgYZeqqxFYaOO7QJQ0
BBbKS2UhVaQia2Xye1a/Eb6Ll4DQn/bmCEl1PxizGbwiSMMnXOLOUIVLFRUbiiJ7bhwMCCRN7WfF
+Paf+mBDAfSHIwJ2Oto/q2PPUvfhX5YaYz9SpEU8+JVpW4GRDbMWiv6M8J8ktqzUNsPSDrX2mul4
hZWAweC/ebvuBzByP1vaTqnELK2OoQDQDrjQWsWXNlZN2dJO+2Ydfu4rH6MMOxSMGMD73mzsxYiq
od6C56SEF8ofEXQ5UoT60gk3vF30emU33AGIUaN4YxLcEy/hldp1ywKYq3aUsKt06+m5RqLj7OQL
hTkXvqV40Qt1YgX0HSaqncxlQCH4G3Fxu2YBfLkyp50IQOW+TumUWPO7xff/ejE2YKwBn7cL53rH
jt5CYm7We2clKc9IUJKofVuC0TkF4GAqRet0qY/FJt1e8jpB/eNOQmhwgDSioPH4H/yn9Sq8Dyub
YkoWStzi8hz6Q0DYCL6m/HlPD0Pe/Qsq/pEz2asAXtnw3D6aWAFV6AqEk8V3LRAtDD7OL10e8x9A
FgOgpUzbSNV+kUjXrlcHGWcPW2gunwgXqhbDwK3N9JybfWOpc8R4Wn0x/8+FjiyyOq9n+M+3BezX
ar5A4ha2OyeDryPcjAy5gNh25t8LLk0oj0i1ZmZ1JOuEoQc11oc0yhaE61r1VGDdHScqzlEXuNQK
uF83gKowcOhuE0RMJrGwFR4PDzzZDGK06DwKok5uxGAovvVTLN+GO41NydHu55f+vdHudFFfgthk
iknmwON2F9hW5zn85iykjYYN8W//YMChNCy8najM42fIu0x8LljMn06bB2PPb8G8EsLQlbVAa4rD
CHuPWA78dzpKcfbJ+2pkqTWB3sOMTvXMoIIUuHa7ISV6Uxs7HLDDRFznyZa9IWL+6N0Y2OY4hZe1
vWoUnxvtm+zc8CL9dIJiwrliip3hi/p5GQTno99qf+JikOMW+EvQEaTu5QS4gcoTsOijYMi7ukRD
HWyjzRVxO18yIX9FRRakLVdupe/B7YbJgnU1jCyHpBudqa2ZBg2bJvjoat480xAWFA5DX+4rYA+7
puE91GQoHxlz1Sj2ipstlUUjVdHFTt89LWZuQytJbohXxMO1/49injd17CWHE2eQwTjS5BX+5sAE
jNPDnIGYPnIGepS5pDj+Lj+mFhz5/ZQ4tjtj2cAxrz9XG17OBlxv/vG0EOxfWN0eQgprFVP1zSCl
t8kOKMh3BEQqpJanFYDvk+AFgnCW6o11LDzcgQzeWArO/DsJJ8fGEzeQVzbv3Ri+zuicEniOJTIy
lfaN0PVvDsBzNYBGvg8A6yAz1l2AWosXVpBuL6uKP6hBMS/RNdBV53D6pMa0RSh+641c02e/YkQ+
hVfXDYNOL48dF60zLrKgod1VmxQocT59wwIhtvhUsOHcThKiQDoxSpL8ek60NroB0QT2qGyWpUPr
pcghSrp4BioSgj0v/ufXl8FOXpmd7CqGwJ/QBfstpFWs0OmUU6s1VRXRjiOzgk/y9V8+kTwM3yR5
/uUNURcP7wF046lNOyadk8KS8ynDuiqkamfIgKvn3jjxiqGXRH7WGI0zX44WOsMHCzRNgCvtQf2R
85Z4F8tbPBFSMsBQqE6i/zazo0EojztOOWYuA7Uh/81p5jrfzSEH5h5rXn58BgwQmeQL2vJ4qqO6
W87cHa51yegtY21iqIp8sV+ChOk365nawSQxOCout64n8rJPEL0CUkSRFkCynqY0zMYx1WjeHsdL
ygYayZJPlbmxdM1HoAzJEnBj26n/JyKdTr2wvBSPUvgfL9hxdoWhWT6ra4FflI4fx2mT5GSoVhZ3
wiOuu/YDJIHJcx2lq6DZDAc/ux6Tz9uGTQ+4Zqz3E3Ag7LdJCYAI9xAJj8aki6IatW1y3p0Dl3jy
7W0PZm38xNiO340HcEo1h6T2Tr2kd1dffiX3e/9kqVKjRfVikSY4uBADCIjyV+w7iLelxxoXghYJ
NY1+nGf3UDnviXNED0iy/iQ4MaX9vlvfmkpH5urgFnyFz6pe4jrr0vCL6p97TVQE1rw7TAG+cG2f
3n/ZL2R4E6QEzUPfhocYQqk8EQzA4i1aUNutk8+sPeNg0ABROv+ThOPQglfazVWxVxst8gLYbfSH
0TNNwncecVKntnAGgRXBoga4Hy/7itkjdazAWJy/uvRROD329S5iERhvqyyxzItXxdLBb51GEY4o
y3rwZZJL2G7YD+rPcf/Jp3XJfgezEt2gFNLFdWoUQMih4wWAsNSeu8D26Uje5jxXswdpz+ixcHPm
mSxEEaN40/4v0zEzz1LF5ekxrJG/cI5d3a0D+0tZssOwhZts9UuFrUwozJQSCGp3PEBGM7M6zv8e
q9hP+BYweKddPMff5pgpJX9og3+nb5aioe/M6kLd9IzqDT/TLDF7/Pg2/g7zsiMFIqefcfR/4Fi6
RqCo+AjBViMEudpvxPfXrLSFBMXTsvwKa6/pwaLiOoRVASf0msxI6XVoze7ivYoKyJkXtsm7xXGh
jo4bVw+fpWIP+i6xCUT6p7ab/MKz4RCiyplWu90LOgA/a1oakHijUgqq3MyOa4m2v6I6vq3qNen1
TgngMj80cvZolSkbCuesVBNKCJABQgWwt8WERgj5YtF4SOF7guzKLNnRIaGh/yAtsip+DwCW4ufd
LwNc77MTO9DOb5yjIxVEEe1V1b7g/xH//IBoyHgJHfR3Gpk2YswWuoj4I6rprjeBWO5nowJa8NCU
2Y4Ao7a+7Nn25NA+YajUGSy/PCOC7tnKEZRW0jkX0+j3lI1OifLo0fS2+bkeEP9lYEZ0CgFozhoX
tmriDEjtNWiKvpyxD730ZSO1YV19nsczE96lKUW45wd11dVZUu2wzCUoAv5Vni4wwtUujiL27x9p
hUa0sHT3IP+IUPMlKZvlld+cQdARAQCOrjow+VHEl0wXxRbn6rTtWjIzf7gptbvvXsohD7cEUAX+
8Ks0iDpiMRHXNUhk5hn39kWiYXhh0VSzXuEJzsl/cTT14uBifoMg/2enBfR6YwA7cfZaG9LkGWjV
jraVyMFFtYVOqTqb4lb4rn3PpYkSk7EEdPlxl9tY08oJIdr3s6bkZ69rVqrqClRce/uzq5flnLFT
w8MgzCZZJJbtDsxJzhiL4jHN4zNrDE1ybvnv/q4CxBCYC07ZhRtYP6oTrrgjK5SuhVqHdxt6oCN+
DB5oHFPrd16K9w+ee/TGvRZ3ncN4O00RfiMPW726TFNLooyvaJJ3+lwX5rCOsFAhFD4ba0XEotXI
x+uN1MLU1zlFDLHzAzUbeU0v6dX2M9wVmVdmyYVvPDwDYRI2dYyIMtXbCc4IstVUUX01XRkIPv3+
qW9u21iaw7XtGFD8cMqywYJza4tfeD9PWOWEwVatXPMvtbSoBMFzdFXa3i1oMIQqRiq1TMfaRKiS
wCGILuOqjI/QX5oqB1F1DmzwBUeKqqpvPml75OvkjlfZfDwOc5nRpaWAYT9qQhndCvhRcdQ70duV
zziRSlWLPhyOFvEzK0AUng9Nx/GLEjoZxNVsSxeTFWEoe/yIGHqmwlAnMENNCwGr8hnHYl/jSTTr
kifa8cMnxVsx93aFPuQ5Zu35BO1AaLVQwXRN1PJen7ps1CYsMEPhS/6k+NHAYmC02tKYTbeFfow8
lgN4PEHQtAwAZljDeVML8e8zcgOuwT0LK4M8XVE8d5ozyY2SO5VU3QPrtf0H26NQB/nidSrym3pJ
2BXCqp73joDj76MgwQnY7GpATuscnDcLpzkOd4FCIwa03uhTd6lSFy50J3NWa0tqKTBfHMaLdEVn
Vvx4vkfbZQGrizwn9u7rMX3hZsoazF7ZUuHWtqc9lztvlHYIxGMIXUb9KIBTclyg1w/BuDFRfOZb
/cPlW8bsuVmwbBeNEewecE69j7c+KUeBFdUbjD6enGsK9tEeoFWWTRBN8yLo5zJJnJO1q9Y/9xdJ
GpHeNT8QaIRmuZepJHLy98pOHU7Hyz5mPI3NRaAJotyN2kyIszfnWM4aJJO7C3/4Sj6S7i17saBm
9sqEHS1ULkACrSbGec8Io7E58TV67beA92Z6V8YdKUj6BQB/CiPZFNR47XWtUkEWtYiATxs5Zaci
TqQl5w5xRLWsbMQDGu1mXhfo2UdR13UuIL/aBXEpV8A6hTZmop+XjVXliS1LQHPTHhOq/lLk4lL0
3WysJnL16MpI+zzcVDwDeg/8LK5XOfYTlLFI/2gsb9znadao2iGApjIhlzaJRf+1AlKYdMnsyVSP
XAnbc8+tBzlgks2oDpw/fcUQfse2OQ8spt0YIvd1qO2FDDbniK/957jq5gtuONkMJevTWiUkICp+
zrIH+3GaNL3dbDud62smQUwWDbjgEaXBoJMVSeh2PZmf6AlBFMGeeHK+efRHmLKEeKbYFkdIY5Ub
HeU4LwjeuZlO+GuZBIUiChoj3q2lEvQn7SlBhxianfboZWs5FgGLFGT9QFHbAdaTLQ1bGzkbeDT3
nJsiZtsn5CZZkb5XzhtfycBShboJN+GjYFTKZiH8Zq02Ne2ePyXAPkH2RjxR+30lJlUZGEuC8XFM
1Nfgy1/ApvmC0+k/uYVNDEunl+mty2+g0cvlcQK9bdMADTTQv/kRmE+BgPxlLXUrDsMlOwYl3hYj
NVIIdmQj4WnI83Zt71OIxoXwmwy24ZwneVUvSN5UeEsiS352C+6IdxGKuBTPYqxW+m+Vs/u7JRHv
x6ENio5qEfnP5p5fsQpr7mZkQoLQpBGFPaRY8uxPJ008KxdjAKfdOAzaR/5c7xjCr2LTD3xDVgPj
WhkEGRd7j7mvVe59C6RNDFs5m/QWGW/om48eF1jh8zPyu1MfFe6xZa/SLBEJo6uLZmhyfbsvPFZL
UJ1BhgowWWMSeC4AaX4AyxUO1IEqcY/+RMQTuk8IgENPectV2+0PsMpQktmc600plwrT1hLTC5Zv
Z/CuCudD+OczfsEXkLMyVWimfftvCjVcnUyaTeuCG0nKUKz1xWBpGKbIqfSYLT2QudS5+MIzj8mH
FMVaItsXMRSJxKDyEHTlpkqX/LUZ3/fu1m5gcLiSjHrdlrWWoupaH4dWHO+f1yepdr/kAYpRGKXl
2xBZdExuB4/xq6/SF7qG0GlKU3v75QAUqsbrDQmWTzOMC/9kDVspzPNbWNp/gW9ZTgLWDXdV73BH
Gzlf5xNy2SfKNKUtA9gGheTRefjS6AyFu4II4Z8XqmU8ceYOWLEIIgl+dPYq2I2W2zLC7Ikfeyaf
aiRLpU8SKO3a7BwgyyXW2Dl7ZKlETc10pnstOQN/fmn+ZDltKYJ91+IfNnyBFE1p84XSP+A7JANd
0vMw614pyLHbJ2hoEXb4twmVQTQr3TooYurLpuadf5EbIobrcPQOjK00+suFM9IdhMv7H9zfage4
7lJjvkZv52UmiWIo5mHsloHEQk9Px5K6BC2MEqngCGEnu4JiXVl4CzjAsKRRC6GCoWFYs4/QYTC8
5MxE406WrZn439MH/dvG1MY6UU6NzzeyEwjdO0xVxOEgx4s57xYMUHktMSkWBw4drLo45YgYQDSV
KNullYBkIj5MRDuZmz2E8d8Si9zat7jtpAYgZI/C8qaeWIv68BWKDAfR/DNPTfFHg8u3A9tb1bUM
xv///YzKYIYPOT+yicq2jp69zWudMJ11UXiHpZuMRZV1zBepbQe7IKtUz9xBLdrtPSsnM93+oqZA
Dr/6gkrT8pzkRwxI/KzdOrUSQMoLngvkZ6y/l1hPMHtDs3OeOj9rN1QAXqQEjCde5TsZT8Ks96qv
FXgwQglTJyfQaaVW7Nn8Iyw0R0giQz0f5Bzh71fPnkM2/kcbkd0h4zyk+v3WtSa8OiKsjC2iPuRy
zTn5S4zIy2kW7pVt2A0n0ceXY4lH7yRYqofYbZX5t1l63O9Kg7JE6PujvQP6YOJ/j+XCrNYqMKyB
RBHYCbrO5DWgTvs00i47wR4iqyzIcwDMsinI/nJUIRwHxaZdTrhr00+VGnz18MdwAUL1sVsA3r4y
pjMu6dWjQFnogR1fxMt8YTjRIAG/y9uN/NfocqhgJ2DKlOYwnGaJo8P9UaLhL9e19sKFvy9+dM/w
6H0UM/nnQZLcrnWnX0WISljtkK2moHNc6PmVdGXW+KQklegT1+qXEbqfFJDSOBFkQh754iHORy0q
EZ61MFT8UyYBVmytFmwURPcNt10zlK62ssWnU5wPS5cvrh9jrlyOgjVUPz5H2inxdWbnv6NGD42J
A5Ah8Q9PJwh3Uz1cHPjPktw8yH1DvttTbQxfRO6kF+ygJNkH+lCdfc9Gb8HCvPF7+8WSP2a7LP3A
lxtRAaF/uStMNkAJ2RVgrSs44MxmTXbL94ZixL66dJcKXUkkUqnEMTs2H1x0lIJ1cBRZSz0iqWwT
hoAzXGNGkfw9SOcWsGzzDOlMmlGcgIx7Rg/IaoigsszEFyPJeQx7Kfi24/EpaqRdcCu+i+k7Riiq
+fbiUO8PKwDPPSrE5EJRo1dncLb+wHhuSv+lZQCg1Knol66a0lfJCvBU51JuCMVWjKVZ1cqSd4ph
4Of84D3sjkpumH777v9gviqZ3aWl4rFkeMBP/adK+/KZaxI1DWU+l9hom2Xj080i2tSZ9wQUKCRA
i8KbAxkcSsccOOjpl4NLZ9ii+fAKyLoAiorOMWFHb2CPmb4oq3+m7Z8UKL+BCV/K0T7K3PynPZTv
CsY+D5d56KlhN016AIearqSJJ5iQ9Hr/wGlUEmxMI/nI408/A1TJlUzTnLPNATINRGxNR0MzT1l4
TlYJg111iRK3mO5hC/Utev1/u+jhoKJMfc9aqFYas5qelNZgHrjtLZIhY0my6u7peCWEG3swyQL+
88BD5oVUYwcK29X+37k3RKQhgX17weSu+6T0vcCquIXJ5212fBRr2LmxWtzbb5DoKkUqmd7157cy
PLoAPnZFbjSOpeq7vjvYYUVoBX7TjD9z4+XecaxKv3EfwFeDYx9tEgFkEPpw+0sw/xgDu0XNnxnA
iEB2krVUUjhhVjbb5wqq6RfUtVw2Iz8T4xECDBatnqg9b+i7FshD7t+lPzRSFESY/n+X0yotpspk
hJc5gIFc0gFaXqJXMasxLk4/No2B+VxA+SUy2S67WueaZfQOBGC4Oss9t9bPKUXCuLbIkghwO3Ec
n9cYB+GF30rWVvaTZbLpgaHCWc4HH/a4ZCJNvmw3dA85gKZ55FGoN9rLacug2h8Rafnn92fpYH42
zcWHcwfqq0o/WX7sOG6CNoyX1ECdAOwx2XQnhNQoDMt5HxyJjryPWLUUQirN6m6gvF0+XS5dqXh0
LdMYRlqNrzViWcBOFboW1PUnAjZOPtPrfUS6/nnIc0d6t2jTq0QJWfKI2Sv4V30BbZUnwgncD+PJ
vQWQZKLLxXnLHMCGU8pr88MN1GV5nA3ikLfXYiu4U4K7kiJJz9Zz9yS4PF771VmmWNahqetObZJf
Ty6ny/OCaVaHToCwkbeR4YFpjBDhK6v8GefViNw8lICHY2R61EJzUWnKZqK/jPJUMALSeHlEnPm2
n3Q1t9kURWc0TA9T4YMrv2G8c3e6wHKEaZ1nxTakakOb/8lBaTZS0/+XSewfv7IEkWRPUFnWuFST
K/qZDv/pqqCjql48L8qPVp8zeNci1xo2Ao/sN4hRULZZPSrAiuLJ3gy9oSY798APHEb2Mpd0plfe
URqT1d3KltNAKmlZLA37UwsVzzvFU5/IUY24DMeI1f9ejez7OEaXwdbLIoLL5ewGR2gIDxyZi1qp
VwQnXOb7V2Of8nvkVLQLJljJIGxX5u53leQfsfIf1dkN2U5cnr8/svEk8JsEvvh7Uz/8rXHQI4G7
o52y0aymKuuFA+dvV+qQfjamYb9tawUteqTq65iD7SPWhFHkSTp2R77BUsiK4hGCg2B86B0tnUdz
SonURACIQqHgSoSIBpbBXBBZf95wAP7Bjtz4qVfPYk3htTJyymB+v8o4iaYL9723JOiuFOB+Sx+z
P82BpBg33B9Wk7eiB5913ZxSyRnzXfvwXCCQvvqgv6SOqb+JZSjPPz0zTbRRMQQD19i9jAcvftFs
jhFuxhpKJt7pyipZ3GSr+QdTaMngmihz+FyTZX5qvFffy9pbyjroL32OhNpYh8WW7ve2UHNwBKDQ
bYTHDM7d1/K9A4O8VIm413LHXeMPzRZQZ0cUy9z6/PYd+HE1XZ5Ek0NAcyhn0o+EpCx/9esqNBTn
XkN4aA5wtAEHAah0olbRamG/AOM8tMX0FIDTUT3pJ1SNl+7OMbvQsWYRBjatXhAIU4iJkm9UODlA
1WLdBQtBen6kpaTxxHBSmq6WIOYDSU95wz8hg0bSxRS9RMCq0WDzYmWX4OQ4kwea2rFSXZ494HsW
DLV5865yLpavtlQZEhm91Fi4Hom1dUUyGKAt01QfvCOSbz2KVvDlOeSfrF6LjI5g23Hu+wWZ9wiu
v381db43P5yEuvHYdB8YTdxmsob3oGlj4cYTHpZU2DTml8azW4NSgSRfhZXmLEAHa+FgELPHQdBU
hzoof32LuZha+tYQwxc3khTLn6Rr3QSWBBmdRrnxm2m7yox2oPYOtXsF4Nx5EYqRFlonILB8Czfu
esH2qJkLhIbaBwmogDHwg2oEPTRL9o76VEYYIgjTh+hwc0H2itSlg8toPtlpmK/1kutAWYyfTF4L
x22IkpsRaGx2pqzhBmsMUNEmErG5/sFWBaMXn6P/bEaOn8Y23lhR7V6fKgLCxUFYmEUUgw3dkTP6
TwrfrJ6DBrwEO1V0ZMoTdUWc4CsaKwCGBdCEBZ7pnG4+yiM2MJt6En4I+nA7IWC0Z+aN7Ej6grBd
142UHO8WZoBuCLFERVKiG7erz9QoQq+DpjTK9i74vvq7hmztV6r0NjBXD1MIuzH18BlDec4LUN7g
qoKvtF/O1FY7/rYllJ5LYbJyqXnWk7Q/MKZ9MHSYD6y85dbcgofZXLILsu3xnyrFD8q7neFgFLb1
BBIiTQodr85+ZlNyWZkrKK9Gb1NQf93kLrLU6fDV/Bm53Dza7R4kSUCOvHq4z0K4vNlea79rw6qA
5o8xLTkBRWfb8TRV6CbyWhkaRsKpJCulDf0PCEhQ6vZDH0ZxAvF4fVCUsSuVUEFnSIl7T3kFnoSi
J71vt4VcolAt3KzDtY0dmCeaB0tVacB1WTkwQS0Y5Nnaf5877PhkvGrtaleZhZIXB+/n7HfYTp8F
f1cNXcag6i7n07BGrnebJfIKXh7bTzxcBGbzyB27VfLhISD83u7Qf9wZOvaIDIBJNSIvQEBiR8Xh
KIugvqqSF/DNZ1Yn2HXTNKWkNm7YTZ83uJxmE2wPtfLB8+JvIhSxFOH0739nZhJX2tNM32l0ykFr
TiPqMKr7j4ZM+zGzBhNpbgmPRBQ4NX/2ma44bkb5ZGxq4O9+SoBy9ksLUJwU+8b4hGhR33zeQnZm
tLGdPK6A928DUR5/gwQQKuCUqaIR4EzEP41m8lqwKPTGJjfg1XPr8e2I+pySEO2/dQYNiqfTWTxt
h7R+oM/94oOjxhd5EkFY27FVb4TThXO0wEJgGMwkVQCqeIdgk2SmneTIkxarNIcQNf6JgMGmEXhG
Yaae7vNQ2PNJKhdcPTb3aBAx9aM3xWM8JJ8hwriHLn/gU9QZjJX7VoOANmtq/9n1HRY1lUPempEE
fMUqzxkcwi3ONMs8VoStf8wAZHF3325YfplF0faKC1d/yQtWwkFED9uHfnR0SwrOt4dWDYuuDrBT
HcaluAjjEs2Ynm82I8BGn6Z4a5mBZSyLmT/J1Ilp5odIhYkLYFxIpQpXOUtGO67UEuNndbCtQJsJ
0mh98xeAiFernXvD8K+lI/zG7+OH6vb54DJ7jnp6V9tTB9tV5hUzH5GRbJ9dyjHPzeN57F1zeSpl
ukuOGr+BQty6rsEfPllfgvPwxCR7D42EHFSLUrYe8xgTiZ5ZxPX1M+XibtqD/4MRLTi+yJpYEb/V
goKoNE1/DHtb+PAwvhqtYgthEdOj+1QQvdC5J9wtQxl7RNxF+Z9pGQJw9nSsYV7TN35jDIiBJ48X
gfJWA09i1SpM+AWEMym/cyi426k5Sohhsu10Itfu3OmDF37E+dBDnRZpG4iOkfoNSZZFwMOefvLq
MQIXlpZPjee+0IVIS1+lBKgnTv1PTJClXMqiq18aBNYoG1j9AGpA9f8bX9MaQ+DDMhQuoGQvQSO1
CeHvoIONiN2cWcFlEwPa7idJtdg84EiZx3Gi5tehi1luSS+mjirWiCUsonSEnXZLX9a7r56kuiC+
CLqBD0IMM2cuizmeZUHxs/MuH0yms3d3TAnm+6VHNFQlwX00yrkeujXewoIHIhWdwOnZNHCXnPOu
3lol/mXdiqVRhs91a9fFOLFaA4Mqxllb4JfPMRhivRuXhZO54r9yr3gY9YfmMnmT2jg7b/fqoOsx
ChsMqP50F58uiVzeogiytoqSzZrBbkGTQtX5OwtZHURqKQBX56I4PTSSPK0JNhNlX0vLs3pXPH8B
8ACT4umqKCMbMdSa8YGiE1ZqMEJ0RfnrU55jsaoLe1MA8LpxWOEmszebuyxJm9v5OevpVm9zO6Qr
HNEBUbmKudsk4g8QqDm/9qfoQ91TVDxCKY/RhzTENkJWGvE3fPCflts7O+6fqoCps7HinSumqAWj
HwR2S6Ee7mk/iPJlKmadMznhTG1Mr3x3vaAHJW4OSxuPfrgQtG0xJAe2fK32HjqcdJfRbVZQdLgE
0t7MgsgnvLiJ9IxXGJ5XF2qkHGKi3iihf+27Ut8aEQTRHdJcFGPBqlbmPFfnoZnw+8iK9Spa6ivr
u1VlmIexszhP0tBq6ur4aBcLw7x/ut4Wc/ZvSj/CszsrmYPaH6u81Cq9sjyEFO/YCrwZX2/X8YFe
GP2ubaeNk4g3Jb2InsTgn9+3Nt5y1Tt+MV5FEyfZkOea6qalbTkj/EINHE0KUBFcr9UNH9V4VdNs
AZwKkN5EWDsu0Kt/TeLdHvS82/cS8lz9YCRHJNzCEl+O4kV3GofN5I+SGT8CFQBBgbvUuMKVCDPW
NZLWyClnbDcVGl7X+zujRg4ccdbhdY65xrA49ept3vtDBdDHE+o37hlsWyFsUD1pv2JfwGJreIe7
5GAS3hPElnyOFiGUDdHXYYBTCPhSS8O5oDh8T6GQvnHWNpCJr1l/CS56uYYhxSkbxB7Cl7nCmNcm
LjqfU/9lwCJGh/ORx8ymuHXC+4VTcbexY2L8ri3E0aVXket+qgCf4CfHGfuhPE5nGizgL4BRj93h
3whl8yuGcXPMR7b6CnftlbnQyKL0KDb6GSVK0zg6DMUMyIwdGmRnJ6DmC0Phlb0/mO7knpqZ/9gA
2tebpzmZO3DC6DXYyM9HgPLB860ncg+UctNCCUlutrthQjtwuZvIH7rO3ol+zLnEuLMZrTiaoyAk
Vlhmm5TtXD0V9I1hyojm5rgv8ZoXu19GGxvT6UWIIesuscuoELrWio98nBXU/AgJKq/UZfg5q3vp
h63i+Ep0cQoic+B6qDlr1XkIv2ZmnyfACQ+W05Ko0Z13oIVEPkA6fs4hNeevPv6IjM0NS3XVaM7a
OaUJ2eyn+oZD4re0zWRhEO2uue2AkmJU36qbVysrlyMFTDrw2o++kWJZ93a0dot7/TYUu/vPp1BN
14bSKj+LBoqPOp04J0pDlqEo4dojbRbYUmCPK5HEvA0nuGXG+K+A+TMagUwQ9xPcHIGobcG8/G5q
HVc6LclezitU788ItoQutr2cG1SsuLGciG5zoXTy4lClZY42v1EGXFMSnfaL9ywfOtjR6/2uzG3R
j8IEZAm8bLNwNw9l2inHMrVuq1A/arZzDOW2YwfJoe1BexvRanx2jddfd0U2nVpzLa7qsSzf7OCm
gAN1XGrtlspmv5QHys9BHd2hr/TXP6F75t33UGMsXEwNUlThj6glaS2zlCc3UQYbZHZ/9s+vJ/UQ
/1DF41100/HnQ8V4ZXqVxIzya/6ZIpdDhnkPEkHXOk/O2fK2UOWBtHj+fJBBRoxbtVdAnHrCow8v
Ov6l8/LG8iejQmtqM6CV+vRw2r5swy+vGmkzkWzSjKuxKLZ6XjZqzr6/vtQUg51FlUiV7wYX8UZs
kDJJ+EkYkhMEH0n4po1oUxJX3CuHHNw4Z1HlmoIu6GIShNcJA/vbBSk+puOjH/SHMskAX1nbXk41
rAeHIGgmJHiMHhZFv5QAKvdiNpqxTUX8oAvItHgEWlaBgmbeWMGg+PObUWspkbaIxTsPdQIqgeBg
wUl1ZNjOBZtgQS1wZrkGjUdNcpm6Afklrq2ZQIJqFAUO32wB47QYbVl3SN6gW7RXV3OsbjgIBk4j
H8BIi/Z1U++DwOK8fXxyuRYxGNKol3ip8EoUd6XYyMUapcJy0gVDZwRIP4DKHsVei25oS5Relka5
tdhbGMDIUg85arQ1hQeuLhfuo3Rzkdpx/j4e9eofSYvXgyPkPN/FliJ/FzO3wNE69O+wjOu8MtGf
nzY0WTTylBAMOPFIHR6roqG7FydOktOIKrdmA8nLP1X/9A6C31eZswL2btMrjE6bBUWOl9PvMKPZ
eNgIOXY4gELJPnaM/8HPcWXlzVuuYl27DaruFhhS2eMoOmMkxyOBgVl9XLce9toZPpC6K3+z86k1
pbV1oW97vY8tOxcR7wf5QFpv91apD6+JMvoNlbSaPZALdBWYw8MWPoF68O5/J+su9uFH0nfmaPH1
Y44TpyW5dOCIr5qTi9F9C22v+zZHiMwowOzpvMzn2ffRFxrworapKD7meLSME4Bdr1XHn1ApDUk6
noKiUCV+Quegrrjf8zNM1yvQGZ3Rt7BJZRzoCLWCwHqKVyihHQmBfFAr6YY7W+yAmFWzdbpmGn5s
MzO3o57TP+vX0pzumCVpqmnjCi4BzIOyxGmMPrCvw7hdnMngfTugtPq3EdIqoTEvVLH+MiFJgHwg
o3x74nBP/wwxrtK1NU0Cb+MgW6MhLPSd8M9HmzsnEzt6vdXIOvFpWUhAMyDx7lHIHSXG45rwqcM+
7sBk8HuHQ+/232axsfuwAhtZ9mUmQPslHnfOJEwFBKFGN8sY5ucDpE3HXP6ZwvTpwa0F3I4GWXUi
0Qc84+/IbiCKiVAb6G+lcnhBNNsRGJUO+g47D98ti/3BDNEUD/wjx1krKTUX3PmQs61egjjxF7yp
buNSnc5HDBCv0EzTIxoJYKR1a7u+WGGSfeIwvsvCfrNAYgHWQ4xurbJh4wEFMjsFjTHSfLoJWQiB
LvGVib7HiagN+zOQlb0sDiXbUZNStJ65ZnM0+XJ3zuoh7JUKSSdew9Y1TNd0pOvN/aqu3DkihKTp
FeK304YwjuCrBDhdo7I2Bnp/av3rzt4hC5qNYyxscHUKapfeSEy7NnYp2i3f6xJOgZHGqNZ9RU8T
OQDWd72oOV3NIlgeS/BKMfZ1TvXAgNpxObQL4F+FOv+FxUNr5GB35QOk3ivplNX2AYCQQNiUGPez
piZNmHB/+r/at+xK7xwx+Wxv/cXFAcP+6WQ40d+CEeSAAxyzBnM0YgnO8+yg7//CBRCvyWooJxbF
vdgFZn1BJdsGxtA/cBttKzs4FJ+OM6bZbU6LrVcAAx/A0Vvz287qgIPqIP5Gcb3YJ5KY18NsZnBI
MkC9jkLosKhfznDGjJiXHS0i6MZ+1m9C8JzLipmMpPW9oeiPQFJGvYndHYHkhOWzkpUPrttgybci
Q2pQlZAD3PddYod+yH5OZk14Hu1w7jx/Ku7XTTN+KHS0WetyY37xrRjj98j6VvzQB3aEbbT14B0J
iZKL+JX5d4POb3v1YgvoZ2MjgYrnaEHPXDZXz4NIqyM4IHU9+Qg55AJVJtVcAGZIuPrMrzyEOCoz
wdQHJSq1FfJIwPUiBwcE6K01CPrP24/f44gNM54loxUbkWszhN2xuuWfZpygbvRYQK1fS6agf5EL
9TSWrbzlTS14l6Tajyukqffvn3Y0ui3pQgW4YdisSP2HOkhbtlwSzoPDdsR9XoUz914puPAtK65Q
TTXxQV7d7hhxOIUytMDqFx8bu1P4Ti2JsXlNug3TfScJKnnJ3bBDBoc81xpWm1SDfI5Y8/kS6Cqf
hrOWDybGx1NUjfARMQpSyF3b4a43lG+KhYLjZn8FKRNynLdrTLS5rEZAMEC+tr4uRmb24823jWGp
9a5oVyAizJANYsPhTQ7Pn+BomMXIrIycb3QYAxymXxXqXCEV+zvFLNFZncI5gyirrML1mUKf7j9s
zSXvcsf2MO+vbFXsm6xIKI8Ud2/FtkFaTnLVn88nPC9DLkwd4MRyovlwbgLV88cT3QwYWkm2w45B
o7xVzxYlIbmQE55X1PAGCbG0lnIYy6IXNFQlymL+DMLO8ujWCdyy9rdFkOKZWNJj2UI25Gv1RlpS
hZ+Pm/Rgeflu8KlCDjLFk1W4vV11xyK4WRjNyVtD8PyL9Pet3fvgkSes7rDs5vQYyhz/ZUOJMbKm
+wLWC3T4kWWb/W/xOxQrM7U6683IXJZIl4KLbPINeCb4+cUxhcbH5WWqHYcjTC5GnIWUjOhIdXVL
bbDUktbADYm3gu9ljbqd4M6djHGj86Jh5oC1jRTZwxqTwGaoXfyInQu20HGHHWQfrcPeVYQUYZfL
DK3iJP/KenEaKvQlTk0WhY0sSnVPUwBRtYeoWMAgZgttzeX8E1Yf16g4hQ6BYrIDkmNwIpppG9oR
I6EHAYLoSZTpPzKiqjJ9RKWMG4feOrHGDzmbagGKtgIbLLdE/gu04vH25tr4ljBVQHKdf+e5/UVq
Wh4YJu9qXwE0hLL+I5iy5cOT7mCp5BR1b40ffWZbYTPTfhCspd1xipgi8QQKkXtBwutSrZaNo3LV
nZVokQkwAt5pAmbxJqe5phZ242An1+gTEwVxg+l18r88s6bSJ24jPhvV+ipdLa9DgbuHM32TL7Wg
qPOirT3yvFBf7FY2nYZEjVOCznU85+O4lvGdSNtW0GFdtgPEGpco3hiaifROc42TFYtSgO5jxC90
luB7x2I5zSlg9jVcs3ZduO5WPgr2dn+kVrtvU8Rsc54isdvrave+mLNl19cqZ7urtfPO0MECQYL/
x3DB0yR0+xd5Q/StyWa6JQZmV/YvXirwQO7hqLXZQme5AAF1ID+GW9sxMUHVNR3A9sRCu9CMzveh
/uDHcPKXUApTUM+ZTSQfwQ2v0/w7GFZYxygzc29Ovy7sEx1gtwgCm6oT0IF80z2a2Gl6/T7ll32d
tlE15wPlTpbFjQ77gIjO7mjPaVhnrlk8T99o3z/snaNpE8DRjzDQ1CdWV8vSneX64zDwSqU5KlYl
TFIEsZ3eMOZpWMzq3gBSBVc2wD1DkXgfGC5FksqlqbOzXZ4w+xD68F8hFvGGRjgd7LjlYE1WDBTi
p4LbaEjit3/SPefJxalQv8fn9ZukDckvuzl9z9fc2B6J3KBe5RFejg6ImbXsVGLiTmapeKxFRxHs
4ZgPTVmogBbtgrrIGyB8iNyXtns/lAYe9y3ZvNMXQHT/fWYhay1bOu+2iRhIC5Tm9pBctG84oHr6
POeRRbWowKNeYHHx6TBrIWCb2k0uT7Lb1lyouTXM49PGOb/QJZSQfbFAAI7S0Nhq1WBAVdY3+YRD
yN93AWIAc/XZBI+qT35XsQp+LCIF0TNo6QYmcxW0E2oZ5QybL9YzsqO8noB2uuWve3jMuaoCXrbm
U3E32nVmXcnIsp+MyUGeL0bofWYI7U5huJDL8mSiFvH6fCkBPWRxJ5xjFszJUDPI4QVk6k16ZuAX
sA7ya2BZ3MjbhebKN8xsbZBDSEl38OMbi11cU+s/7vDjDS6b9wLs29r2we0VbHiLp3Qp01GxEXb7
5pS7BmPR5oFgx4X+GfuYXsh+5KjBC8azcz5/Yf2ps62Ptezq0Ox6slTW1hFAryxhLEFgEdM0b21U
aRtbAnKJNecuSndQukRHntKI6i6w5eRNV6Qp7WPqIjyH48c2bteLMnNPqW+LiAZrDesoZFD2ASYf
XEUAqs2m4ImLgHSbjQm+GVupQ/rs1XA1rv0+nPaRHO3yjixQarR+cYyHAflmZSNb8gFHK3V9drUm
owQSZwFjTHIYQGe9DTUPo4JE2LQ+HYKuHAk74LDEzbtTxFib36sNquHlux87XgU2CFzfpp+ZeQ25
s5Yn72xCbgjrzk5oxxjRod6GPE1fg4tl2sbvggcO9aTzW7mYm89MvjeII+XGoK2nAARbucO/9kVH
p45yTrBQfvMh8UVSaHCS57aQkb1JSH2Rmx6uPj7kzoOnJMLQ4XXscRjwIIIP2L/L8pbTjrDAGxRx
HkYpALxq+Pel+AIfCzImkBB3HXYlYOsJG77ByD8D43YOOincRct1nkpT6PD/QbDINDZ6guMcZeW4
U8AerdCtrJz0LaUBNE4fo+C3K0dzJuhcPT+tPWHNC7K4qnMt0bKIRkp9zdDciUXMMs+jd8o36OPm
XjhvS4Kz2v6rLI9vBIfMYaCEGAOYXqLQMa+Acg8LomzCO0mB89EHgq0CKSFqKfs/VSPg0gp67Yg+
Pp0b3rrN4T88FN8Jk7Dq8o0At9kBGb+jwYTFAVjRC55OlQVHf7MNHV/M5i5OlQWJlHoaBhdkPjYG
oOTNdshFXgjc4X/ORk0fgXYwJtc9tpUfDqcH1J1JO7QlLDAndiCfozC2d+3OjKpaQ82cCNimQDnp
zbKX57GLm0NaENaRKMiAVmjD3/0qBAp+XhcrdnHxY83EzxpQlFiSzggp4AmCqCDo8D3v6RHDttJS
149eVunm0Q9tjBMK0Cc8OQUdF/29+VMHwznsb6zox3NPlGFwF/XPp5MjLvAmz1zYkMoph4s+QIAH
DzqoAPxFHUIOVPMjkI8Ju96AcD4BKATNVb8C3w+Fv2ydvks8UoaDTdc34arBbRTNiJK1uozXSxsY
8O+wB8SgcUrC3wm4Ni+iaVnpKBWO/aB2VVdZK7XdM8lJV6o2hWdTlSJKCWiWqarCmM1gUr0B5F7R
zmTIwkHmun7Bj5W9a2DyzxnILWa98Tcv5tfONS36nIfU8ltnYAgB7XcYsS3Un+ibSlUDa4JMFkED
lyyvleiNlTt7BTZnJqG3asLe2RdZt6McCDXHKtUOyVjQlTLOI3etl0Bwu92r7PYUIuBtAh/hUGAA
h3+PYsk0c4Xx4x2l93wqMk3M9lRmEjwCdzhRv0KNngMKr4NF2pRtXcl3AzyJfI9VwJwFw6217UYp
hCGah01QdN6liko9Uiq+nENuLJ30tJQItuPfSBXokjw6L71r4MJmZWVxkvqFPP3/8XQAwSGNRAam
Rr+uYsHlb4zakzPPiFoj4lF3J9tBJYaPrN6s7drIyKBJKR/ll+80TdgBdpFOIUOT6ZttVZSqKnMv
e9GWeBplC7C3C2SllEx1T1MAB7bkV8ZiwSPiicO/y2DWzK0v7pYwylnZOB+FeeSEI5kwnjrnn3aw
n/iqKnUGHFShNQOZ9D/F/+WUAtU0a5Js2Npdb/Vw1BMKQm1VAU+inSEQbcT2+yvT0BBnrQ1pDQfv
XsLnINW2tol6QJs/jQMdgOqiUvr4caYtDfS6ryzItPCPU/scZHKZT7RtDkQw0XKtrg16NFtaB7v5
kkZ0XXB2pchV97qbjRTxaPJRPpDU72IhxHKe9+DJu7Qr6A7DU1Y/hDpjQAu9hB3mtCaLymNx0Tbs
pqU0d3RL5mC14pUzbvLgvONfjnyExG/lhPEXn8YE6AEBx7sHMqlqBTnzePTOKjz0ip5vTPl4bVn+
M0RiPWJVZL/9+K6Z2XIRK4qtRqXoERbu36SBDUlnYLt7RM5arZng0rxyCCOvr+vZgT4SbYRZn1bU
yuUlM3R8z7gVWdilipRYu9oWyGtFjiq/0Oqr04o8v4PAeMsLDxQX/r31Jptw9H547Qr0CT5OrzaQ
VIQYBC6ZhfG0Ch0C9BnwzWr394PfNlV7U9P0PlbfNpB8ge9R1wV0AWfn5zlChHuYBWbiOto6Fiaj
rsK9k1a5InKTjy9Iv4hBvDdRPdC+XXr5AGnSNykqafo3QgzrTFWojZ/9clk+/W0DF+Ph+vsAi+Em
WbDzGI6P17Ak8g7tgLHGPXm8W2fQpN1u6DVYpiAoBC4xpjNb5qYfCz+eKSVPAgLIJvPHKzPWutet
lgY7WH9UEBsFreLGqZjOOE1N55StTa8KGzUrToHvKRz8MY6eEqd7D8m1Ri5HZ2OJf/k+skSU468N
lWhPvvsDKLr93QnGltonOveeMtGM3YLGUoofTMMvRvjgu9KM4nDjCayJfbUeIg2EfT4upbIMpj0o
9k/nI5Cv/8tzhR5sYWXQLyfa/DbwQYF9hR/lFpideZj9/V8qJDbpPBvIxlzTKy1oklb4IrRST/br
Lh+Zh0e3ESTDVy8FcL0xP9Hu1Wm6p1Ms3PAytPZcpiYg9peALkhJNU/RLwM2+w43pQtp9vIsc3dr
0564Yihna1cNFR97duR5QQI4qF17FMjds8xt2pgk0UMESlXChy7nZqa/9yqnZPdSOvO0jfmPnuOJ
EowPCO6pM0+Jw6j2QYhzbfRXo58Duz4i888A+4VukzcrZKfsiIeSO76xXhG9C703T9o0oUUCrk8A
CgmDWQmlDPka2vADpRkW5nHF7VoFQ/8YUT61n+FNtNHV0Nv5ciDf082asNvAlTyKY8tZaztIVml2
CKN3gN0mQaIhxAhvrwXtK6+jXHOU1ecoVN6jrCmSzpk7tM5eQ+VncksPvDl7+/FNmHY5UNls6685
Dr9+moC60bM7fpKUghZW8hg693Hjqa9s8IdK/2eFn4YdFuI02X85Y5daWdNQhVs3YhGx0UFQM/1a
xvvOrhtTtDTh0jHbdnqDDoQFuk4XDZTXNZQ8bLOb4GONo5k3zAr1y7wnz1NGGJKrO0P5U3n2TmuY
6FguWFHK/mty36B5vMnSnE2tkFNbwWm8W+5hDAHWV0D0asPeq50SBcx1SsbWUjagQg9GSQAFPa0m
GXywonVhNahgyG+JqkG1LioNa9xnCeJ9lpwYKSFmmW0POCIKUz8yQx3B9AWR4GbsUB2/SZ/Bsgd0
fJ252Lf7mmHGGlKHeOccKxoX/cjpt3q1G3VX97wJ2BW4EZE5mI+7Si/MHS9nz174rxWN9IbNRRPg
HeygOkPCdKDmJvKC7iSVbyiCz8UCmR/xgR6YDpkq3Y/XxorqXD+G4Bitacy4zYLpCWw9nbEcho4C
OHtLnklel2t9lJFoFmHzfjV/OEf7Ia7bDl3mJdEjvYecQyBuG4vVdChg9v9WN9HTHM+gUk/xg14R
GExpiDJwjWQaIC9e0NlZr8VIhkNBu/jx5kxeB7pqgLOOQLGq9onoZA5Xz6ejnvtGf7TraCe28Ijx
vLsET+3Mx8C5bn+hNkmTpaaRE3b41AtB8HO64EBZESwCuGoTaODAXgEhLbjW0RKTTVqVDNDg3u2h
bsyyH4HMdIMcktkWt1ImegHO7+32cJPCr5oXubvLa1uPEAeKr9Mvp11GZc+XvimZE0z2rc18qBek
6/O/dvRHTikQjpsuPvW+6t9MO9L9x9P2Rb8Z4GY6OrGydjDzrVEv/NFQhgE5U+Z7qrpD2DF+7osz
Je1crMygE5fg/u0sCFZyaFC3U+hHWUrfAlDfsdhf6AN5LG5IatIuXKllFNFFst3KJLw0WfhdzN7K
cJwKJ9syW4SezdqLet3Am7f0ylDLcaWYI97Yc/XWv4prbzNZyYy3v9pDfE4dI+F4jNeGa9RsPLlg
PsYTJ6B/GfJ4dVGzXUkdj0+GE3SL0WkYYOrcJs9CTQR5kQPK3ZK8I/c3iqjglv8/l+nHLHnaGCJW
csDzHtsvkfL5sWhN46zuRfHmFlQiayiaedcMFZGXvmICuicee7mfsH+FiOLyaOKwkP+bde8p633U
HQVOAbRybOGIDF67DWvE0fQvQ+f5B/jZsVlIfvAZAoRTzse+NR8ZuWiMsEfuS3L4Aetw2o64Qz9B
nMrhK17G7q479d600tjlaGIpy7ZQN7bveiHyxbBVlB7eh66JRJRmND2nU/VpkYN0oJaLgHBHxr1h
mr4f4s5GEQC7P0NqlAIKb9A0bV3A56PN7+ij/sJj3fiOqZI1SVpethQ76QXYdYYxCHxonJjeu3s6
5sfA9YMBaLfD+ud1zCIDL5QGcZf+F9bEBX0nRk81wxhaqhucQENDg62i3AGEhL9Vxd2cvCv50kEw
ISXNinYR1P3/iSCZQqR5oslHjuwdVVjZqQobbgAbdJwtPNWlcQ0GkqwsCpSyVG4ug93Bdh9CcJ19
gJZQeCFPmWpwdG5NWaC4KT1OJsmZePr4jXIcGheX6NEIaMVisDrEFH1D68704er7kdWfJOuysTvD
S/NBOG480d8L5wwgkxTDOFyVZuA9spMIn82lTuj7VseS3yXCeWZhYKaFH17AFsI7oA3t4lPFMjo8
S+pLUqsobZ8D1wHNprIuMqNRKgh8yAN056cammJwXDX8sNtHslbf4uOqHDyZVP4xTuQGOQ/rZzde
5nuCu4qnCdFpNMHQ57zl2bCtdlqlAB3IGkZ5idHGUA58/AKNxju2SZqCSfb/+xkP1ZQkapdaUHmj
6KL+qECRLSiAF48k8y/YBNAKS2VTcekGucg7d9pB2PsOJcyB/TkcSDIMfQr4djIxvsvjO5iPQCn1
gpXJmSjgGIXwLy3AzToxmdQyTOskhgqu3zEqNRKCSGv0IWUXSdyvqGuYtfiYQvKdnSV6Dn4GpDmW
2MyiJkVc8FWQXvUs+0KoZ1981JLDihGk+Un7P172p7X3KOVYyuAoSgQvNKef2zi5Z4wuEOTVrxUl
6i6r8dTpSeLSI58y7xunWU26cCx2jbxGLeXAGJGw1JyJYc1vLOoavhtiIHzA3GDaN+tqnbUbSFPM
9jW6UgOJ7qGOwbLw/p2PQ88wyRxgBmElKW7xWrnO05Mwl2MA/cRJ8tkjDtiK31xjyiZgzJvl8IIX
dE+5eKJzoZBPs95ISVXZxeaQB3no2v5RrYnH79273MD+u8kLh9QpADzT1IxKMWKLYD1nZqaRkPne
KBNRRJht2e7V6WWO4clPMIyL19hSzajUqqU5qPbIgFOV6pJ6FbTMPuPfKbikXxbHP3BfBImhcwS9
TNLPxkJhnGl4EDq43f7moMmCVVIEmfkutE+uJteLqiiQNqWIPRm8s2JM9AQC0/AKuQ8BzhrEnuU1
9SBFx7XIB6giLl9BSqkbrtO5pKno9RubzCcPk1TNmGiqchPl3SMVdYa3atHP5EPDZ7xmHWA7aHfe
nLmX+zxumdHqZBNi4ZzG/0NnpiUfqy9fM328IVybVIZPUc6e/KUTnk6p9DwfgPcDYDSJMoWkeBn0
FrAFialZQ6ZAj9InTaVg71R7ozq7YGKUODi5wpAJ+JhAo2z23+VPpt2k+VruWOik6NZ4/EDQnHVX
f6CscYCrnVakmz6hNfPmh/1vRCFhsTQ5XV2+U6yO2bQHiai553RF6joOL4+WP1KFAFYdTaLa+AOl
IlW/i0lxr8uXFj2zAZDqLRCr92DpRXxnIUrZ5b2WeYEC4riJGu8l8fluCh0jDPe3TSfzCWdj3rUW
0oh4CW+csed/UhzWE/79G95DhKN4y23TcEkLXHiNpWPYpguA/HMxQU8JvPVf4CX1eQ3NhmnwmvgT
fxKm3b6KxAO6QxCmdqfWCqT+XaAblRXN5Z6LpmGF+ph5zeUil74xB3Il4bdCT6rb0qIfrbF6VbaH
eVF91gx5Gjohy/3WTyyAmeGRb7W0X27PvX9I32ZNaT1MgwO1zRSJgYcN7DZ01//uYJNV0mrqZaoj
XS3/lxX3XOmaupKZ0UKEy5iYfem0hXUhrMWt2avrGsRyZrhabOdBK+GOnPk9rW5NLvtMcAljHAJi
eyLF5MA3f2117iSUnjeAsf9J6husxyoh4Yizps/nuvODNXVRmewLffjKB8m14EEaFA478hetE6vV
KDzb74bZkkuB9NH9eeE+CrB9yHzctGXCpIBVke8SPf4W0UM3DOyFCdlFzTu+4BmJS2AwnBNJfoWB
LWZN07pGDM2kIXmJSBW4mtJh4jCHnSc8nDN05F0+dRQ+05bemRYTo2gdPtZlymDn3xDAJv+MSAwH
ck6Jr/B5BAaGJC2ciM/QzQbWdfXcVhEfC12BYkkARWQA9aiNxOmo4Lesj/5kONQuL/XgeRjRoQya
4Sa0qDnTMmsNFxL+BQ11EQtQkoCzDupaQAeUc39n3K5aOiJVCv+jfWosVaih4w5UkooQC6qVEqdD
nTz5k/Fr2Pj36OKzojBZpHPS0P2MymR34iTDtJY8qWdza0omKSLScb5Vnu2TAQQnAhX+VVNyg+UD
AkX3n4w3Py6DAlyzLiIXLPKFw8+eueC6w6mLIl8fW2/QQJFnHe4Yzw//dUPO4QSAY+iRD2J85cTv
i89jElUANaywlii68D9/h89dLMNf8hbaRpaHxULHN+ioTmFNKudxYNW+TBqEoJIS+g8vCb4KfO1H
fCuHLHqrveAWmHAV3l6G3uPtsiM2ws3XmyNhSeZ5A9fJTJfos7jk2V5aA0KPjQZvgvTuz5Dcahfh
aKmtqBY239SoOT+lnQVUI7xycFJaR72WoLXAa3x3oMPI2wkmgkWXNzc7FTnxVnVnOS6qtJoC9+t3
3TsI8BGCut0JgOJv0OrM7CWxwa6YYk2LlRT+w2PyPBldkPZSYQhM4RfPDqxRpX8u7OwIR9HUcKWD
nKAHmhKZ01uhyE+YdTf1A4yd0Y+6f2p3BpgNgsk40shsei5vy7KpnadKj6VsEc5o5mR5lToGnVVm
04nDdwuvbSkkZyyrXrK2S+RWTqOa3MMsskCoQYq6wEpVCc1Af7an224T5kgIPy57NRcGXTGjPgdz
YXXRpfNyGawFohXH2rkR1xS+OFNNcGiRApNSxz4xIzAzdJEqKLpKOGz4onKTAAji0rkjz42D0vhJ
BBac7QNuW538KHXuOnUK+19rkGjbBmXyfWQ+QjRXgTeLCXUueOUe6kX06w1kX6sU49zij5QDkbSq
ebaejh7trn4VSpvJnDFsF9phpXECwEMt9bee+v8ERwBb7gSsSmdnqCLlVkWhrvRp5l78nMYqh28K
lBVM3t5aB6fRUy2yO8NWFJ65oZz5gThzhtHbT346c6sOQedpvEx+S3S6MpgjvG/tNLwjvACiyWxE
g4YN1rkZude9CJ3gWVesKekcAO5ej+FydnegcjTCpZQRrvhjSyK1ev2VSuWNsZhgPlhqm9i3n8sc
24eCT86+7ontkP37myg9C0nJXM4FQBXu9nBcuwEXmg2M0sgieI6uwcIiKifTyGec4fJV3ulEAEth
Lkq3od6z9Sh8Tsfqlc8hVgWdEGClUS+w9zSrrxJZfyCXFNG/oDZIm0fl7h/Mj4YTqup05JgBkGZI
u3T5XODO9x8xQ3SEV6F1squfTC40D80XA4Kcz22jeFAN4yWce4Bbd1O7UFPRzKJXZ9EVsfl0HZRw
c11Pe4xlvn2AwU6Obv7gVbHTuSHvtB9A3Gz55MFlEQq3ZwJcaIYSO47D7LgRuBhBSmNX4vjyTD18
mpCMUN8/ftM4+QS3GcP44G+uDOtNxhrzB1nD7/ezltD7JapfjQ4yK4+vgbMw2C7ntFOl10VaUuvM
Q+ovc6fGUE6SIHqammAB9c/gYkp08v3TGh8aUJEHFCrNiMP+BruTz/u/SjVuh84tgn3yWyfr2ZtA
YH8aJkP+0eflQzY0R4aagrdLu3ju02soF1fBfWuHp1j+BSuMFy3jacKhJ03UaNFUFplxppZSQmCq
TRvxdz/fHaSs8zcqsCG+KU07xvwWA5oUwQoWXdhBRgPVgwN1/Gelg6qt6UjvHxPA2HynFzvjv8oa
hndca2kU5qEMvyb0RJXeoM4wAFk9f+BzMmZSFN0kYc0TbGyd3AD1SfdpZQvnQuEbhiitn6u3BGaM
IsIgnU1qOaqFWAtywHPO6b1scH1jJRtY+yicL83GuY+ol4RwdkiTs9nRaIDb9jZafTsNV1KKzuOM
ovfVFKDRQMCnK15S0aIJIhHhSzmRvdPjrQF6E+atIHwkEKO/e+5R+Lf9WKyzvihqAJRwzy3NQdey
RhNd4CPo3jVwG7fhXMW3ZE9TQ+AHYOs9XdVwbXVMbwEqrHkK6DaxG4Ho8z7Xg5RCTFfSRlQwoW/l
2P4OwzHMLklTm2xlNRUKBDc6GicKTqIMtTBPks3JeSJUWtpniSN8545SSkUIIjrB+PXbkwhMoPuG
nXZiywS7hPtF99Hx4kCRhpq81wrG3rfEDrTJTnFBL50F5knn1C26yvpcJnlZAVXinHqTeg4bcuWU
bTmwNIbMK0Bn1HRUyUqcgM1LeD9pqKMs5oeh+P634NVe6aPKtdTLft4BYlfhgFNXCzKhjyqyBjl7
S4RewzzbUboDbK1Gi+AHPuQSd+N9MbGN//ib6RJ41N13TLfvHNTi4LUW9BuLDMxOubc6YEVpKt24
vXSvh/wMtUHgKO91WOU21oW3wwVGNID9/eM0CbIwAasDUO/YNlIL1pWqwYUqJa461ddXtSxr56gr
+MhvSNsjRkrSnoTfiRL9qm0R5cRzp2uJb7j0xIla/MARwmTgR5wl2bQnAQvhtBZkOv+5rZwsXtbD
MxVyZSLGEQMPGV0v2Ean9tmYjB5xHnRDF018qraPy+OzNlWELWLyxaLo+Gv4cAfLesHZG3JPKmkC
y+A7YnwxYxj/asIju8fqvuyND2nRHONxDoTpNfc+1o3F3wLuGCTu0eICB0qeiW1+ioTZbcED7lu2
LstQqpOlvXdH42qyJh4JyINkfYlw3Gch7zXgSJjOfGyg1Um0MKLTCbP8dt2MfmA8zkV7KC11f6w0
ZIE56hKMO4yEyeG5Y8tUX6uLcYvG7X42pF15FLh0bXu5xc7FUyC/ySUfZoPX5JwvJSiTR3wVWdou
WfOlUqLI2P321jcenQ8gAiAsYYTa03aZaOt4pHCEjv2N/UbVGLu+teQt/WiVVPn4LexpY9G14xFo
fATSkmw20f6YfGtRytaUm6DS33KvAFj/J8wqiUy+/xXfPPwI4+sKnd9R7pY/63H09kF/jY6GvYD9
Ms//Jk4oPiZ8jvBtdxq+UE8//ygHNiJsvcFy7QJm2hX3fo+n5eht5iMTvlCLKMwcxtUezzQRTum9
wdEL25u6bMBDb/7AQuAusIi8IKVb/x4Hqy53bDQLVCJ6mfpy6vNLT8ZG4bxN0vczaW435Qx721Py
3Q7eUFILoU4EPRcRevDjSFbbYjOKD8O14zZB1N02F4Pil+7ZZ4lEJlRtoBAIB+OaBrKgZwYMBrUr
yzprdd1/4/EQC5Y6ZpjwVv2ztFgkqvoAXoRvZr2qgPQgh/U4PBwwQU+VcVG5JlSj5v3utQ1dwAgG
xyoXe05Z0WSJ3ZlzT2Fb6AwDGF/Qkms+78TivORbD87sMMrWM4ZXE3iVfEjQJ6BqST57Z3UyJoK+
VqnNDcnNvqT5phBL2rtWT51lmqw5sSGK9ZkmHsGjWAT6wrJRRrvU4Rscu4NR9XbtYS6+e5/H8zRo
mumTviXa/YGf3AE8yttVI+CcKRDfy2aJUX/MDQm0oxpRx6QkXCFzN76QVZpeJi9PiBDKLuenB8La
RraSj37A2I+TW/Uld/J/LqNDIfalzOzl/QWqF8SeDkm6zldl4KUASZff76N3Y1nwbuzROBJc7B7U
wo8m56LGWRXjtqg/uYM6iEu8wLmoVUqQYltKCEvzxU2ZVwQft/O75TI2NalJwtvo0v4OP0UDtybZ
RJCvGFH51LbTgBzzZlRfRuLLfsmd2iDVEq9/GRDN47BxUdMMMfj4J2FoM3DbgqtWNQly6IBNUwN3
UOoWlB/iSySMhHLGVBpxvWo6TVnLAbzZILBQuWvTFnoQkxsQ24O1gh1X4Z23vMPtmfPiVuWneREe
jbgqQ2kCSIvYvsi0MY9hcFqRpyd23dB1cQ7ncJ48Gx0PpMxjfmre8SDL60QDp57BBc9LOc4dySBm
0YDGThkRZRNWAakkfyrcWDrz2kpJCfC4Y3JaLIqLzLCpisXvoCqRA38EmzP/ztdAJqGV7YhRu/MF
cvSw4alERCAdMcQmTtWpOP/cUFCA1YwYFkQwhKmU9fbdqeH7sEqeXIyLOWx/SVjrAMMHyoHStnnc
CmBEqVNWUJeFR4euGHrqq4wHO5y2A4aTT5ptRItpAkwcUC90FwkJlnKDtxjNr59RJs3+Rr1z+uwy
t/knaI1Ko/7zc+zJpsHFJwzMJh3UFqNn6FiJ8Ie3NUAPN3sedgcxXbez7I+VcMKYUCXMNL9W3/u5
SmlwY0EsDriT8s7cZ2nieVY6giBjiy9I0P2aWpiuMJ2oQGiRr84Bpi4nd2SVtXLpk/5vEfSpo9PN
M0Xm0WodGUuEheQmBn7RLmb2iKlvGtHIS1yonFntF7ufFN7135jOta1Pov3EDiCosLsJ+wP6aeW9
895UH3W2C5HbXbaWGQr8BMu1LFwtlPj/BQwN+CZ9YuMwrrUL/4ixqtxL3qiLQjvuUk3VUVDvRzCQ
zMQU7YacCVRhLzpXgcOqUy10wBxXgs23raSEPiwHN75gLhLmJojhyUdzghYl7I1BbgKa3F5MG3Mb
0impFbVoPZppOU8rqFW8fKGMbGIHBgX74dViqlwtrSLjoNL4WX/dTQ58sXBeFHiekN94N7oKzr2v
h1MZ+fs2J74aQcEdAAyStTMCqaDmyQ23/re8UGIt5B4odeXvo1p7RJzR7/4nDBDuUQOjX3IR6Zto
N5o+RHS9RCtX0Cz5bTVgFjxQrffOJjSB4Vn6fHBKv2Vs1Qa1du4qGai2k44SGLbmt4KV9zsbwOst
YtBZlkAEuH8rXgWYv2xcrXBVL07/+g7QwDk0hYzBSjJIR57rDlGOkTW7OrLzh2PZD9LvXYGR+/xo
iBSiCJvcIIltjSX+Aq4yvBhRq6BD5lyAxQdm/vlxr5Ot5vMdh8mck8ESr7xYEElRJs+oM1Yk8Wbb
u8+CkuOLFARxiqQb7mserXFVeGSGmSC2EAQO+0Bhq+q9/72FAxgiiaplGkYR3+cSm5Me6qFjvCnQ
3OWWcvM9uZoJ+QXdNlUTIstsU9SOlt0uXxDAJyAxms1bnt5A4DD3t812Xbi7mfeSM6Wf2ZmQPsHS
WOddh9Y9YE7oMJIE0oyH5iIJJXVydAuu6G58AGJOEUpcpmbRJd0RZ9NWYGrgzdQKQRygxNvmWD2S
gLK1F2m9QkqlDWWzrUKegqIIKgyW01tMFoKRhZJ15o9nHh+JLooIuao94yut/AxCFNSlM+dqozYX
CUPjDq5wrwVJ5g1MK43Dm0XF5GuO2tYZPP/i78/FSwyOy9D1NxA+atjCW/AvS/isbdB2TMv8swFn
NK4WqToh9Ssbvb4unzwzN0plpO2d/PkmNqYf8OG60+xv45JcmrEnzOVWVUi9h9Eo0jsTdy8vVN18
cWv6YzUFNsULcaeKkYZUBkNN109meqEo/zflKxUMz6qCmClENqFhNNYgxBI/0wEm1nVtPRxmDdii
/GE+A0xHjFSVXCHNnvZffLY/L2PVk7zO8hNFFSI8uu84cF9UBaFZl9fT7adtuIE9hv0SmF0QPJ11
aTFTW2tacvnnfA1FNISPww1qPua7igx4QKu24geXLVIkYVAlH31a9LMBcL4//03oRnaCnlQKiIE1
nPKev5yzeZygkNYwdheM98DFG4ya+Y82WNZt6juopplMIe2GGJz42zMObhycxjRQqjN3Kd3fLh75
/Mea6KmrUKX7Lpgpg4e9oiUrgE9gJ9DiHCo5ov3QdcsBxt3cnyAd38xvZrHwbis0JqRs7pwKr/Fc
7nL8ZKYwwL5/e1SxzZ7kgrsmrZWy1OT/NgZn5+lwuKta/yPjhN16+zngTCjoNgEc6snkUdcUx9D6
8qmukeTDyv02+vQrudxPLpwWBpmEXuoX5EPsWJLYA/qUwqk3uO1D3lskP0Zu6wK4gPcMRWwEOFz/
izvHGrWx3UDGNHvT+Hqs5YH/WfHGcb7R3h8Nyc7NPi+j7wh6Fqpxjusn9C2NbgJdlIY8GyEQddG1
hhrZbRAeZlhHbCRBihHfmhDE8UwZF8Dcc8obdYVe/rA4GzcO+Jrae8Tlnxhp03dgVOFEPekSBlf4
urgUwGxKP/5YrCs9b02adSbcUADivq82Xd1IHoU9LKtHLbYHfLjYJUvycScUt9vloa+cI0XQXFZt
kSgwbpnnDWWQHn2mfKzWMbOlwuKomUcMbLrArL60Kjvik27nZNw5AUUdwTuiVycbLLOnQdg1953m
EXAMTN3xUS3BUzhbYFBazHY0nxiaOGDuFluBEioyJy5xBO7GwzKhGvEyNs/OBrmgSVjKpJhKZSQt
5o86tQ6HZJwhQzGNWjzmCErnBwPTiiJvDFteQBxAMG7iN9GmvXm9fAFLjlUXmpOQ2OMo/OVLhYYR
uaR3gIWBc9p3bbUe3C5z9e2GaFI42x+HWjwRh0NMKKt243YR0k/yxbzQ6CV+dUz0+Nlz+zPv6b+z
v0A/5+QTjTVdVjU8uJH39qAoRzpNe7tunwx8y79FRl7uO+DEfjtEoMt7GTW6AHWh8CFGd11LtAz6
RFzlWXGXFVubThPq/Hg5qsP+haacClArm0puxPM3C8fKpUF6XraFweMelJzuMiEq67EbpckQQ4bZ
O2HQ9SuGs5mj9oI56TTnceWtGSYp5QVEUsdOBg2ZOYJHUsEBzvqUjDC+H84UMWumXAr2Abml5b0e
dnj9QkydTJIrjbryAV6v+quMSaSok0ToEKjDOm/T4+3hnKaS7tX/DCE0RLvBcWvSORFhUIJKdBrF
1KVpNoDq7bd8unechU/LBD2B8tNdQRjx60kw/D0n6XZOnSei1444zbLuw7C6qZ82LQh5gGLVdSNv
lluT7noWZxHt7BESjP1GhZzwlM55fQVTDf9RC+ebKlIBvb7N1pFFhhLZOwRb3WBVoTbabZsackad
Qg86WCgSfZUTrjed3IuS2JiMctmuIsvWkKqt4A+EXd1b19PRqloip5gJ7OE2yVDL8QcWYRXpFk5j
vbm3JcO+ykV4XlOnh+0a0SvzB6fdHw4qa/3amAdSl6kW2MTA8YoZHaE/GdE9rre1JT4bNO/bqFRn
Oatj2KcegFu0ADGCPpiNlHUF6ngxdEIvO5x504UbKV+tyeuWmJvajl9PqgmHYMyoFzPiQGe4aztA
+6rmwUGVWa7Eqvg2Q3Ff7v1sE6EEr2SvB7ehXNl3zJ38DCLjwDjunA4ZPKX7nBzi1J30ofUmuC2q
ErvdkZeI9b44In1z3DuzRLyM1CrLNMpbw51Bio9wloPHGqJWuVDJ6lSUjUJEaGfrdJDHPHRiUr9i
wB6YoXIv+nQqwdHLNVClvNGoEFnF/ZhNhiSQNo/p3Vnqf6eY/3aVgrYDD1ljATRpUCmKDj/a8xyM
my02zFeD5FZsOIauW+KS2A/HcXfsrSuVv/0zCajR6LY15QYE2pyh+gY2MBB5gL7SW83VNEsg5HqL
g7CFz+ePVp+We/F/3gYliJy/8XhHgh620N2skvwMVdQqrVSNeEvDOctJs5p3vWWx7XhllGomS47A
sa4nv5XFuQD1gPLo6isxO8s1r5ESHreLM+xrtyry/Je7Zx3mBzKYL3+Mp5Q4aXU6s4jaUrAx95P0
U+BkwNHRnkOSvWPtbKOzB5JRxgoDh93ujfSqF4/uZ05EGuu7DwG9Pil+J7pVa9t6sEPNawQQT31v
4sSSi4jYmp8S0yuImmIZEpnw8aVkXL/g+jgHiUl7dZjagvbKxl+W0N3P7XuukcBom1aOFMuN+2Nw
Ziissz/04miO3hZmrE1v+DH49TRnI/Tzb2ouxEiwpOr7cb/bfpeXlVL1QOBqiNOxSSjNyjKETTAT
xPBBTpgcVROkPYiw9MvNTo+CxTPevcZyT1279/ekS4FjFG+2eP+6c3nqTY/CeWjFMPbkgF44i5xJ
ALPHjBZLtwqULPmO98u8MF7g7swT+E8Fnyo90mC098Jrw+witO8mXMb8UNj1O+5qO9uoqwu2DiKI
jbjkqDZhGvoYgc131PvDVhxPjgqY1uaR4GxL4m/otv+bhYZznN+xrV2nD2BvJPxweYFNYKApfu0I
e/od/A80Uhnj/ou8c3Ka1Ttx9fOnkGnn8PmvJ5/BXukLD2+NbKYXJcRmNwONoJc9tvAyciEzOvdg
OtGFE3Pm2eDnhPvn7P14U8y6Spiks7iamMiG0v/luhLxWzeRi1tPaXxOegXso/2v2B0PlSxSvYbO
vOr1VWqcSqbbUcscwjyHkAGEh4jzjrUKhJSunXpNjNKQlqg1ODN+75GBlNbCme6NrtvXdbi7SUmZ
J1ISBU9HZkrFd7Kc3UPWfXo0zbEbItneKhCmUl5/iKk5ZDDELdMDiuhfB/qlBzAqefYRKYTKAdt/
Yd9/+RfjZGuhmU3VLvNcopHNTz41dfHLdyU9kyuUlIElE/s/TD6looLxgj49iFUM/2/CXP4lDxjk
2sH5LqZG25jl0xd1BB+hfbAnGzE8OL1tCDhNI+iL/OaDR6dBG/2mDD7Ovl+e1eh3dYlv0sWizzuY
8fV3IEPhPPciT8rU9brocVeV+hUzSIYweOa2R0dJriXbbvdMgD5LHypi6j66UXkocJMqgwbdxWGi
Ho6f7YT5PeJ+ny1eFm+U//PyLLZm1pZZtfsuhRAuHH87ClbjvodnZy1QjD81Ux8ppkFkSSjvuggi
ua2iw5AuDhpPk4L/TGEANNC00tcLcaWnAKhXgPPKVCwgtWzj4BinrKewEZM/Tf3tYSnEaEd2RXXl
ZpPp2KkSKI73vYXjmtrYH/l5EGlcOfyr4Nr9WOXkFI+tEvWxC7J0d48eK50ak1Lhi+LB9N8edPlL
ChElGdeD+liJ0xPtS7IVw39cMjQ6oQ/sQvJD8UuiaXZHRQA8se+a6bNvpG3IgwQ0aE9ZzflXlh5y
3rxJgpvPwXdGhEcnsEMSE8LW8DpWT17FHFU+uvvSH7hm8AZd624Hap/0w19H5wKNr4RC/t1/S4rU
W/jk/l6fElQJe6KkopcmPp+oE+08KhpbNEnOYXrd8C/cwHqOjQRjjV3zetoNwUANIh6q9GURb8sp
ZIVAl/R07o8bQw3wzMh1B6OrjoS3LvW28No6XgmqZBfrTTo0n+xM2GlIQwwHAYZiSuG7/IBd1jTM
+D+ah8my8473204qC6xSlCUsOeExBv1XY6lXPDWW6EnUkn1g09JJAyUMQahFdkLyDha2vIAY3pX8
5KfCa3VdUJtAFAjJAZTmbeP367xgYuvoOLBvWQbTO+Ip9J1vx0kG5canR0Y2rueAjopcAGulD9Qq
Z88J5dLIuP3AW5zrnffZLi+5FRiaQnZsfYiPWI5rE63GdsxZ6DFTAihlI3IASumj/15S3pQl1LN3
bn17IeGt5Eqfyd7wQ6Ob5vWeC8xS18jejdTpsJuzIhXVIb/RcxmHDRh1Xgy/H/pnKVDcxLmQU+0c
umrXvpvRYBuqaNaMpW3AY2OtETzZE6w6PtqSt12ptd1d2/LgVtXRwhJ/QolPGHmLs+WdH9ezl7aW
S9i54zcv8WvgYUbGmd7aSPYMN/plmZAVVA/796LvCWkfspcQ/cXyYR2fTMnINCiRRsZ6NiJg+qcT
JBkpbj0Ktm8rmORAistJKECDq7kbYQNT0C/hilV9GTSG5hBdjKxdMwf6+mNWnxtn8w6sAQWodcTR
vTTDwtHODxW8oFEWaljwBVrLG7x+VZSd6uzFx7uvwjBrlMttULEQaqpUP6S2TiBUaJmqTNH81WRl
EFJrMX5rvF2daeu5jbnMbQnJmZPCRDzjfGgrxArCqWtMQHea1bKlgfmzSCJdk2lk/QlMDlli2MpM
dObz38ks65M0EPFz4rd5wbfhitfrdUMzO/n7wNtHFojTReVFbseVhtd1xmyzQw6oPk7XF3Nl1ZPX
EHdocYRKbNs77v15nOuQVA4IgVHwBlznFKgIX+BIysecPwx05gvxtX3HfZMHroWGu+ialtl6trxV
8C/3oTU/iE5t6GATdg7U3Bwqdx+UL6+sHlJJAgDUJOBJ3JP1moPBs9ZLWn/0cKZvS6skPOFEdYfP
Hsrr4FGhyy8dqYWuOWDU2qD5dtN1vLl2XJNX8nKeAyBq8MsX7lEc31H24ySJu4dZgI9UNLWFn5Q5
RF/TeJaTf6FWzueVlLYafl5/he0cf8GOcmbo+C3SDaf1CxgPfeNQUQh6S3NRy01HEnyfjIa10ic+
WJ7Egmi0H28NgJAr82taI4M4z9eRRsG3jAhCbz5fprj7G5Mq5vUxrHyvGAkvPcLDiJr32eb7IJJX
BjN9+0eN/LxqiiIWqPuj9wD4xWfT8wTXKoay+vFA/A01qpWQLlCXa7oNowLNtBlaO1b1uj5pOVjD
5qkU5RBHgNZDiZyd/Z/NQ8C8CikdzklS1AGPhuciqqqXWfXiyedkts6UXvrDXXZ6SQZJ0lp08Xa0
LMyUf5X8QFNTTe9yKuzjnlnsDiMnJIrpHjpyJtD7qPeUKRYGsVVEw8nTvL5vPgTznSVLm297sOiq
CrdLdfe5Bypagbn30iyV479RnaeC1tq+r/16I0/3q5UnhpDDmVQDmeYZ7I3iRh3O9JNzz9ICUyo+
8LeC5fd6ttzS4zA7gUaJOpwo/zGT8MxwQwEOVyEp4CByYWn5INsr9desWyBMzsPg7dzZgNK1PDv/
m3FC1YVD/bjWru3eMvB6y5YHt0Tk9czWFACeg9NYMMNiPql2kI8CRtQREoNz5svg02oYdJjn5rXx
ehs2VmWADJ1QpxRpLTYSVjjDz9lRsL+BAIccb+ywjFWB1A9e5fa9xbz3/+ROJmRTm4a7wb0zI248
96tUdhZVvhTEvncaf2wk0b3idLpGdp9LX0O/eFerwpOZT4dTbF1Dd4m7YsK9loxjsdLQw1sPRL8o
t7hnsema15keKHbEhrKQNiNtr8EaUbD1HCJG77/uOzg/RlgCI2l43nbHUpyTFpucWHuh9B0Ol5za
AXDjPKXg6d8I1KS4I/WkWaqQ3rx/WayI8nbec0xjvqRCt94aSzI+VtaZRSsCIVyo/sRMEXZTBwbs
jbYgUIm9fZffgBfq27KgPzVkxWZ5F827tIs/jaUdINVVo+Z1YUy6kpsZ87COgEOth9CNQ/7aKZT+
3YjRnbcWrjiNoP3QIpYb3lqq46kWfUCczUlVcilCDePfrgw4errdPXaLnyC7VyljeHV0Q1flz1e5
BiABwCSFex3xUW6JuYkTcoR8i62lblbLzE6Zm0/XBAh21hxINsZ46OsmUVhexUbXoj7kG3B3SbDF
I0TugL6hCQnCYSg/Uf93pB11ZbCvkuVXh/FYYlVajZRDsV/tO5ClTEkOLcIemyFzpuHFDBDHa/Yp
Mw1Omc/FEWi1wgHk8OS34LfiasB3ZYwY4I5cqhJsd9CWBRrXMGzUnBt7I1Kf9cEx/WBeqZuwNWso
wVl1NAmWCJl0oZRPonMeCoIeIs5G1xnzldkcma8ARHtOyfGcBkCBf70tEC7CmU08e1U662eDiSMy
WFV0nAnl6e/ri9y+n/R4tQ2hc2Lthp8r3NoDiJrjR4x+biqMpYM3HzqPf/BKd3ka5aRFQwx8xo4E
qVFbPBFyDcboGgVuUSbdSw+hM+zIfpwyMPFK1n9H22HwBIPIuOjEq603o0aqY2ocOSf9/4feADhA
tLkl7kavMmc5GktVT7uodTFTrmF8SSquXoGFN5QYmaXgMBiO8gBVvjLSxg6DszPEsLTWCZGSvdaZ
O/jH3ca1MhnQOZtQK9+oira8mpJaJquKK2b6qV9aEqRXVHXahNsTUhQR3tBWSVnV9genaRoksnr9
LF58XZ7otb05fC8FlyZH8wj6qlouDYfF69dHk+0l0z8dDsniu4P/WAKeMnsP/l7jGK6QSyJQmtHr
Gys6jLWH18UT/a9ZffnfWwcD5c7yi122bD8G1AZ+ny+SV4j2oNuMEj558VsnX70g+mnLu2abX/1P
tZ67R5lIo9mqZ/VtYLqNWSNlH9xugyq9xYo3FUnZMR+jpVB6CaV5RPAg/8tc88uBrKTpUTKlLj9o
7fuukd9x+com1ucaLGXjul6zs1J25MCTvpoU9Kwibrw7kpQ1jKkPSM25+Y9lYtWrYR0qjIeo6W6A
aAemfNu/6/oCQik6L9q6+eZf9xVWy54HA11ng6lUdzEq/lkVj0ArsJRlAcq1EodusB0ivCRvwKIf
Hl4N4X+H87CBbVmoxQDIA/xzTBeDY81E/tsHcMyIeaiiHjEYmDzCqohF+Nw85CRUgwTQKFI7g8Zn
oiNiTpHtNE04SkElhN0QpUGH/S9k3pMCTlC8prge0Ju0AUfN+4TQVDvcKeF4+NLEzA09uZnwl2Z6
FMrOBPFHI1UPG8mwEwNwBMW1f1Fsh+PNmJS+zAHRWTo7LuRAomri7z/mAvsWUFu5SUkwZFjCOO8x
aB1iWT080vYQYDHJmbgJgc+kEKC7c0J1tFId2zGKssvu4aisQdKw3LcHl8XyajX4GnRuYJ+shYgs
qEeek5WqsnkIFlp7sIcCRwhwoYpCT7aTM6XcKtQyNdeyv/FIW9Vo4T31Dh5g5dKHydK8awp91/ux
9DZrQTpTGQhxqFObhHIYq36G8O4m1dmYgZQvDtDt61yXUY6oxXZ8Qw7tvd/RpoYnbhSOusgYidpl
elHW5yOEbUG1mhl3yKeWEByH5JaraMg4NjRsoIWQNi3kRtIviDKKbXORBtz32w9nWu/lb99ulBG3
oDTvFPHKqUJy5n/xUKuxUnR2HKY8pl49xR69et7CMqMy8djLoYIBlwOGlFTdE1ZfBPWpBRQ+9Rw4
+yFbDEXiu1noVNc2oD8nlUds8pbVc/AjuWGn0+Ja5M3+UwZvePXHFK/4J/UgySHkOcjDLiyObuqy
6QZsrv2oXmPvLINwn0ItyVVpwV70OxWKcAPwBc84e2bRnp6D+Q/p9yVLiyIa9hXjc+V1CyWD01te
k7GzdB17bNTvSdCMQZVaV5bB30/SroVcknhbHDHwNa3UeKRsUV8N42ooZSPnIMJlcMgT8O/W3PU3
K8I5R38YWIsalYgjo8npzDRoHfB4OERP3fp98QMghL4hlHC6NrsRIOUsrH8hkQYOq6VxLX40tGuL
Lgd1tVLP764Wn5RqOTxiXh0Eq8vnS/u0DD3umM9xkGQgwzO7T6ihVHYsx1u274xW0UwEbvP8X0fu
lyeMmeRzks/VZ8bN/L9JUmMMgE3g+Nk7hAuYozVb7LmodG81PxJeG7DzSaWy7f/Ow1ikQno9E9pu
M5QpHzmh9qhpLuuYoxjgaSZhcqa2kJvyRFpeMLFndbs7CqvLozWSUPIXdUkTCNfMaRw8kRzknnq/
WYWu2LlVlN/BT7oFB1Y6MvN71hb/3QhgQWuTnp8gac8dQzD1hFjmhkWJrR8vbJpwT8DnEGJ8RE3u
DAU8ZNxbU2+kyU9kGGSGr9gWfDbs5cUlvHbxilmyXiZJfXeQf/WyBSKJXz0F6DUXST7onvOXnfje
4lfO+FivDmR92ci2lXcZP3fQGJ/UFTdvX0lFPPnVz+evd9MsaH+zCBufZZoQ7s5oFI1qDJHV6UFO
y2My2+c6EJBStrJ3LqYhriAuVq6KdX1vqdFsKFM5sAvjARYT939LCwMolUjaU8MkFxIFzp1RvpBn
phQhtMWT8F6wlxiUqAZWeDk3ZW+9/sTTHRTGHbmm68Ze6JqTVAXGo6EIjzGMzAXKV+RdVaj26Z09
uuFyG+z23nNbzZDQVB8/TU7GAm9LmbzZPPJjxVcUWuIiJFkjEsavUIMF9/gwsSXzDUClhP82h7Oi
ckUfFb+FAHzJzAVAzhdHyft+Q6HqO9HP6+B3vpuZ0kaZ/TgqbeVidiHS/jHhUtu1pqwPRTuutm7Q
sASjdqoDVsLDiQYL/HBxjNKgvovpDIoZ2V3RsfIcPh9FaMqzCHF8w7tfQYk0Kn6W1dpH4xdDyy6k
qsp6V8y5t4ZVjxTwr8pfFxoWNFPx7eBo/wl7wcqIiljFwYRcEPLc6i+J87k2aZdwPJijUKNUnJOW
eszMprMeNbwJ/QhZuBxsuvTJpxjJl2QpqbATqNkr42LdqaRUD4TY9oamkR0sZuAazizkCRTS/l+G
CFjEPtMlJ/k7K0l3zeNKyUTFnpqDRx2Sbin2MfQ0oLDDYT8hHuTvJer5giY3cdra02K7mGjj0upm
1vdB8fJ1HOpRZNdWA5NFnIGGoQ8QQpLb9bUsqG7S6NKoam0oFJ4XRe9S+r1eC/TC9CFtHQRyYZp4
no/NEk/mliZJnSMOV7Ku0RX3bA++I8iIdS7tlmrN49DhU3xkqkjaBF1897NJlPMRVrSiHeTJTl2c
CSySIpJZskk5sv9v3rtuj4cNasaDY3GqppDYmxJEAfW4Tnlhus6cziCx7IF/b3inbZcMikNmmH9h
zmSVdQJrbf6D1NoYBTlI5ccJNIF3i0vvt9OZDUOMu5UI2x8I66GIE2SvcO9/hE4qTVNG66pKPjZM
jrQeOVELxXdflOTv2SjpUNWFs1UvIfTxBmvV4/+Vb9vaISMp0hIV+yVgvTkitVowxoauRCQ+Z08t
coleBCxXiVm3sIo6612adCmHuxDyThIMF1UUWG0jVdMCV+zIDwSOmq61vx3/Gv+mbbc+DJ4laQmY
i2vs9CHJbRzLjBVNUaOcwxQg72Oou/rm7rK3mpdBKMm9EPfZO8J5bYcXv/8BOon/qwrMA9elPmLT
565IlM+Fixvo+CcOl6L8TfsfLIiUoMEgaCXbzU5jSrnuLXOsI6lEKVpGJxXZfO44lX16zjbJpx4Z
9jbxlUD8eS8OjYYJtKy58xrPNBpnrZCESI/HWKQ0ykvc2VP85PeckADWRnJEdfmnqcbN0HN1tmQi
ca1FX2f/tkuLc0hfo1Ayt0EZJS2Rvw2hMB2RKdIEyda6/ez5kZ7bsUL9l94eIWoqhtQvKeQgFMWJ
DlTp+WbZwEZxOtMuamMFzmDjOw2bP5yTueCJnwJ50dGfqlfQscKMmLgXgRBn31yDas/zv8PoqTmX
nUdsv4r2ausvoYFPq8Vn5oFlF4/6Z1zRvyHqspbFZWHUwwh/ChtIGaGC2kt5wkEWnULv8LynZ9fO
BK//Y9KteWYm2IjDVQOLgZc2lOxP6zEeFDqyJFc6x1rbUf6Pae5KMAnT45LVYmgrkx6qVdlacXdl
6WAXdkR12HM0A3wqPNACHsqlDu4Z+XY5cLE0ZwWVD805h4BROqJNbTot6oLMz/OoGODHkGP3KMBm
CBWzEL+jNOpcl215KXu7gWnb5pjiTAo+WLWh2PLjlywz7g6x5lIO3Thy+VJzmP7hQNqC/RgXvcFm
6NlP+6iE1S2GrTTPGdxpbEv/w3qel4MPUQuiT2caEkAx5Hb9vW90+IT46tLReqG3iOY/7KHN1ooq
zsnwrPypnVDx+NfrWn+oGKHMervg+qveE3CKbCg/zYYqCZqif698kztSZPhTBzGGbrJWaMDBs/N5
6jI9q1/oBgtRJtg8l2AOzvOjcNaTk8E0+QaRfhRRdzzdR2x8nwHJWTjKKEWquwVquWP9OlOYnWVt
4wsudArwjUbXNOaNf16qg8/lmCtQmrlki9Dj3w/HOCrRel3rpSTbEtejbfEWZQ1IQvO+FvnTflWX
qA/+ZEhok606mOM78kskdfXr8PXpf90mrmWNSaw5SE1J5pdB5hqh2NFiqEaOHIw4hNkKq23oIgSE
nVa/HhaykQnU0wGjev+8bvh/NoQazZ2bUj4yFtaDONbySZbyH8Pa0SAMTebRPdhCJs8SekMIwW0W
jtIa5MX9Ro2plC93a0Ij8/430uLuenEg2tCXPyy+ZBMit/Fi3fS21Ldj7A9iAVb5/7YAT8+kThG4
qqHzoDJAqFVqApwgS+dzcAhS86EzOBTfCS2358rnTT2sgHsBUbgLbwM3VTs8h0lzgki+Pdg6aXw3
K9O9wVNYtHw40ruYMOR9+uRK9u7qLpk8MRGaGwQ6rtwUo7b2KGhmFN1t0VP9CX5dGsdJykwmJGTX
pLc4lkjTi9caVP4eAbCHIuQT9Xkx4wTQ/iN+m71oWzqRdWgE709SOI9f0dHUkX2kebM7vKGkT9kr
w40Ci6hPUc+oam2GERNVlK7099CfMiz9ipXH62XUFiC1uMspsmB91xhK3tKv6fT3OG88xhsz8onR
a0w7kQ/WI3OLiEezqNYFFDO0MiRZLL/loiIGTvzIYpQ/6wqScimJKimTf9cWwX1LeJnViVXBeYpY
ttXMfLa+5RRUFdmKndQJn7Gf3ncwHqeI9DVynEzwBl5kAsgzropXL/wxcWna+grYs7FOGxTrEIFI
kxwtdN7AGHn3LPU0rCjRIRnws+6HuYwzB7HtdcMExmyaOVw6A30GK3ga89VSs6jesq9VoWVuRJYE
vlyVA8w4/VQCIA8u9lXNJMeue3Hg3PlHOaaRyaQddqP7GdLPBvbNcx5FfEE+o78/ZNYmRDdf17i9
pQ3wsmV8bd8pkVi4J19SHGwxZ5R2zbzkZ0u4qhZvmEw8P9qP9I9Eondoe+DAn7oeSFJ5YdRqjEHP
MOQuAhwIc/XGSHIEFhC37d2OktfHhmroA25cY+HhAtjRtLoHv68aeUfLOnCghCAMjMHiTCx+KK07
V7oyHD/IpvihRZBhFFdEW/qJrZPYv5UV8bnJkCW716aVyip2K70xlDTyavqFVxoUgMA8bhGRtS3K
pt0uRupSY141O/lqsDi9cHEyRGH1TU59RWS/sfJI11/d75QLlNG+WzN2hXuxSPrhWAfm16vD0dbH
Xe5IeIpNn4iSLtZYwGC41e6dzR/MvYyaUNTTE0b25zc+tqj8rHH8/wyB/0MVG/BeKP9N2TCsOCZ4
OlxqKJVeAe37uYd8cmXKPYporHILelgZU3tvN71ccNVgLSvsXwNOYbaN/FfAYlAnYa0BjMDQh6ek
Kez21lXODgX/NDaiO72KGHN8cmI2Iw1A9mCfOskLkzhECXk4pDzio6erpJ0ZtTHQxj05JsujFI7j
azQ6enqBk3ttVnmdE0Tf89xYqMF5JNLy43XmehXEo2+hI7PcMA0gglhns3iQTppcPN8NZLSwu9xv
toqobZVDmuOf/VA9CFCKxwLjuCXauGqOSqMQaz5cutyX+AOH2/BSmK9cRVybieZnnIeFgnOJ/NJ1
0Dfj3m/vnNphyCHImb0ePftIyWvrHFoOC56oRT6jscM5X/sM3PO4jANhzsGA+u/OFlAXzW/Is0eq
QPgR613Mir92TLczXzqFZMnidVld3Er+L4rrKi6R3xMscSbpMQ+UAbGMu68Cta8EZfyWoLHpe6v0
F4WdhZbcsXVNSqU4mZj3LirY0bEpV0QDtLLAtijoAhmF4NoD5YJEAX8hJ31DahrxIVlPNYdyp/aV
vMnKFWvFNF4C5RC94HYlA86r/0/utwMyAy7hRZjMKA6kDzQPjk/88PAyNd0uznD0wfa6pOAOCHdU
JF2lGadNTokpBD4SNoQt4H+lk7NK3RnxurjMhP+7zZtSM1qKmwwf3AyuhjDM8W6gM2BL4O9/3r2d
zF1AEHkOcxkg+Gmc8k9N6T5in/vDXK9lSob7vTlkgMjxX3XmxbRWse+U9IpSi27yLNWTvfOQTmFm
SlSYHLOlCLr+PliXbft29hCJxSG0qKJmh44sX9bDfZOrPiKDCBVGNuCgOtTq/JB+l770iOW0k23c
Bac3UIhJ3cKhfNpweH0KZez+QT0pqoA+zdX6OwgvEHEFjAqlc7OUb2DkLW4a4BYgTVL5JLnLC3N+
b3fqzCFPeSGus5179NCQB3nmOjlNNqbC5p/g2CyUZ7D8sUMi0+KQQmQ/2HM1AqA6ZgJBV796HZdL
xFvZ1RAuYV8yFNIQkLa8puVRd/Vkq026uayypBa8TffGs2vCeo/zQhZNtxvEfMZyS3v+GO4XFQDh
FWyTz7/To9pXddx8A4PKdOn5Dz4mGXmVN9+tjvJQ378VDFkkyLEd4tnBUXeD2tck6MDx7q5iFBIG
KmoNSHrcGJvK15vH0cQsPrqu9O1TkxtW0RVjJKOInYG10ZbJYEBfE4o1G43j+dDdrgNbwJxgyESn
RfyPWnT/LP+H1pTwC75/mdZ8ARY5q9KyLuf5r8y2YTlhwO7TX8qoXKLcI+ASTl3f8poYM7lr4Szh
cWvau8A2B9XZTg/+kmsLqGQEtHXzLAqFVrIMIKBUwiNbxc43+YxneyPo+jOVOeO0lA9pkSOexgsU
evEYU/Yx4BnrZfy37iCMj9yuZ4HXVR2QRlxV4bhLqeMw7xc5dGgzNEXgHw1kXYo8WxEQLZ4pJlmE
xJizmOR1vq9KQNy494wd3NenzfbBKAxgWBjuMtl9NqVSYgjq88muZLsalXw3wkiMmTMOcDItX4Gh
wYwhk8Zv7sNo4XWwGSdy17mFWjdky+aLoGsoXoNXbB7ZFk8QrvzRdDPvPaanLQClv49K1W3E/zc1
eStMfd6IQiD/vuI5ljtMXKImetAKI3oIex5FAskO8aC9rE3vS41wWddIOV4MPQyO+puvBJnlV7/O
X9kdGr692zP8LW7XICadvNoSvEEceEOxCKwhK5OZhvi8VBpg/Ali1LKM7G5xlvpFXqoZcPYcVPL8
mUqcnSaN4ZkJD0U710WajWibVDoRGUvCD1aKBgE8ajn8TW7DyxVZ7JhgX01wxUZknk7xuO1kV8AN
TCJXNKmy5auiJnG4Q4UuGU4EsH95TAQj2fKXxjPsrenI8K6XqXv0ZJIlU72mhUtoIyk9Uw5ecBai
rQHY/wIn5NUb5Xu6dHtqbSEv/0mzyGiNh4leSmJAdQshu1oRcx6CG1+90qy5jlJhge+f3qoRct7R
llQXQ4PSP06KRnFwhQGH+0+QTKPHVseIusN21mCkIjt8RkoGZk4MzQy4XeDhfTNzlgxdzxAcivuD
hPLttA1yIjhqrHQKrcDFFbVbXY4ycrOQdcL6vWujzJ0m2JmtAna2PTMxwBf/xEj8oH2T/brAcl9i
c6qEvMyQNga+1R7Q2MlIPshGjbcitwZxvcIyD2le8t/1mB9uE/F5Wqs+hPctN4N1LBM4nbsyGJOX
IsmAEVVTbvZhebKd0hT3HVNsY7eWX9veyU/Xkju43bR4MFsFQmjCfMBrFFwDRkqTwV7SSPUN11Cq
XG1Ggl7u7pkNGUfez+iU5nPRcADXx1qpkQmh+k+cWffFKD5J/weJ8a1NzzxTDNv+aP7tu0fOhwSV
upKa1C8km4ZtOtqDWr0hR7/1GIQygVy1v+KmO8a7s13MUP4NhHnSk33IcKrtrYNxTFY7nM8/BEnK
9VpIYf0XJTxTfqcX+6lbDZprWo7+5M+oDBUx34EqMVP0os3NLATqDi/k+ERQa266YlDI+P2OlGEN
uYYqvegWBNqh6s7P56I4JbUbG9gefGcjIkyrVf9zSjUV/78QujQGvv+g9uZx33v4AWYRamlA6h99
XuiEB9uDRn4Y2nBqfNgZ1mg7hUjy8fl099bJ1MYUbhaEidLiv3uvs5PeLL//lNbD5Bhbgds0+wnb
Z+bf4pHqrAxTAXbEMnZ4O9nKFbk3GlW6q4vf+dSP/zw4uJGc/OEf/yx3hGKvB1vWCzuCrYzze4po
yqSqiZlZPoisYNoILq4ne7urtpAlbrh7i3jjsRd4rNOREESBvT7VGvT/wpjRA4DNuoHOeyfqFYZN
XVaybWqX1hriaJ3/8Ww1GUFBbnoY6SXkENE21lk52x0KChXUElTMDYsoR7ecpgB6aPjJHzcJlPgA
1fqY2zZd/3L4IwXKmVFmceWjl1TA+vsU9weMavCZ+sKEeOmH220WzuoM1djTiSYiylceHrTVFo5x
6m4s5khVTwOEtGxuOrZWGvVuhRUZzxRAbch0W7x7S/ffS9jRyDYCOdGOuJ/Y4ErrORXwBYzsy6LH
i/pYS7TCu9peWWBpJXqXqtNiYEYDKpCCUDeh+Jo3gI2GOpRLIK1t3lVcL6v4NoY7f2WOdTenNWz8
Vu+tErh1Qu9QsQ/2pB2UUPsbcwdn7Q7Pop73j9D54DobdMMbcYLnX46dLYQ+SYiTiMXbzDBx+pUl
300N6fMt5pwrhrQKR1Pa6R99wXmZng+tclhqeNrhkNRHg0OA1T01fFPLewgBRvFPlLdy41EkdPFT
lQTPOVvVrMHRiyI7jXI9jO0edptZJhRshXgPzaWphWittI2qMSxmVc3Kg2mXJlgK/dkl9kkNlnDu
R/Yx0BuoZkgdRYs5vCu4xnFA+deNgSWVUPp56V6GSNx/Bi2L6WAXFVITc1XS5cbkti/8ticdcERs
YkjXIyfBatVteaKwggVBTfQjEW2KoLLekj55g0jDrJ0niNDexamcUU6YlT3kbsPvSEGo8p0KopkM
Js/fqOB2BTrjVLV1GYSMNTrlU2prxuB35GL9ewGR1pv7DzD6OlTWbxSZk3WDeAWq6/11edJSzJnO
3yPVb1uCCKszRNpPX6ti/AgZDiYPOlfhMkgsoGcGUVjeIc7tsQvRFa58CuZgbCu6zQLXWvN6l1+Z
h3raV8vQG8/EGMaJ/o96WmroYaIbyRTwz/QhUnVppkDsAxGYlGQLtMpGdksu2o+zWmmwmzrmX3Uo
Qmz4XHoz1iF2Vo2v+oufAti36P2QfzlrIaJSxR7+x4eB23Mg08XCESmyTgT4+MHeSrHWREjnwKuU
uz5s6Z7LmUdrqhKqzdJ5pu+6ExAAckCH7JJPi+OfzClbdeVZ1i5/GVtuLfl9Y18l+dtJAKRXyKoL
pns/TLU+rCxxhXX7LGKuZ73ar2OTf3lsPapjVFiK3SjFRzy+KmVplHn3j0/ylr9ChwHD5atmC8ev
ab8ZWKJXq8lcxaOiVrUiq4B+RF9A/uvZE+FvxjKVZ56wC5s9coV/UYtYVxmZOuo3a7WGylb9Kx+P
6SNUiIDjnGmKTrvrXp7aLS9EhMi8sOmq720KRW7M7hA058IqwKCRW0xKp5z2d/3Yd0CtoqvtMCnu
Htw3aD5dfVBABiw0iwIaOZWd59vW6KfaSOKG/2vf83Mn7X1lOIv5LtRhlzmdfyNA3ZSPgm+Tj2l3
VbgLN0wL2OUO8dkQUxepWG0UevxxLvtEyBtWgLyNHMGMQcEZUK4S5t1ohU74dPUJLNk4LYVzJZGY
zkNwzNfVA1zX74tlzvijwoBJ4t1vhGuCAt0Ot8f6ID48yTSzwYuioIiZ9NKlxUsEZDnGkKzyOlPR
KXhWyInD4NJg2FHoQsfHT0FNkXV5d9lHI5b6gVXi4IqDFwXvduGr+yfYDTZT0az6hcvn7vU9l9gm
Auz1EDkWqM+dv/SdFskhJ2EFM5nNRtQwJjZveYJ6cbeba+AiOUN5RX/A8czxjp6kjv7+lkhDoh5N
cTqW6M3+upycHYs9+5+XB/4FralTG/Rht3NBnpoPcypvX82S2Tz1DSeOCCGmjx0AB+VNEqBXRvr3
iRgDwOERxn0wIhFSHxmSZKkqwgfxjqUmSk9bNYlO9b0Ef8ObBMv1k6wNFi49orHqjUbz+X1HPigy
rUtWoyUB1olEJe6g2D5d4UJmKAaEA04IA1ynwSgdPigqhXeVVsSv1kBBdqz9E80RSKbMZRsNG2IJ
GFNRDyKTDbRJmbe9/Hov27+kDf6Ua//YchZon5KBn8RFXGkZ6AzlBC7//TtLsfzQedrrjckCX+Mr
WqTtVwM4eMKxqqiSp79LCKP7J9QxjiMBcPMg3Bh3PnLjhIx968J9PHqzyDRF4f6wSo7Cb904Rl1X
MKv150YMrZFMCpLmDixDkissD+pPuxoqd3s4HQkPaIFwPtik3uJvMZkQdfou3jRlw/sk9/0vpNPb
p/guvyoqtPIMRKcI49xLwiG4jlLxXx5r5DNZG9yQ79e0rLqCKh+kXGTqg7VVqtxqD7nWfnmVYsCt
5km6z0Wgo2o0k1cjX8pEbs3KnoiAKdfeK45DYwarU8ftVQDihTkZaOxMB4LbthRJ+dHxmn5Zaukd
udxPug+7zGP8ymm9aZ2jci2DeXedMJ0eaTDVUTzM/b1bmin3qUJX3PHzr118cySBf8BBL4EL8R1W
Y7y9gVWJWRI7Syq+U4GsHtE8I4u31ovLP6rAc2NE6PXGNE5rU5w+apeoUk6h1nrPy3anxMVtKSzX
i8QFtKpMv1Jy6JCK9Lo8zPSKm2rIjNg8qUBD9WlQejiyelcqYzzmYsgbp9jeh+eh63WGEu9mkKLa
L6Yto79qJ1wSpvDLOof0gsIWbV+nLgjqEF92Sb+C59UGBpYHLh+4FcbinVO/UXizEI90ec6a9/H3
zgPV4mLGlWJD1cO9UMiuuo1w9Gu/qvjCyuK8c5jIKo4yBIhsu6nPLpNWQJxDg8JOOzmMA1KgxQOY
FcJ7vSjOA4a1v0/TKpplgxMO6zhXjE+GR3RmFuIVFq4/rK3A3HhFH0lfo95pYnr/oli5Ayahr3PI
KT5EmvBxrDE0rLGJTJehMugNllXb+nCADDD3E5tTbXvoxSJY2jfnsiAqqd9AlJVz3xV/sQN6t/d3
OW+S5BmM+lnxeUTK6BhxEGwJAktkKmD8GSCaZE7To8wqrdErRgPYlYaVCSbmvQyTB+7b8Wr/772S
tv3yu6/pRr/1g6j6hiHRnqNcxklklIyTTQuINb7udQI8Gn2jd+TaHFM0euklj0Nt1Em8dL3pIOse
bofyZajVA381QWCQYTTC0OcXYwNeUz/IbN8cgErqbQ5oPD50XfUzhawC8araG/8383mTNSdGzl8h
R8vQnO/saowBiBn36H8iitXr3vSLdV5Ucxlp6NgMeLHSWoj7U5sEa9TUKewwLiKy0EyZ3yjLwZ2f
00UZ/oaS7uWCF5PuwjTaEaGDW+CJBWe/iakMmrFI8OAALB+NjP2SKN+ylK0CftnOoyg1VNr+5hcN
QRCxqIZfMahAuZwkrWxg6THVYOxjS9eol7EZPJ0bmiCyCsLBBEEK4mn1eyqcmdESe/7/yQzPBjSX
Ssz/Df9Z7S5dEs2YFbrA5HsrDI9crQ7413DIIwz77KQOqU2VEC4wwjfy1AXOLG6flGW0+zsbO7Fw
pDiYwxwuSGkj0zgoiqWN1Jan/C54/RLOUH5iwidwa38zbcAQ7DZ9AX458G4jPy3e5j+HlgPZxB1N
CdJXFkTNrqZJyF/QSA6j2ST9sBbNKV2qkeDAmTcULZvRQyOattW7nrvy8XFsqOSwlasT7fZWxRbj
BQkHpOhSBZCsA+25tbRLVyl7UnogtgpUqaRcoaXudl93TC5ouEs7KE+MG9CmvwGldX/pjRGvcLDa
VfZTUhbGDiUfR3PKbAqk8HLxQgMIFOfhBMqQnmKVeLJ9xzB8Q1vnu88BNRwWVCfVwJr28DQ+GKE0
vF/weZQyFjrM+OyHTU/k1jlPJJ9LPwQOLpP86slDFWAQy1cY4qpFgrFoINc//TzlTOwXibS3xtb+
HjpL5zPRG92WhlQPw5JMbSM7LsmW0IQ9cwp1kb0xC98c2hMbDjf5ajJyKL1M6X7y5uzQosSgeyNR
SqSf8z+Sd4lg/gWqZaE1R+f6nYTA8UXQbapjbFaLziDFRI9z6THv0zesBa/8fEpg2Oqv39NYf44p
LOYhkieaAME4USyqvdVxoVcB7i2oc61qePjJY0rou/klXqWm8Eb/uplQYJ9511jQ1rkUX4lzu+Ec
fDTAquvPkRObm9QwaC0WeIN/rXr+Qw9Pn8dKEdRrtfIn+ruA8kRRxtW4JyE3N3Vy8vv6zbnmfWf4
RsADGSfQt/+qh7U+9yf7tU/LQWSkxqHqLiKtq3DCKzq/p8vSrcOAZdcnUlGyK5QFoestVJPWvFT5
ivkQTNaAzOGxN8kGPY7Jy9k/NNRIbxE7EV6Ys3gg+9hj7VbR5JMsFOu9451r3NqyqLt3lzI7XcrM
C+5b0LD93vfv/EkIho6TkmvPIPGLnFtUZFvSWamAOSUuctubn4XHphjUBScmk2UK7bixM2AdTWC5
WQ8sOu1vyHgX/Z4GhyssIu4QhDqQX9MFUkAL/9jizTqqFYaBjmy6FqKCKP22eK8MwxYbDgCaFnEV
UVJCUveoJofbHwvslQQiZb+i/wBVqY8aLRo4tsVWH4T7PEN4zoxOBlgTXpx+rsMMaBW/xAvwNscj
SukdrPumRRtKjHE9l6w4m2NV1/iOBx6E81HsXhf0NEYPqM06ZKILn9FKp6kHukkYWbp/emChEgG6
sexfAw8jh7LDo0+A8qsWBbJwYZIN/TiYenoPYf7k9ce+vnxONJhRXQLvIhwj9useeVK2a/sTK2LY
qCrtxA9Px7y45Zp5oy3R3FClv8Hfqq+ux/wB9PiMSm3FwrRqbe+CdI6u1lV2KMBL4/d/YT+4dGJh
gR9Aex9cbMCF6Y9V4l4sNModx4mWlQx02hLl9JzsKu8ce8m9JT8k41kI0hzyBYalZpn2Z1bHg/pE
S0McEMCs3V7Yn4ayFQOJNC+6WYqRbO8IZgTBuJQ6drXYAEDmLuhZm/mrG8Jes1STHd0yT+Ujx6bl
9wrEI0qK2n/RNjgUfmzv9LKZ37ZXZjY6y9zCDjQOGDfg/xWC9Hmo7KGZLB+4YctiAlZ5scjiY8oE
SZHwR/CjhBruoc5+Aym0iWMns9zyy8CXNJWDDol5Nn8TOQ5tMrjVbYgYZLTIvmRcP8Po9XmDVl7F
ivznF7kkQJQ/pqd73WB+ihjPemPoSy94DsnQnxhKOf2ysC3e9Fd2lgXZgiBZBykSp+JIg5dPW7Rb
7YrMPiK5JQDe4i//t4HhE6E3tRTP25mKsmmgPmvzSJQ1oobnIgNofTJtLZQDeFuGm/l6kHQ8kj+9
feoY1ej1Zgi0VxR4uHcMgpTG/QYqBKdoK/NNQ9gxsAGqgugvKQDUlZ8wbjROgqDB+gbTCuWqCaOu
EB4D1VOkWmOH3yrPkFEskDGmskLzW4GPG3vQf++4JctvfMYb/VPEB4o+MPeyhy5PUTlq1Yv3Hpla
zcFlm4yW/5+DOAQdvW88KguhPxTYOwtJYGraHFVffh5vu0QE9Jz0nNPNmgJHyUBV9ssE0+znvoFw
gnEGOVy8jp9wFvDT2dPcbDlMeUFsUZm8U/G2SrqEWA5RAFCE9bPl7MxVwyRGn7zQhKXAudKJdPQl
EM7qk3CuZ+S7Ek6nKDAryufBNf/ytkww6F9NDarnkLlXqbRuQJeoFab3GWbKufmk7zqybmMch9Bl
1JIewTSKrCiDCFps4TzjhVpWT/URErvB4rhWZdCIMEJvUI6KEUaakM9SEs2oWJFEWl5B+OJzcZLk
RHM0TLzKk22JnCgA71GYwX8ov/goKj1lLc9f3VGXbk8sfkVlbXksglif7XjbdJ3nYbCzEZlUV1NZ
AJK+x16bkHh3IRIFIpdaoLMuMycHhGYU20XTO9pU5X0K/EDHnDSu9cX/hqgkbu6b6d8C2HlgbjBa
75/54WlEBSY5htmtd9Peg8DQIrnrH8xaNTRS5jv1L12n2e85tQPYP0l8OeN7pFAgP2kZ0czbzhcT
K8gmUYa4RDPyIijZevApSsEjuZ1FcZ/TlNfgdpKaKLk/L/kOu3Ign5z9bkRadDOAOmXL6Vnxp49m
GS1DCZ71WlU5VDGvy4tO4IYvla2CTwX2HoRgWZQSmHTk45kvxvGbxMKeU2tpR1Z6jes3sR/kG/d3
0fAduGZMMCQkn3WHe7oLx0jrTZ2EgQbf81wedo39X7KXCxLwFWcBXkFancx3KZWXUtfZMZuQJzO8
THwCJ7stgkeRU/1T0q6nv9HeuCTvz96ZvdU8RkCm9gjvnZFRSoCHMvGdtLSh3SHpC55sEUoDVtZY
oFjxWzpgoE7jZwhsZDnoh38EveWhgjeiSt8G+1YIGRdr6H8M1sCj0iHRnM+B4IsppoYyiMEnOUIP
HY/Q/IeZvfEhwwJ0fiXRLnS5nUIdjYHZdPMHkOmB6yVIfMegJBJkJsDcOCxZZHSL9NzpLqh9AhcU
dSvavOLXcrqwUMuCGbkqsyOZBum05Yhx4iat4I8f/vTuDt2ghSn6IrBr7/LfeSl6aXUgRVrV0TT7
9yHgSwkp+KMc0mZubz4YpX++R5S0QK5CLxaMHaZAASzpx7o5NHZqPNfXNHr9w/HKJ0rAcBOKNwUc
txi7/5abRUsFS/P0+dv1+UzVTaloKLvREzPP5+q2O/4Fo4ncG+tKzgYgsV8tvBOQlbjCDTccGcjJ
u4idiVT4gG7r5swD4GQwpJFRBnMBPqh29cRHghIqjMYbgEjPg4+83ygMDZI0VaQJxCpRqpsIZ7do
PjGSns9z3R9nugm2S5mKKi7gJGoro2GchCay1cepuWFK0uJ3UyZ9EAgEjXg1Xe0Gi9JENGWHrF4V
bfJHprmkJhXAVJxPdfCDsoi4OGCVRF3ry5/+3twVUg/eCG9n/PtBwFM/RDUhNJSin2RRqZC2GRu1
Q/TTBQtZprhhQxk+3TCb3hH8zGZ8SeydpqexhJkiL9hvz/F7yg33LEJUQj482rBiKubcxOng6iJk
Q5OWDM83W6bOJWZnuCxGdOtPX98I71LZbHT5dgHjM1jq6okFykVrpYf2yQujNCIvIZhsPa6FN/94
ka7m5S+7GKPlLzXCLCKxOt5CROVsE1qVlP3+3LxPLZ1K7HPPGb8MS6RdX01bxV4INR3A76iT8LA+
SuP1Ssxh73/BnUJUQkQM3yTOeFipw/6bIVPmjEV0XwzHQyYz/wMvsPazelO0e2m10p7YM/I+m3TC
zBb+eFHt1GP0vB9SgWVgm3OJp/jLOqtvAax2voa1teWhTpYAia1ZXDn77GIlgA0aHnMAiZU3uxiU
Vx+k5z0HogXaTAFhsG2dtEnuJrhfzw78UstZp1Y1GqXDXeZ2HOJoc52eSZ0oRgFqZHgWIOGTuoeb
xmq0aMCqNHyPFkuOxUgwSz57dXtAJBVzO/6DdURW9UwEwSl+Rsw0Dzr23TkI4BJwJgSpm2s6z37L
KKbuBtWntqbHk5yQOhUohUy1evWG8pKaXmLEz90ihIofDRjBuZQglbe9iasWoZxNgolUWxPIxk/a
ekdZPq/tVSsmkDCziPQqjpD4C7pxmyQADGLQiUsLuNQ82AJQ2Nu2GFWUezCelNl1Pd6sYQQT4pAj
Jd9zL1jYuPXKT/VRRIy+pdEa5E3rx6WxdbMXX4MR5S5NGwQoZ6M3eTCkv3JDmRRIqhP0KeTsYsLu
fP5zXxQUJAOjNh411wUgWGMXPKfn9k8Sp0s332TM1Zq6pvC/IHXmNNWjHF0X8o8kbMXmXph9v8z3
2G2MQ9OMGOV0ssE0u8eOpkxuCA2JnATj2g/C6KM1BQYpidYOGaXsBR+5wy0GJsaI37XIxHnccQ9S
Mp25NUAgEfCs7FbgQ6vhMFFVC1cwjSOffyyPHtfhXKyzFP/bbPnR/g10UA1DDHHXKCdi60IHq0bp
jHEF9tV8fVEaIxBu0o2oNTUptO/ATY0lGryKPKN8vBfRh7HsjBG2RwkiUfWy9Wdcq003zcfcvOab
2S2JUylGrLiwNXYDg1sL5vgg3YvJXt+8FUJ2rsEJMukWVLm8MdUJ8nnCx0uxUryJz/ISk8wRDnwx
gvj1wS8bTIh26vWNE+NWDheSJS0UbewAdoxL9yMdQLuiF4mLLxo5rI0dGdNfmMAJEK/G9YY/Eokp
Xtgs00VymbzBoUhg06/bYY1Jhsaw8DxHY+pDertRAOyKHEzt8hZ4kE7TC/nuWI++uQ1oouoOKQ6O
xlqYGidzxv0RdTcm9hkvh6oR3HntiEuNKd9HOblG7OMz2KDSXmm594SGH17xn0WFmLPBoENZe/iJ
joZDZySM37f+6nrlpMIRm0tTvG1ecofuZ1VXxSViIlUZi2nw7UK9qAytorE02tPWf+1Cm3IR8dWi
DKuge2lsa2GhsA5/KxThYo0AUFElWCmPjD8Z8tRQLvhQ8+8YzPiOkQ/T0JqqgFFVMYZtqHKmIp4m
oEfQjEC7CwXPjGd+JheHRew+SMjj8ey3zl0g/Qz7PAkvZPxxrXpFxQPaE8pAZF3+w61m6x/eeLUU
lgIAO5LhRnVJFq2LZAAi4nNJuW20QAgGbHygS9DtXVM4bI3DkADusGGVItXs4xNw79V5yEtORWuT
/ryoQ16RxrDgoSrAeE98zENKAWd6E4qL/jjrGktRUqGMwtZznodrDXz8HyO0n1EtxblRJxkaahSQ
fgUMsO6afhletBccCT0v8vct/9oMZHeIdgNxh8oUFtFswQ5jxrqod4N3ivwbZpbWXw3tQfm0NsA2
i10M3bpYoF+8CBbwmqA7/jzA9J7p45yPk3uiXi7z6qzx0RYbdWKcgU2Cpn7J1c2fa6xiq+edcy0+
sNMmnzetkr8A5WHbsRtIC4NG89vd+JnrlFYrn5Yy6K+lgyywyVqoROwF8uONI2PLvJDbUjpf1qX2
UJi3FegkLWViZu4AbMHnVkdxoRQ+8jFDXvNYh/tpeiRHa2mjpvytljAjfBR+LN31VvRr35k+Lc+s
Q4HNmKDZnej+dB0oVARbDk1bE1a6r/25fu2BdUE86rE/zSsv56hEQAteKL7Mekp0M1UwH7E7hQry
gLwpBipU83ZfDG+005k7I2quurNqkedR5yMG3vbagHTcMRfjDr27B27hxOedHasr9ydRyuoXQgE6
QqkhyPuvVny3F6MVcXaNy9QBzIrt3BGIpZ7FPlT0XrIfK3oUXQslRYFzq9XDCe6xTnUR3eclzVjq
Uoo+0a90KhFBkJSRlU+mcfA5R88nGHFYfhNDoAMqsKGfDuDSNEcZonAAVtqi1rtHo7WPtfepPoX+
hgelXhPVVdfZLHkOy81njlmyjpo6lkO9VOf2vDPgfDGnd6RPCSgWKxzK0B8wHvOkfzbD/I/euFRO
v2WPFY4acajDrQrWXUMzFtQZ86FUOrsqUB6mvb8VpW1yPVd8NNpOaQur0JazIGDEpeCQnvksi3Rl
zOGuwQaeWKpwzSLNNgEUJYt6C4kPNtfmrTjD3ua7iwNaygzIGaAWntwkeUijEn1MbjnukIk0SEla
jUKca3YIc77ugq/Bsvo74wDf+Js/gfQElMCfZQwcBDT7BxPIinulUPAAtSv4CymxCwOBLd9UAUvm
32CTgSuXsoMKY0GOGBHRfEMQEicjqH++3rhK/0cin8SP4r87zl4DFrAPDwAdAICkWGuN+me0WYH0
6exEFXkQ0XZSeMkJCTqehby/HJK3hn5V95LC6h9p93FDn7rcULwvk+gXyD+RFo/b918aA6aoTSQk
fBMXrRhE/uK6vKshkp/oTWEg8W8Da9BqOXS1uKHEyIosnP3ter9AtfY8JJRegkj4KtmnE0ErJU+k
48ri3xTdpfGxhCnGKWmY0gMTJqGFfEihd5P2ch77ymd4ZhAM6AHtDaKuteW2HwAVpjD+or0q9Ekr
SYibiazbMmnB1uP3dDfgs7c7Z5+8xtYvCnv6ryDAfgzzi2AwU4qAaI4uE/cz+gBqlseJHh8RYjum
zvrCNQrcWWnCmvVaFHhXlP7tDMIC/ZFEm4UhEkpRljuB/lf4Ne3vWV3Vv1sp5Op2eQIAqPpDqFHC
wJkV4huqcpxqOVOgdpChsu82Lj2Lapw/R/aJFKl45DFtc/aQVxQdngN1GR8uBbUYj6mCkehBUEiU
BF+oRMal1rHBg87QBvHv0K6PsUuaLoNz7eSUec+jmgSgfr0EUEKk/6MhsoW8Zd9+xRMARrCYxJrQ
NAnYHHUFaHaAxyk04Sa8fvExjzHB3Vq8V5kAaWVzyQnQ9Qrk4fWh0yHhxUTPwRseOHgr/ao1w9hb
unqOkV7WaAtIG5OUS30e9+H5q7vJ4Y0uBcmcBs0tHOn+YuEoeGGVaqC+i1fpRqbY/OD/mN9tLQ1/
HCmIQpJ/YPgwnCEwrcAqot+U1UKG8CaiWEckyE28EV0J+yorL6GRwi+DCOiBb6zwl5CB0b2cvHuD
gOIxXsWeApky9juZVLPWVAUEU6UDdfEy78jOlO0vZirRbMdeblU5Ne1203QVnTHNNzbccb107321
t34ui53Q4tynJ2AXlGRut53l74ccjsOAyj8XcLjOzYFBfP79wKzcYPP7NY1c+WPTZp23dFYW/qam
Ij93zxptjtWU6O2xwEOovY5DUuN/S5cxNe1GO8AC2I5U5X6KGZ6g0CGQH+C0TDsrsdK8dJW65fZq
LOr2Jp8antPpdEIkGOTllaDFYQUtz5VUkW0vWGb+lfo1/DN/Ra2K7n4ox7eZvniUKVhjdxN/1mWc
R/g28IoPxtUZzM6i6Zz7bteXKk5TjgBkmKbnbDDbwaI888wTyQEpqXkYoAEZGbmiY/1w1t19U4Kb
I1XO3Xzrvr3UaHIFXqQGB9gZD6EFysjDBGay9Q80VCFviKRmfbP83YJjyPK/1QBgM49B2Ope6g/z
rRD74IiooHeU2snmiLyAOHnTQ9geGYjmow+So8FopAEDFjipe/7E5puuHq6vleTYR/5umDW4TzLv
8GkqBBShVUyS8aEArotIvGNnXSk0onClUHuIkKj0WfRTLtfRo95BP8XCEY+Lb+5YfC1jbLnYVT+e
wBqCpBzlbhel2QM3btpUU+AyrbsDB7R9skLcMnHm0+3zFLsDO1U5UkfbgmR/6Sh3w9fvS6GgCJIL
23/nSqruSk+FzmBRZk5fFrYCS+v3UQKJ6aRtV7iOgonxvDbMlvIUdPh9Oc7YL85u32h8xh6372Cl
YIA8y/GcV7DuWJPi7+meO89hCMjW+7baN3zVALIcEUsmHUiPwcJ8ElrPwO0Ky8/SpDqSwEhjoKFn
WRA5Du6a5lyh1pr9b+M1yWJBMZuNw4deYebf+kVcYlCjF5oF5Mr5GhtLtTY1/BCkCTMoRI+muR3x
MpSrlBfpJ4lJ4SKURSWEoGUn+CE+Ci5UJ+sU9WJ8MEycB8p2nAtLPuYffBA5OXThc7GaanMUbHXX
JG64KQp/OXfoYqEXnUvPgTydopoz6+wxZFkBihbanPlWWnzLNcYJkbfDDPJ66G8t0Mv3zdNMI87O
GY08xs4U00/BecCMopW4desc7749FSWMO0jLGns30kuKCQYe5WeESdvC1pETzim24ZrJ9XnAZxlK
6Lo76CKR4rxDQzTKUhvKSQ8cgDUNNeEeFIy4SvNQfcOxuzVOIxxJ/uEQdZjqKUPFh8KpDHMNbR5I
n4XLuyKkvFN+fy7Uo+qAPRVF6vYfmTzPwmP02HzZuCYpuKEhBem1iUM9Km5mYK1TF36aOsN3rN02
QK/3cCCX0ss4bkiDgLTbxgvRepu6jzVtLTHYDytpcEpgB3Wxp2x+tGxvu/hZoe7NJF8l36NVwFVw
fe6/QtyYckuPXNFdhzavYeO8+0mDunC23eh2mXCy2h4TQEx3+K6jnaC31Kb1ESAqKpL5gYIQir6c
6A79TwZHehAFKlPvT2mjShpPLwDaGX+qK/k6h4HyEPS8ky4xTnPbhIq3Nym+g+pipY7UCE7kFiFQ
mXLfBdKddaLEZbY36Lw3p4mXCUwCtSe9Q0UfVZus9GHB0z026S18GEGbHKomZo9SkiklIuzqYJu4
29RUg3JdSm4uzhDr8rjA1Coxda+jEdEgupBCmPx/2hqHQceud7O4cYwh8gBWrzDwpR8QZeCEqsAh
zxHPLyuQGEebWtnrRthQGky4/xZ9915IkxBforDC8n0hemo5f2waVmFMmpq/8uAWRPceZIpVdf0D
jKqI7lnKsfPT/sPZPQCrZ4Nfo450Qo0QefQgX9aJGKYlSx0b7UeqDrEmPrQ4cW6Rld4Ubx687U2d
H2jlIKP1Cmi46VoHkmHQVONpYncnYbMAycXz4cZ2OtcMwExK3o8aYiplV51ZwGtypt+jNIgbyIiQ
MCGS4Dy0gqkzjLD/LSDITROlWJJ8plibzYhIeNK6DOCQNytEhJToJde8Y8BAMoIDdz8vjNi1FhWy
Wh8pfJV1TQxMPcekHeIxiI+9qgwBEUu0u0VyOe4F53k6woa6gQ1DEMfj4eKWUo7lbobMVzXGHQr1
WbZxXHTDMtSOnTPjLmVWBRmPl1H3oZoK0PKN54MlOgH7Txb4YlDTnX9XSYfu0ufWnyhYctRQUp9l
/zTI5wSKplI0wZpoYIJZM/Y1Rd9R0b+IMwM3OXMkpK6SAtfZy9ayE7Cg8QUt4vjVJMvjIhu2TTrI
0HL7TwAPJ/gxzdkriYGb3lDGrhgOuATMZQJYAuN0Mz0GeYq3+tZHcpD70hXX2UPdeu0Kb5FsIc9c
mCcB/z9brgTdin4dbb/ESRE2rAW4B6ST0c0UInKodW4KIwnnYc3CLlD/b+A9Z4yCHXF8e2V8h4AQ
SrUHG64FWoKIky9xJ9TGlyiDmoLuJ3zYvGiX9u8GcvNs56qM+4u/r07wzsykV8/TNhZieQEzS6vF
wq1b8y6QjUEbzgVvUD5j8jRYISUODBSwT9W7nkOfjAr0MEuzuSX3QP7HtdiQxiJSCPvUuGz+D/2h
eu2dENkT0KVDHLEmYcHm2Nh6aRh8Y4DNxGriedi83GoDvFGzKSXkhW7qI4FvmiEJJm8UKzLXa2ys
g0vUyX3YrHhpJ598GP9ywbayZpXgylTRSpDLIhh8ZqNiXQAJlQWhTUvU/jb9sAvTwnmoJp3r/sNQ
ULNa6P10r9yxqiIojeWvHxogjTWFGV0QZPPw9j9P6r6SFk3lO0ps3K5xHc8rp+Y6XDZvbWNdvtdy
zQptBWxSv8GVtbz/tCued9WmOs7dhf/6z4QeKpC2aPuZuO/AWF1o6EXffU2FCtWtdV08+90fnuqZ
oGmtuO8E39Uz7XD2RZ3n2zeG9xo4x0WCdbz9Z38OyEZTzGhZlfC6TrsRfXceJcxZmT7JwcUxFt5F
lKnpkZTs1pVew7aJSDCCVHlXJAP7bJWGoWWFPevnwEID5dPJ6A98VkuAuqhLN39Zv0TiOWMHahdP
bo1JS6el1Kv1AQwGMkNEzjWz/cB6IZnckHH4TeuGfawtmSXsc8ZJTSf1tWE3rGFHAkyn+tT5WYTS
gaTWXOl3tsMeoHQPI2FS4le98wD5Clo4KNtNK+6TC1J1H6gXW05jgM4zmbBNMH1c6ADuAQnb+QDO
0+RNkj6q9wXq4rSlYx0jkAvngK6rakbcZiAHZMhpDn5DH3GgMZyC4RbAW7IkhC7Onr9HCoeJmgwq
0vfocLqXKCIidKU4tKESgUEKID04ut1+qt5HlMUTGO+erdQBGO37ee+wyzb0So8HDXctdW0Tz9w7
PT0f/7hmZgIIvqCV8wcUv6qTKEUKRR2kfB7Hw4b5pLHNkpEszdM3ptWQp1wzlKfjR0UJmFTkVOFt
4YpJ7gTx8Z3sHxM+v/8VHzE6Loi83fjddcAmgxs4H1iapZsCB3r0GaKIZRUjWI8froBCiOxD38j5
xWhydxmsIdzVUYxJ7zZHII1qHy+0XP+c1H447cYEWaXhTeyfOJG6JFdvWzTqSaAyfE0CYmPDHkgY
1GPOJdi14g7GFhyz1lGTXoRYMEOlBB2UCBSI4adj47WsJYf96r+RfFpQ8Dx6OdPrA11adETXpjox
xV5OrpJ2j7BxchQMy/yU+jpq3jPEAUPPZHfHeCqaMz4EuUD39cVpFVRfEk5ktmEn1hIBayKoa6Mj
cRRLH1HDecM7CCRYe14SpBwpavg7d/NiFqgyvB3xYfgiXN5d2WGNYGLZM0i5LMy+N0c0CD1khTHZ
dpPb0jlahD2N1UgNAw7jnPnZM3+p2JN3WL8DUCIS04o81kbCYAHoEIA7XUNGcK1mXhXzsdPGFh15
w+Tb3GevoyLI7cR56bNO1uhakxFgvsYLqZWGaNLEo6hxL4yw8PJAk3Zp20GG3Qcqq3EuvmR8dWYK
Oc5/CAJ9jZyQdLpLuPVFjb99zfvdfHNp0QSvJDrh3OcO/AvCE9AVVqFQk33oLnKONdKmNjZlUEkL
knoiEMr9E7a94l9XBsaAfWzv9DmK9GaXAJ6PjZgc/dpPdAnM9exprQoji02fx8dWKKoqHXozSfKZ
pvyzWzXQssbSlDp0bUberqXgEltWvgMglXvCVHU+t9t02Nt81NLu+OirsGdJaMb3HBiGM1sX3ZKw
bWyoYbJonZbqmusYJ69t6639TRP0JjLw/lhk8ZOGTZquX/FGmi8D1K9/JM7eattZjREJ68ekRSwS
Q5EnfYA+w655GlYQZ2AMM3SLyrF+xI7GUZYCs0IZIUEbNsDPbwIKrWKHGgD6d2TmYT2iAy/4Ipgl
myXEAqPj+TbLVQAw3KJiOBAgskMQgEUch+dg6fQO8q7vghO+GoTppmJZO87ethOhAAa8Xieobr4G
/q4YA3klMwXvR7BjGX9kZs6jAiafhFJjbtLYdduAua27uHfkwA+TlcSNxn5v4msCfWldwPJuZE43
WWvODHYW5phptnfHAgeboZ0h1fh5OQQeVQz/akTrRw2RqpNggivn0cQyTwg3mJX6mlxn8e69TVQA
gXRAVh9j++nOBANi0t79PSkjJVFSwvyYdJyavtQymUHKdQ7EQR2khlMfR9eeG/Zhiy6c2Yf6WaWD
9F4g/H+9nR1rkYCcX2j11xiPIyu4tNoA7OW2HCKvnt1t2tI8UxBSEoc7ezN/DyG7pI03lZgLDAcg
QdDLqq/uDOqbWqNMB4DTDvoKfzSa9TtL6eWrivwnVcC0li9kBcWeY7E3vrvlqNPKYKTOINhRODsh
wtbdUvuaHH1ykFF8ROeRBd41YZHk0/1NCmYHcoG6EByvoedYXG5YAxGzi7XVebU1jj3j/07c3pXj
lTU7YjYBk/M8Uv1XzjBMQUYMsHBc575E0CHpcmseHmLCohIVO+Wdg4lL3sSP2Ce3oW41FPgtQB7m
iw1oA0EuzJJT3XxzsSBiWwi1E6FzUqx1tZqyBjBpXEWWkv3Bkxv1BpUMmfB3ldXcJz/tkvDJMxhx
ws04B47U+1sAD3naWZJFGGJnlUj1FnOt3Om1ELdCZnS/IV9By/6DSXxMGjFS5KLfHFoEmknlwchI
wfDaI7PrNBqQA6ZtmRrv/IJOVnLq8NESuoWc4TGhh1TaeRaYUvBYUjt+mfQnRZSSumGzBGef1jG5
NhnHwD3uRHMb8mmVBsNtthwjXD/0cjZo4pJruppa3XHlU71G5NXhzC8ks2WLRULDhgk8B6zH34dl
88tgsDaYH9+X8xZN1bMG2R5jEjtCA9vCYk6oubY9n6kqLH5WloJHakYHZHh22MGSllhJByxN2H/l
g6xmXWCpDVvMxLKCefAKUNm/qT+ImSaS0V4Zf2u1JRmWA8iz4L/EIH/l/B45FlrEdX4KY+Bn3Qub
pr8M9SegCx7flnUo668dU2r7tXwc4KfKTKL2k/vNU9sLTApNshrLwvmlImBgPlI7Td89uFpf2a92
+QTEp2HHQWcV6YIe6zrp/7tHQn8bEsCKDqUxEEeM59bQcQHTam7LXxeBpb12lOQOhPaUwKD4p1+d
vykCLt6qJbwS5TUhAms8h2/5Sgo061TNWHu2BFUHj+u4D7WXm4IZ3EZTzFnvQY5mXEbcaS4cHx41
3xOctP0fq8eiGORC8fFtfCWgGpdDfm/LIw2+X1a01o3/kYVUOZl55ByXLobdvb+rnOmoUmQewX9p
G8FBAqlftj6uQLyZsYVlI/qBfWnRvc6fO0Ip4IQUK2WPvgkx6YH5SBCGwfPCCC84vnNw8xXjaniq
513zIaH6F0765e2RpNv9Emc5OSPYf/17f//oHRrSLHvGrDvm5HlQOmMgtvTVVitHTonQ9suX4CCJ
lMDrO87DG+I1Wgup9wnWLti2QzAmI4q2UvhgEVDHqAdKx7CiAR3YlWErWHKl/lqQ1mGcv2q3vcEn
48FGllVKa+Mh1I/v17L6TbKhZBA/v2W0wHYWe1nuE2yyrFI6uYjpiA10J1ujCEOdZBdOHP0GyaMI
naT6WORjka9Fcg9iMmXcN5zCY15YDg0pUmI40nuOEO1RkNVCpb81Fwnkuz/mAemRZGYzSdJbe74P
z6lL2vQHu+uyBTm/xKzb9imoiWMM56C326kj3CCZdbjtxF7m+ZUxv6z3mcVgB0OmfX8YcjM3MjRb
wH9n3fbjeICisCSOugChc7CXx1/H0/5wypKVlZyoQPaEim6l9NWmB17OpaEBENVcHUfyWbbrkqlg
6trBkXo3iIlPktNWo1Z7R6zOkWOQNElgtifKQ79hf3pc2Hup2DPGK8pIxdPunaCKOQ8hNfI8yKkX
4zpzq7F/uDtjhWLyPLRni9dbNeQsaYQz0biKpBOSvnvBSq86OQ6MDFvmzQMr5Ss7BDTHeNRD1/yg
PNLR4lmrSIHPQoCiZAeEF3sRn49ZBKur6Qnz4nme6QBkS6SLdScQGcElidtnYCJiyO1v5Z4hD/+W
Jx+FNlZIiRVTwzeTKcmwCyx6pi5uoTDtXJVSrASx/a4+69ZArEL34ct0r2MSVSlQR9MirxXf4YzL
LB8Qtd3BvzE3mAKv9bXefrupvVOxEpdTW5xdO7TRNS+cEqs1ZYBXpWL0Y4V0UhDESSuC48ePCONF
jJ2OaWEgy4i28QU3V2mOkQE6ii5uM4n1FgFHl4o7FmI3qG3fb4XMzAaJo+nJBej3kFusofIcjUZx
5rEBIPsmv51G9uhwTTIqto88x5z43J1QYPoRa752RseZzynV7XJxKwkXoVD+t4JDsyzNQxiiT7Wt
T1685klbcJLi1nZA0hcZfAfeMXToR5+FI5SDuCdveqxnmS8IIu+GUlUoPGqhs4aIXIHp9CEvDbFl
LE+kIhGOCrBEd6/cf96HGKNv7lsKtJCfJv1LGAnwb3i4HwokyXd4SchWpHdoek20qBD18ocUp5nu
kI43OEgHtdxNhvdnqsMPKqt83ULDOBM1VzQp64T1lfsTarb+ov9UgcpcIVwlnRLoidcp4On87axy
2QftMKeDRF+29veqXs8Tsp7nu+nKQlE4QQgiJaLCztr8J+ghMEYlBqeasvbvJCFB9RMX4FIEBNqj
U7gIJ8r8bMYXu89E7jAfDJHbSmpMvROuusZZgz3vssKIQpM2sKhNOeyzEzanK/DsWcwuAqWHFoRq
qGd/N6BR/TI68JtgdGOAuewh0QugilH+b1FSUC7YGTItQ7AM7WPi3BDI0QdoqbOlOIYEifUQYbNv
sl8zSjfha21oBcZpdTiuGl3dhhe0shAF8eUMSeF65cdebmz+UyoS023FBRhuSkG0GetEbYZ6jNpK
tFBzLuFn5L+OPKexOLi2M1Dq5hE6n67hI47JLrYOOVAwnbGEA1ZRUD15sO7Opc5D8qX1vezguIU5
0+adRNDgnl1sU9xK8ZgOOO2gZQdzHkPanBBPdglgGqkWx1hqp80gXkAHcH81DSqiJY8h5TwAAqM7
ZGPwBFKrydnjohyJ7j41lZnd+6JvBYkxtUDmTqKBcdV8NTM/C0YAN9ws1/Uw18bPJrAK75vER/0y
jrSXXsgJfAHitHBLnkhiAuh+bYA6esK4ACij01t0v2FfjL3np+FMI1bK4bxxYPUgHxVbbib1zD9p
GUNDLETvoRZLBpP2cHVnzbwR5jaTfcAkw8rJYrkjeAerLH2ot7mSIbPvmDSgMdnrrKwYzqfQob+s
vAab7kqcvCYoP4pe+sA9QvHYtGQroAHTJbvnq0oL48FbJ6UUyk/eUC2SPuqdroe2lUMU6nSnANiq
PojJxtit/prcpW3C5wuZcPRBQd6uZO12/PGpPStYRt+H7IpkSrYa6dWz6Kh0vp8KZJJrv4VP7V3q
rxNp4YBI4nX7HR7HDuGgCs8jl2XszQ5iBJdiOYSo8lldBx20mKX2hUrdbmikAy+le5XShXqzzHnK
qs1FX49q0UyPiD/3NgQ9s28C08zbYY9NClekSf3IQ9Wj3eWa2Pqk4e8AB+xmd/j+6hNUNQYHPE9K
D6FLasCI4d4si1S/3EPRZYSHhp/i3kjRxUntQLebebXPHidKPZTGVQu+zZaRjJQ4HW76P7rVq8l8
LObDDklCv4BUDhV5xIs1BdCrZ34ZnOUg3NsOQMLNfUb4yyiJ+Qtt8n0dqAC3x2Y7wzVz5k41pKiv
uUq+y3kwnUPKSQiTvaOaPyyGKVluQLBxL2TSofjR1hud8AUOHAJ/6LWnSyz8rBv9cRbhYSsLYgHn
kJ92q1YiAMEIIZhKIFnrwS1CxClChmIIKwWVllwBxrZBmocF/2zHyw9w1BKTJUuN7pFsVC7kLj1F
mTKzRexHO51gohCBmOnsmxxF/Rhz2v3NkzNsi+i4cxOvq3mXv1EU0cHynwy2BTG6O1n+Lh9ur0io
SRPE4C1a/ZtrjieIkY7EKG2L8d38g6pkKDd+XAxX96hEYHk99gjdzmQfeDxqcdlbqciLYxKisMQP
1S3jfMHhcYizbfLzA4fV2wGOkPP34aHU6HJp2rt00HHuLsq7djCqrFSA7VVqOMh+RMskRPC23S17
BDdyj5XSof4hAGqiXC0ky1NaPWtRgxzPnB8mBR4WC1Yv8ZRFq4OWqKdfVf6lZFGfU30fDL3ZxZk2
3bK6GzmmCyl8kjVzuzQoxTgkoJz8oRl1My0rB/uPB/Jj4yA4XSLWrCv+U70EWuiA4K2Kg/AnUcM0
LOQ5zMSu4YUDHbmPnQO4seeQtnW2xokvYj7sqYVetQMKsXdsWuQPc2TF2BJlmmBBrv+GUnPjxXZ9
fWKYrlk85oDfpaq56hMnZHWWNoMfejOgg/umaIJWYFTOBXBwz4rSU9K3gaBAISjWteHeU3K/VrMR
N2kLgWRhmjyLweJEc4UvJokLFjnndUKG4klQjKdF+3J3zdUslZUeIvpKX8qu89htXDlHQbBc7n/x
dckJF/8fLNmFVjzBxkKN+YdjFqHdaPnwva2cQz9XS2GpuLZKL7KlYqfWLHErqTbGN3Xc46Z5KeM5
MedmP/rfSNhySvRnIVFT+lIW5C7SfbRtnfYeaAbIyWTGTCseYlgejGveMwjOeibvpilIAusvk2gQ
/X+D6K8KUUGku+CO9EGgMommcGYDm2sgpGXUaBz/SlGfuxGgy9lFpjbGrfx/5vb8o079ET8rL1KQ
CWSWHyKNxsN0NhfjYJS4qDcPrrC4Kjm56z7NR2/ISGC6zrKchyBTTUWk5pq4iixrGJAJB4L0F3Kf
AT5FalTB5BjfkdV3/WMkA++GQqqZNN0rjUZ5lOg8gdhpA3sOAxG6tK5gqUaD0qbEsgW+2mkCqX/h
EUGFx64TBTYAJJMAtmVomHkLGbGzzPd0lEY8tF9mDgK/eswntq/SSR/PsFGbPxRJVJBhT9yDu98h
UmhIdZ9OIUSinOmHTYw9Csb0ni1Ut/V8TUv95CDowwgatZxOV6kYT18oc4RBYrKWP2SALUWiDAV6
aBhxxA7im6Um26TxEJyFSxM6VhzmgAX7Db0P/ZOQbXp4LB4ode+OSpsFtggHJxaNmMo8EbmU/SBi
xj9M3xvBXvDk/xAdcuUgDftD3jDhU0xYizJg0vSIQdBPxLQBHx3C4+/Jz0SVGB51Bploq3bzNM10
Tr8wZhYYCqxOl1nFO3wbSD/O8bq1AR7jciC5i0RZnEeXbskVkvCXCshTbBu4JkaNugaQq2jhe3wO
t1wYZm/qvM5GtyZs519ibszOuzT59ABLdcYzpmTTGqV7tUQQOt1xlYd1cdHH0TRh9UUEAJl5CoRE
54KiO/8VzWYTQF3+97JHb/CLRb5ebRxYQh6ONIDckCTaynfGkUJeXAlRhb9vn/LaT1SFJB9XNxiv
HMLcq75rNo1/D9P8+M+eFOyNVar0t8m0ZnpUZbsGbG3dDkHxQP/8vGCmbdfaiRbTFSbp8numgyAg
03GMltEq/qRUnVr2s6AtU9w1Lbj9GyoAikOcnrIjMSErIlRwGjJhz6klBP7F4DMwuQfpiU+siwqX
0Mr+Ctbz9ApMO224xAslYbNl1/QuoTtqQvNa8IjaS5296E23GCjQ7jVYguVWEglLbByxO0YHZELb
u0Xg62KOIbcATABNNdOCIPHUe2FtRbJDCZCUTLtBTHOJ4Ubwl0HQN9CwNVdhP+uWXNb8Z6+vSi/n
pxi7KcHqf5jJyJL4DyUM3WyD3+B6O3WnLRNEbiG9erdpM7GXHltpc4YwmEA4e2SFx/kBIdxfbEuq
+i/YS/FHS2X6j3uGaZxSDY3m7LlqqyewgxQuCNHJbwjlsYGTWgDJnpOmU3zxPb24ZIL7AE6X2lQC
+nNncGonGzdV4hxpWuyp+ywJFCeaTcf921G3Z0AcithHG/LQHzN6u2mt5qJePiK/fzef+MA1vhST
eKjveFkSNkIYOIW9wNNZEErNRf6DRf8I1Mx4qIDqi5Foh7oOUAJsBujG0k4ftCRt2S/edNU22tkM
GQxpxK+rBzo2gjJrqGQPDhl9jGu1vSk6Adaxs+odAPsO/vLN86enrCTXjbKa2byvg/aPGgyZrcdX
4WMfiCSOh+l//6L+a2yOzSMVTd4vPuGHx0lEOQ/sYUfD3OsOvTLdD3t12VPnAJWqUdV+QCEukJft
v5VsqPBCdH/7egyLdzFq1IIoQLZTSJgKoNX+z+Fy2nJR3X/rnnesnMbQGCAvay1Q54S/tUISJXW7
PYkNSW/4QjhiLIxe02tqzS5Tx9v3WKOWo4tDzyUE9wVrfMIXApVQlWaY9OkmICQgKP/gKIbKOMeW
8nzXDF35IVWum2o42m4xME/qpD8LE80Hdg6NNVUeNV0UlgfnS80oamN8liOoVZBxCYLAYq7WHC9g
likK3aNbNVYe4aLMmpd/df5+ZA8iHAtb96V0DuUYiWZgwz/ZWNB3+7J5uXGinHnbdoHo+ZkGzxMD
jFrNnNfGzEdK2EWz3TKQaEZMDlPyVHtnbhO9Xx2PlsJPriU9D1NayW1AFsLEKY21SMzc0y9lSWtl
nxNEqGKxsLQ0xdnTPnQFWGdUIbdJaJINPruwxy8yJZb6BK9UogZ6/Ad08HgHv0NRYV4cZZlDIbXC
RD/t4ixOnoEAi9uxmiM+3mY1WUIm2B4V9oM9jemLgXfztUuvI7IwaqM4H+Bxj19BncyWo/1n7qLo
A5IMCNK7R11FfztYCXBAZfW3M6blRqs4KUNMaQnKzKL4C7rO3/c2Ipr8GpR1inlkd79vykomPEZK
i6+bl0oxP5YA7c0CLn1I0ApmUBvJf6708cn8FCGekmFbUA+rHtvuHG937WukDRHL+n9reD36t9jl
4DaOtpRz9Kms8GECpZ/g+AIVdqjHvJhOsAKX2oAZU6EnzyCccDLb8pYOZjpm/b+zaxDgn9bae0RL
spv7PbV71eFkpSD9kMV7jF/J879tU6GP0bdSx++82kCYMkAgioXB6hUoTr/GHftyAXanAvEGNOHz
tL5EKNHhEqXJ7MhuYwZflDjpfOrtPRAon88CuEpTn2BbsG8ihfyJIIYK3kYDYH8lFRGGdtFHHImk
Vucy6glmoMtejYOo0SPeds9Zg2gtBTJeFdWWzbWN8rp357t1WrkW0Z23Cnochg5tr9iLB2bxsIYu
vbkoo0t4X2qkEw6gk0ByZrryW3TDLhgGc3Ob6OfrdOecMlDRBroy+9L14dXZ1Ors2rUD9vB7Inlc
ZvDMvL53kWKQv9vxcZyUPdcEI1VtYIxe7d6iL9ui/czFzZ/oKeDqsVMWkMX/TjtaLCvJFfwI8Ced
s09Xc1m7aOtcy1XPqWHPLe2MEm8FDLwhgURVmGm/dFVlZNjwRkX54N8PUIOXz+flb+rCnEcKBRZX
aiPhdyMoLeDVTNSVidu/4f4Wh1Pdr2m6skLMWwVU1WRAhGQ6lnZtgMkdXcDja6BrlhlyNQONFYBv
EAmjNEipAiAohVG2r+4y79Y0aQ2bZcy/0O3IzYb4yAsDfioXxELTlq41Er97yI2KiFGKWqVpzP0m
w2Vp61GqwS2T+Qr7zV+hXhO28qAx5lxu/IjWF1tujyU3cuTJRNGpANMwMQDdxvmiXEQBIPCmbYLP
yGOLwU2d9I0U7AGic/pF+qpS4Fp5958UEM+nqBJIavOyshvnbS62+Xe5dMfNdo++VArSfllJEGPg
eBY7eqWsvi/u2SkAIkMIVeY1koIIo1XpSmti3QJ2AcKyMOZAV/6/WWtPedQKDEgVj5bgzrI1M7DE
0K97LuZabxBr3z6xk3hC8pPqJbg39hyvwqsCsKqo2Ifgiw3JYqrHGrYQWmcjcxFNrmMthFFGJG3D
Gdh0zuLxK7/XQxUqDlehCPeVgKwUtPig2uyWIOFCVdaoJkbxrZchPjT2qpr+PN8zT/dBeK9gG3M/
CvkD3St8YNtoBizoVrRcqO9krLkJ4iB1OA8Bvzk8M6qWML+UHKZevwl8A5gfl56CFvuacDqhMGcX
o62rb6SSibyt1lPIPUC1Ma6NUrAUf8PDWpPdhB5ALh3iSNnEzmI9YvUroZ2j+/RD/uIdqrThISk5
Au6NNVwSjo8w/mu+d0K8vnpxBcTo9+3INZ3pdb5cmPM3hFLnRcN44hu3W8/oGmoGzVCqyUMockGL
xPsm5oPvD+WdbHr+FonalTVFPsd2jX+luaFczNFEYRn9VC7ye6iPFFRA4NIlk/gd9pZBvdtSALdL
mPmCdadfIX17BX/Vf9Hh2c1pMPSzDdNVEyr0cy4H82LYZtgmk+yt0BQNXtVH9B+R5EkPUgAlM7ps
KRzW6p2GZKWSF8ogXLYqtjaFVdUXuG5UlMXChE3XOod2YuB/Xm1x9/LP5zxKghrc5/DLdW6Dr/nF
Fkp0Exuk9pRpekXDs5JrAsMBd4M6MghFZcOJ3crzDz4Q1AtwzktJdVFJU6MRSvGD6v+799GrKFaE
8Hdk7a9/FApaNLyx4JwovcUmAEuC2xijqGIM1IAoY1mVlTVgG5ACd0JfEXbX3XMM4pFv6zm3GYw8
p3+GukKVHcYVVgj4h4hFdR0Wu4pUeJ+pPwuk40KNc/AT4DqT4EmE/ao5ESqcuC9tVUqFSPsalYl7
rHV1KvIXMeTOOjgkr1Q9jhWnn2YaITVxvTRN36ibSR00mnWUo2lgIO5pviCYxUopZ232nW5t2i3C
XFm/A2Eoi5LfinWgGFyT1wJhg+4CcEKrQu3LFFmEirAp6+4BNmL8t6EkneFi9WAAqhUiIOTE1Nd6
P7zmSMblEgdKcq++wWVghxJXWgLkIf9KKHDkuyQKfduz8divLx9Y8Jtft+ce42ksoPh0nfe4ghCE
Raq2aGyWqttiTvSdqMfihtPF5Z925SEgORJBTgb09iijjLFDUtIMA3XsoYKEOKoQpMcejFD0OMA/
waExJG9u063/dN5Em/kVtVwtigQj40bjavyz5bsKpMd3LecUcMKCJpOgteVYevGyfSAV5LrJfEWy
fTqAaXaXbGiPx2Q06pSQE3rf722MATvZpcW/UE9e61lNJN3Tyc8a840WkQpn9oNXu7k0Wb7nElrI
H8CvyILCLEw7HDZ/9B3n25/joodL6MrttLdBrE84SwZw7wkLUzwKvSEtRYWCufmDnfxJpExyc6YD
SLA2E8Y2EJqJ9FMHbCOMzIyzycKL0+D2GTbql7AnLR6vQoMrAKq39X8/WAup8TeTx6Fyxz5ZIvQD
3vCZL6DmyITugkLFHrMY/EZpLcVLrV4VqUTyalhs8CuoGvkwTBMmp7g4FCYiEeZT2sow0hdBDZrm
dVF/WaCSjZvb+KXd3davYm6VKmaHaVhEsCzfC4+56M+3k9RMp8GYWESkSo9//HfLsB+sVlIsBV6h
ek5hIymx8pR60wJL0IrFu62tXtkpA9uvZ45dsoR2ibOdqwaYJJjozhaiXMhqu4/b5e7L8+29CT1a
Clvsw9MI2ChrjxfodHgPGv7G5Vz0c5dd53TEvpKX/D0qQEVtPlg9aT492EKuHBMVTxXoUdxBFMqP
Q8lvclOmFiVrLVSfyaNdy+ppzDI4j0KhKxmCcHdrjaRc0vsJR1Z0gYYLV/psc2B10f1hSfsQZiEu
i/NFAf89fGwOgO2QV2hyjH1yhB9ePPd0pusNzQ3j/x2J1p5u4YEZpaUOg3WsFpGf+hBur7T5hrNV
8va7peq+C9HAC/4UwofScLvUy0wU+mQsqJTHOMP5HanZLj9gwil0ZgTQofh23nQCptQuHmsAcSXA
rwmBJLjEvQSFXVIH8rMxQyeyicfQk+MT3NCjBSu8HeXhefkRTDmImruasGZrJJlgTVs2Q6+JRoEU
KGmIlZPVqFPJ7wHd61BiVa/bxSU2RTXTz+JggU3ei2zBV/NicC5DT1JfjdFhPUJaqdvgZ9GJOfxz
o0qVLeGPI5UP7Wj0Wh+kwbhwkuHbHz4LVplp5phRBKfz0iHVqV87mR7DkBUGRuGCwBn1bPfZTUiL
e+ILpsgHzE4JnVDuiGCA8fkXV0g7hrtjSYsQ9WqulCVu+39TrPypRjG//Ie7VeOqQZLzmPe5jXGE
b6yvNr7pn/DQF8nKR+q2col3lUo+0IbPRwK0RiaPpLaR5zls2XbG36mEQcFyAbUp9IGeDhQBQh0l
53oKiEDE6EX3Dhx4Isvf2M+U7gw6Xeq4C0cVXQBZhf0PbPuSFepeXBAs0djJFHn4OJJeAH9aVhmg
S30Jlf16Joe53gaeRFZOfDEwT19TIdvSyi2nu/h2/6cH5w9VhwWO+t+ja3IA1LjU32ja/bdxadJy
UkgMYFRFRSMxfzk/nrV+jA2D7iTWQW9CXoQE01vHxZs4EipPhrEm44U2e2fhYAHzksvgxRM+p1xC
F4GdWn3v+t70l8eJEwQT1Lk/6nfPMJkYNJwCAcULsX9Vff3yT1kBwa+PTTLtACyXHDhEQuNoS/xg
lKj1zVo5mqjCDwQCJYXs1LD0xoIxW3G7eM1d8wq5c0MLaX528tuqgHhY4UpIT2A43VW3fexW2WVi
4rv7mLKrHEvg8Fwux5Ott6YbSmHqk3+PRgSY6vnz+UEiX58YxipMRLskEldqA0caBxj+Uo2kHqtk
JwX0WeVVSO04k7/BSgBXxTUeiXYYyEI8UYDhZxgIm1+0w6a63aFvcTPfDJEzKKny8liLlz9W26Bx
VPsjeiMNtEtV6I+Qwzya4wsPqGcw3vMamcgdiChrlI9ClRKTqd0uHuwZF4Yob6UbVB6JG806PltT
8lfjAgK0hiKAuYixkQZWrMH4mX9B5bOLYWb5TkCyIKbPc/TGGb4zgwcJX/9p5AZdSFcN0mLmRmAJ
hUDUEwK2JbNExkiYrYhoL2uDuSGVxe3eCgp1r2t/deShFo8QaEeo2vxX6nkoYObz/7nXBl0sk/HH
QMcg/GJU/GJBoUmhavaxhjxKQqJnkwlb+hy7Bu2fnrsxxXD4r3iyRa+hF+5pnvxgCaTM454YiRIR
Y0bVNwY7rQ8JyQttZDdZfxxYc49FWgBGQgO4GMImOM4ncEKD/61/JC95dbbHqPZNnPlbKJ1RKePV
tx+6wOL4SLiaCDO9Ycvivw2eBa+pSjkZP5ZAL1YCmBXi5eIawZFROqK8cqTv84PClTWkiyAmu1Pa
qPjT72SctIoIKDHxWbnvscUstyfzcaO0wqUTBSTNxFgcqtIuIse0ltxgBV1ZL3Pj52Rb68wJ0RAA
he3pGPx/2CVhIfa12ep/6tVJhuuhl5eZY0CsjgXh3L7ctGNb09fUN2mGa5VwkpZX2voDSl9bWDb/
VJsHVMFaWID4Wi1fnOQTQ8KwDAIfe8s5FJ2fi8+uwZ8RmtEhh7K0vUEPg8kisyIkjVW3mnDt8iBF
IkCoe0EoW3qEDIBIN9xbefR+BpqPvDLSb/Aks+D5X8yGCoYxgrIyzVpE1A/TiCMgjxwwJ1E5EA1c
lmGWqYZpro7yQoVyaTY7IPY5v7t4s7VshxmsT8xO1Si7ygOcM9+Veh+uOx+eZiBHzqSNJ11x2DFw
I552I90pzOpa5v1V7Sgq3q8SYfmgyp1ShMZz6gydazUHfZeBvzROjpaReBkrqAuN8bAdrEiJI6Vu
ADY3ZZ02ABHVArKr9zjTFkr/l9R0r5/Bx9yJTnXTzKt2pzGPm5jAzs7aDCoDx8PcCrETheCqk8fq
DyPj/onJHDPrOkpsMncyB9xHaVOXgF55s0ZQjc86DVFvNwQLQ21UQak5oNJrZG0eE+H1KyPEmctr
ZlzVQhqs/QZc6XQlaUmKcmKWnPlE+9HKgxIHMOmGFU59BJpwg+1UFpWgV7wVgqV6LUBD6QJf3Ytz
TboaiX5oIx5K1W+bVgIz/6bNzB3eBp3JTERG8BaNEwDgRgwcYxpyYgd14H3p+jtqq4M+kqEWpSET
iIRcGFimzhk0aPX9xpJOWmqFk1dv22sdzOR2lCfgAIoNQ8UlI0jmkSqrB9MKUcHj3O1itvol2BsS
vr/PGvBHjahc5qIZdoQQdp2xkxiX37Ghrj0Mog5yjB/Blu2UJsI2PTQWa0JSGDc5J0r+SUM+UGQv
DoF985ThDUm/01cOq2kTGAlB2B+PbKZnPRQbrqaMyWUOXtbvh8EAbqp0T0aCT+8qE5jp+2eZpU1S
9FuLxbaMmd1s8dSMyFQoHZZ5cBiFQZnGcnOO1ifYxrW1jTvG8mLUnbkJyqnspl6F5LEpQqFmoSWI
LbVO2U7BUojdpcVeVFHnO/Mr+4dnNR4YJmJJORmYSG+7N/oEp2W2a3BIpT0AHYCtTtAB+wXLr5C/
6cR/Q36D7hLq/RjD6ZX01/AXdH8AkhaCVsybRqpb08BwCq9VK3AUCpb4LK14g2VRnQnD0+U+u7IV
hMPfz0PYmwLCXdUFCt7rD7Eu0u9fOMl8SGG6RLODaVN9VTg6LJ4IomsedcGGxrcOJtXBkVGhgK5m
yV/hISqRYmg2CTWFDgrelnmpETXPy3+hGW2RN940BO10u39G32u7YH/gn/GBNB6CQ7SZ9SqwSsaV
CsdCYBPHeDfgGOSsw0PytnqyfeyTIgcaNM/YrZCrN29d0zHYGZhvRhe+tXvgir6I4UWkDg4aYce/
DYkFPW97JiubH5sozGKpx1zcJEZEBPqNZHVC9oAXlY1hvqB9VcKekiXn9tgFAkzEIccSfx8aIQqN
ytU8ue0ECnGD3DfU0o3Ss+eI7oPjXH/ZOmVHoTqC3qtzfDwW328eHH16SDwx1FhsOr9QeWn2C0rw
WlIlq1cJDTw39DN9qY1/WZSLCkp6m/LycRJLu+4JBDojfdQeHtaHmwyW8rfTr4FkUal4/N5mVbKR
PTT8F4Z+6nIu932hmRGXRMmM1oKYTjmb+y1b6ePYRWeLhlz0Y1K/uiADThPH1NTx9FKzyNv9O4Im
ICFQccS+fYTp2ZLNDG9RQ+gANa6NodsCIFaeAiNAewdN5Dpb2rmwOCx+KRQYvBbkzXHzJKiUjsTm
YTH/U0g14kt4jxRgWa8d0CQ++y8UMDFF7RCMOPqtaqEjW4t8jDvv3egScrNhcS7IWpH3siGiIw+V
aso3OWLAvaZjZxRQoyRK67r9DWEV84ak/X4hhftzApIM1CFZuUu3zu4zDazmc8PX2Nx/bbKFeSzt
fhhDqQ7w+Kah0htviBu/wf2Fn/llJx7r63NlBX1/t99bnZ73TsORV2LGonJkl5EgRTmwEgvxzXEn
R+QsDw4aDwFOoN6mamVm5y0KX2cOTO2XQ48JASvwcs15RHvg77d4V20jhRi/ZFIyNnorX2KwNlcS
aHJOGlvz6038v7Ila57y8KE8iKnWtimSoLhGw3yLb7D9Vxt1yPPXzD8nbalTJI/wSmYEseS50P7F
ekkaZRWlCUA1/ZE2070aRrv3EphcaAotviBsRdyOnP2rmpnxfa3HcQ2GmhLD8WyaVztA4vdk3usw
Kc9yeKgCe2Vv7aq3vfymtQgFeiPzGcS0Tiw85OcHnkUfMZ8lE3gHZnQKJ4/oO3w4aSbWLENC2EVO
91z10mPXSP/L+YtPzGe7GL/p5I3h4uMEYPB0U3Seq+W4vrStfxb4k9KSeKfXuzCJXlygV+HLWd7m
8c8e8XfwAMDHGBNbW9Wjuf0fkdwmPyfx0lXO/aYTNd/+jnN6IgjI/bJB/cZ+Pg1NZlOLfBK/VuN/
2knsMHAYXZuSTgnzBnWVENXmRl3u3EZIZwMzVNXIRQMPN8Ksf8sDN1MTdJ2tjjP4esgr7srlrrEX
GI+HAAPu2bpVkrHyhIgXQl2tcmk0iIS+RcXDABA62zhHGkzg3TvxhYsfGkIahTYtqfVY7mqS6FLw
OCcUe08hvJLE9YUf/KSMzjn4elcwXntmVaxu+eRpMg8qhCMKDfFVRjiCljgMYgXxkJDZPOAeZled
zbe0g5XRRTapGmVj20jLXdnWsCo59rGNqu8JE/1QPd0enHRiUvYFJNP2Zzs83GCfN+Hsuuj/Vkv7
+lVaPQ4AhoIrKnei12+axciqx6u9/h0tuQ3o9AKCxyXtZZivkdMtXJIYf6J2XE2kMq2jmVJOg2n6
1NA9UMamUDEKL5GPqtzEhpTNfSwu7FU2EzQW9yqPQNE/hacEydokUmK3seydSHxrcRfx5PLFLLxC
5JSwYwPxMkIbS3qDG9WrkVCTVQQxX/aiSNjSOfDsvFIxgiD09+cBHlnoIPmhLh4z5ck56IIoY3fo
wyxXgejz0aX0lv+UnU+Y41he3CBLgQ2e50nk61YD53oiHdBQE6x+S05VvEAY5kZ3g7OxI8WB/GMu
0c74m2AWd+BYzPYwXLvz6rcmirasrhl+dHwK2L5wzPIvU1M8MNllOYP9WHx1cx+5BBrmAe1TC0ad
tn3QXcS3gV//49RvJST6fkwm31DVR2qxUFXJk90p+RDtjTYRref8eKVUQM25KQJgQCHmlYbmxIpT
/C1eVnu+t+UUaILKh1uOn6wPCOGIFgv6VVR/lZOKCShaP0iSTZ3mwyMv7gvTwfBRm/C0It3FbkMK
AIqakR5Y3+fISHms0ma+8XfgpEHISnsdNuNhapZj/C57euv6e/F8BtZnA2Ck31GuAjClkpvkTEWx
ua37OjewnC+1xjMgRNigTDX94lmQXiDzYoHjc6a9o3hbbntARvJMd8XIgfUlemYI9IvohKsleBYK
NCsN+BraVBKYvc78umdABSN0FizZyAwue65ZJf5SjtACBs1yBRX8hPm86qSzbYeJRXKk72jE7Ddp
r87Vcl2Jn2KgMxJ4LF5LAjDXE6utdbND/yfEOlJMOD0aqYRxP49wnjYZouCY+lDHTq8sW6IQdKm8
/7oevWkOlYELcv//hY+o4KOizxO3es3Iqh3RJJZfz28IrNGhy5DgSPFwT45AhLIZeVOXNxQcS8TA
nTeT4W6zsQOzF+PzH4Hd8Q4+8JQACOXUbunyZGSmShHnhDydjVrgxIxpA6AXanCLVLuX9R3MLz4m
4YU0eE9wR+VpWm62I3+ANlpKetLSMRktFTWkBS7Ns7kpJKXqhnvAyLK5CtRYBV7EgLz293TBtG3y
bcCAddicx8Z/GUx0H/sYZsvZn3JEtOllX6+HAKIlryusBGiZHNXBZQOSKtF4osdY6eiVslEI19ZG
FdQCVsnqesuWccVhpdGC1sVO9EAh7iVdayqnAc9JhFhQ9mYp3o1T/KahQ1An7oWnELbcAw1GrYaa
4G9M6XD8GMFAYY9GJgNhq4nuinSdSJ/Pi+DaZ/gxsTfN9q9qCwO/HReLpxtygFaf0hhlzgEZh3h4
9QYyXYy1tdP+n4jjwCG9XWApW5u35vln3CgpfQ6uHs29nUetVCRcKTSoNBuOSAX/EcEe9kkmdjgs
8q2Gus3jouL2PeWHYRwYqDtCIqxVggy2B74jn88wtS7NnmArk5/3QdnTpEUH3HtW2d4K94g1Pliq
acaaoFom2Bq0SynqZ9pNoRxuJA8Ph5c2i6NG/fPxL9zlINakfiTxpACXtkMTnQbC+7h1mBnpVGhf
M6tQLLCWZ379pjXkczNig9d925aJpTyL4mYso7NEBaTaaNAt9dw6NunCwEUXnCuIApOAZSucrLAI
TFcFizaoDCK2Dvy/Y7miwx2oz5aKMgwIeAsyzK7q6TwkARajZ/3qjaiDe5I6WdEVrfUaB9oQ67EY
7obma/6NLx7VrsZzFH99Ll2FXyKcoE5LdL/spO+Jq8fzUYRQRctq16quOxAXXFQ8QN16LGlqGksK
0TYKT7dI5qxgHCV+TZr72TCpC9ILJlbEbMUAdhF/cHF8ODA500JLMOQPjJPIdQ1wQYZ+Yn4z5TcL
R0CXMTHt65kVG0hdI79+P4NJ6NF4rLXinVw2/n/KupdEXeFdZBDCSE39EGC6Sl+8W+KFRe7j+e6g
iuTvfnZ2XL57DFDHwDXXKvpT345DanDUxmoFpp9PGIY648HBcFWlJrR+kjZWJytspvze86zzd9rC
cwmBH6hma1nMBHgAVq9gkTxCXZGsodvpmxE7HZPGBEwRC849VfCikBxAW/9f64fk8fOaXdk31s7Z
UIumHwdjcTaZchbsAf5AamRMPIdHaaW9fgNmaIIQ72BxGk8Wr/oC09/Z8gfvKb+mJPDlq8jbX8F/
HVk/JO2hdKmutRA2M8aOz+G0ifvZ1Z506ID7mwh1i7Aw6IKAt/FSPG4ZRMUtNXDgJcKSCJdGOA+9
sguIhkpqHUTyICmpccWGz9mDvYgCHO13hmTjmGp+vu0PIkQdCIocCrWAFZeOZTpYeoEwFBH1ASbX
EoAYf8x10PKSDieQzRtJyMd1Ky+VLYo0pV14fgnMVTI6iaAsxMTh/682IBZ4wCG0595N1V5jpHUw
EvQ45sRAsiEs3jRcn9OI//kTSCj9LnvMDdsmxd6Lebv9vI1vqho7rUBoHj3rBNCgUi0EDIWE+N+m
MPoLeN7KYS1uf1ajdLSA0oL/75c4LfduVzN4qWjLoPhN1TXOz8G8hOreXvkH4JLT/dE9l1AdM2Mk
c4DLNG05GLhQb53EWayuC9msQW+LpNRBatYNPhoR/Ri65LE56KUkn/1SjZCMaaP4yetuyVxHRuMl
ecwSRj1ABSAKEobJQi5nTxBtEZzvTlYnVFcgFDlaO06wlzsFIjMpcSMYNDLE3/XE2tgKukb48kA5
xZSRiNv/i4WC9kUFOqV3KyvQiwR36g1bB901RFZCu+nffOMRqmGvxlhj+gk2xWGw+DxwcXwZ3pEp
/UPxLcyEwO5lJ+Y1J9jx+JZVCH25ZbWuVnWDbjGwIvqtWGsRqqfestyqIO2AvpspcyzHAHl5xvq5
mDsuNdEbFtYE1n5zKJMGYzZ7Jfl9z7/lfA/lkfdGBLyW/tBhMJoizE6fg1/tb3TfkCbXngPRweE3
M9N35nKu6PY/T8ImoZBLQtIbq6kk/2Erdi5dkhtSDel0KxNKm7zvTRUmocrzojPuzbRTmFMy0Gpj
qUkJDWGneB+vGbtcK+5FM9ysTvpSP6q/lQevFRo1DQBrf/VmvRv0dCO2Uq1ltOA4wfk3i8R1YBAd
NFxeRtBjZ4bbbi0fPFmQYGFkj42ZMdyCZtEjc22nX1INqRr5BnyvqiylMgcouwcHaTfhJdEv5lnm
o+hVUYkE5/o0n3oXS4M/9sC7j7q6WO6rTnwKqZVFYgYD2QlX8BhWON8MFk+HN/h94EV0VgnXpGKx
iN+5Sc63WOzuw5EbSmdolZPyQEj5TRuP/xH+S6H2STYozaO05ig/myr2zoeWaOKV8Z/TTYC3j8NT
o4eYft6X/e1uZ3G8dQOLzFxGJxoQ+Mwe+cJpXQ6p1zB3Kw2ZO0RO/bkOyPFFTm27ICC0oGbQ4gne
JsNM//mat/9muR0KODU8uKIwjzAdsIQ/djBlrUnCi4kDCLqbALuwPOUDYbdqzTgdsHAc8Yo6pQDl
qmpf0xR83uTkO6yU00jjKoOlBJPhE7T/mWbm+JgCJ+f+TOpboUmCAJggLwzuoAVwQLo2FBVJfFyf
+GxkieYZgmdu7GzfqB7eCyMRIhYOvmRy5w52n67rQrUmkwADoIY42XV5VR/1l3aNVeUUp8HsmSKF
Rp+xPim3hioptBUPnVZxH/gTftmo4Y7aRIhokzAv4hMzxNLjRmiexKiSCARea0Pwsfw2yUBr6JUM
1gI4/dGNNLyW1nFcObEwiKwICiKLnffrFiKa3e8qz4YtlhN4cUUVw/J235VpnDPk59tz7H7NPu9g
R2S0qzpHx2pX0GOiuyzfpXauPt0Xna3rCwRNUbuowX0r14aRSUqA7rM9SErSic1jp2JEvPx5uH+V
kv9zZA57Xpau9vYPsq5F6rynB1Ol4nsuLka79wq8V4iGlQbr2Zp2zI7A4fABSU+CWQNAiWaB9JWA
K29tdXxv5xQ27Wqa8PBmeZlPdLfli3xpYzdpslE8B7ce5iXx9iD87LrpUZbvCF6IHJIqXt/Q0ZTX
lHu1BK+yrS3DV0Lk0mPH9prw9HmiyoPxMuKRRelUxF8cGyuTfYlONBZZU9StOdrBZODmt62zrkLT
bMwUG1xvliwqBMrEiX1ZJtPnYQYctq8Kwa8Z0hkcIR+rOHE2N3WoWy/1S3cVY0Ugzh6SYe1eWrjV
zwAotMprBwsX/WELq3eOZceukUZZW2G7jiBDD7q7X6lwio0XiRfD6v1G1Dn2MGhxPcA/XiteR9f3
rTRUayRY5QFyO9tIXoPFcAnda/+B5OhYiXQRi75F7YciClqjC+P4YJszkth5HlA5AKyTj5UfaZba
xfc1yj7rGCLF4DGajL/F+unM5LG7KCEJ/UinteNkGR+mUlzfMHPL0g576NhkclQsXELuGZXdtVc1
CTQIHn8vfRuDMkzP38Ru9xbSwePlWIexccvZYbx+U1cQIrPSr797Gxemee0FVm+gG0N4au160Od/
p4TN5V7ucOqypoD5AUMhBV5xDiMt1C03KqPpYEHuV7hfqPe6Ja3WhrT3thLAkdFhxOXFRugsgkK/
1YpSFdCv57uXAeHJO3cbeaUwVG4xRBCBtB2COQwUScOP6dKaUr2gI4+958v4J/RP7/p/P+qyqY+C
r6/VR80E1UykGTGxh9NJzgy2gAVjwn+ao75ymPsaSjB6IBEVHxNf6sqedHK8GYbsTZ+uw/NLeiws
mxgnTEZWhcLNe2raXrMwNGWDvToYcnnqDG+adhIE6kSIV4lYh9iAjeqvqOeAt+i69UmA50pPIBsZ
y59361SVHyC3dsmBe46q96rYtuTvD5HlsvHq64Wxtc2fn+C8FN90Ad+BN2mOFPaNVesfdaJbIta0
DvOQI9qszxZ+P0Qo1wKOosNDslVjKPsFGsnDhGO+2ru4XD3jdisgrhEpCHG6yg6fKcr5IAZdP631
Lz+nqHDJKHpU6dEhrH0Vp1Y5V13eZW4UPTLTiIdrR0FHFZ0yhpKRRG/DLb/NWmDfZ2+NLZl+/IAm
2wI9MzTHFWNEAI19weA1GOF6ngE9xswcw9j1gtkh8cCVRg1+PKVAUAdta40gTeK9lPi+5wgMz5NU
AA3QIXLXf+CeAs2roRFTGucN2Wmhyv3y/MMMoMp1Ec+FpIVq5pG9cmeXbyYKsZ5wTGDZ30LZswtx
pRxH28z87UgnBJey7Gff5hUN1SxOdBfJBxVA8HzdqI2RCIJVhzNUZBZ6lODy88PDT60MoS2n36fH
DzOJH2lNrRIknCDKeog09O6Tcza3LypxPQnLHOh4Xf8tlDfvr0b3raoIX6t+UeKUSBdyC0QrimBG
rQgDbF67DWmxBO50F+8BZJq4XB9mFaZgtGYe5p5kxymzhqSrJZaSxzVtrpwikigaKw3jLJDtjUul
6oAReNpCQrka5USZdHZZKPOaPp9r8P71QInl1mcg5ExvVFWvkyaWEXOvuMvxoHtkUtgABpKAPkYm
hDxG2hLpUQ4XmbEDv1OAnU56Fx2HQaBG4P5tIa/qGd4dkoMXkTOSsDUqgUqOf1kiPo9A07TYnI0K
98GFGmUujBwDZrlF60vL/SIUYgFQVtgCoGxF8wIObqXZMkR8LCTRM6wsIxn5PtwtXrqoUEKMBFHP
qbPxWTMtpsGUCqwUjNbyJPWlAFvXhFji5rKdpyyqFxVxSdoIKE709YtqOkzV6VlHrPSsEDJ6/DAj
RDJLbH06eErf1JI2j4bYwK3MQLsnzShfDDtKTq0l8qOXEyAekc1j/hHh058YIqigWbowU2/ZAxFB
B5yB5HE4+s9ZOUM+sUO7FEAelg/zuj/GwRzWT7UWipUwFuVLHBXFzIg2HpDXiF6ssEklxjuZ0rXE
idvV6IKQFbbbZnW3Y56jYWGm9wQb3iGNtq9Xp4IhgwLDciPNrteBhoDHsMkVkpCO99UQ1caoeb3L
apNlePtgPnZgyIzx+PSonpMhm49WMzOYXTPKWjXK5rtaFP8awfo7XbAlWO1/60qBpsoAXcD7gbzP
EwmsnM4p0t9OUjsAlRWx+V0wE94PN6NQqxhKu0nUMi4NDX40ErlsX08H5UG0O/n323sTEgurfs6r
3+ow8sCcXQhxodHifSmchF+Gy6teBFI7JIY4D/O8X1Za86rAwZK+84HJYDt3frCMGfCYIkwUtMs0
YGi4bTFJWyPRTkAgCKY8fOIlJZTwLEy4eK9ZmompV2YCpOQ3VdeqCOLOmdZr3rdFwPkFPLnf/UHp
PsBtGRRQjiwTAGgl7NzM+C+veDNj8Jvzn1Y9Ds4wQI/0Ek+DHKQjVSLusY+C+KYxhlrlW+PKvldt
m8aTfowZ9XE3y0mKgUnCB8+JOw/CZp5j4vznMT/no5EMw6zXVSCO31PavTBk1nzg+mpchM0Jk/Kt
hlAtq4iMcKsqWo3l54Qs3sGLQTb1Mn26rtdkAN8Ox0xb0qLkOEoV5gGUk21vGwQA3rmQciqWdkIw
4xYe+xa9obX4lthMpfcK71bZD7mc45ew7o1ujEi4yB3y4WxRrDnNZoRl3QRaz0uAI2LOVAHyRPxu
fqczpMj0PzWauRy7jWrKbHQz0UmT3C2hNiS4i/ys4L8lBwCwcd3udRn0n6c/WcEDbFgkvOVa1oY+
oclZhpcOR1Z8eCVK/e1lV4Rnd+wss17HBWs4ODVLH5yAj7sTHjxHRiZSa/hDbVVZslwnSrKhyw7E
6ded3Tv+al2hg8+QR7tMhO8qeXpsXkzsTGBaMiDaHlgCVy7P9nfbyAht5x+fxKp9+lHQyJs2bOlk
CoViYCbDc/qIJAhW91lf/DoO2VFFsJf1gV5t8mHUlbFBWgxOwsSoysSZnHrMYLdG2amvGiDLII7l
GITAI7CKpZI8TiXbRj68X3sTOvFM5Cp3RjSqRT4g9TGXALLdwFO1zjC2cgOoRHQDlcwLfTdMcfx+
pT35lZo1LScKr3e+sULI8ARBuwr5BxSfQQBP9Rj6WxZpO2h7CH762IrcEwjF7s8hOk+jgHEAA/XK
MgllKkFoMBahAXnyM+osHRePiwrD/fJaM/CyAukrnkTje6gZJSnaw+HyFKC9SQrXbbpw0X6HbFci
1/8L2bTAKMMYKTRPs03hNUiMucKToqcEjC0Jjr+oaKtkuyz5oK2amvp5ci93e0RZm8hHueqgfxLq
1nCEdIW8Aw8dAM2ZNqaQLJ/yky33zTImFG2ejoJ7UEtbwj/5s2KQssMqzITNVIjs3T5J+SwHq0GH
6OA06CZoerrZVseAeCQOKTDhLjYSAb4Yx/Ry/c4ge0k4jqrM3yHjrqIxf2LSCJyBi2FqlVJJMiZV
VZiKR4W0flQsfPYKbWJx0HiDkfMRGXGtC51o7F4zK0ixq1AU34B0CbaddmHjAoFqueqMGGwAg5zv
GD2p0TTmqjztQcZ63Fh9RVvreREvV3M+AusWAVPRQbre6g1M/ewdUoL66NhGtKqbvXM0INPhL2/W
zFoOReOXYD1OrkhKa+2e7oOqb43eG7Px4eCAL+6neLLwe0m47SneueU2sBp1TYADZZamo47VPtqA
H41tjAFKUfrrimDes/6azcHmOngKSz0WloEDRnPeOKWSVRqwgbrYP/hXoxSp9kZ0rCmU0re56fIT
GYpDM0Fy38cmzKJ3MLOxPDuXOLZso+ud6dQlGzaI8+KQhLZCpNwYXELo8yAEMO9grdKZepEigzBF
CewNgk4kygy+mfkXEAdJZEO8Wi5hvWuB4N7Z+L+qBJwhSn3ZppjomfkMaAY67plNz6ThSw9t/fmH
ADV4vRGiHgxCddk9ix8zvVTEjcKCYwTCxIpvm6Zf/4kR9Qb4DWROKRTleAthtevUT/l6Zyg5ofiK
J+/5Fb9jws1XBMKAR8BTrCl4GR2Uhigk+l7x/DaZGERw/+W1oavhelj5LzwTjRaWe6Emf6hs9boK
WpjiTRi4xqNMwWWRLi4RMUn+qDWFNpJhW7jB4SVlHBkirIiDJE0X2CPIsNeDlDIo0bPmIR0dXrQa
GtPoX5YoHwEaFaI2QtPsW295GK61zASqHFo7nHdp+fzPUaR+nXEHVqmVPYmqxrXvNC7n29M81Hoz
9fcdgyW5CFTPj4NixrNoQSPuPfTRmBQNu14en7rMBhqXU9W9SCiRn965L0hlco/GmeOf6blb7PYY
2kRSRdcd+7TYWjgpcbxk65yBuCGvfTh6XTCdvfkkz2Dt5yLHDmGFwmb+HFxriQFoReXrL16/44YQ
wceaKd1JqsbJ35GnPkBzFAXEKUUBTLYCAbDcTlpxDW2vsdDBRK72LyR1TYotT49sXIUQiPSQkRxI
c7YkmDBEqW0g7ISjqnwrtri7T4BvUZcSn/UQwiiKOmd/WMaTSIZliSnrBCmcvg4PpjYHyBhO/j+y
bMC9DxrSwiNdC8t+8zVZ/3dJUmp6jNm30WoaOWNQW1N5mRVYMgoM8tIffIdeAhehTFvsHy+tcAm5
9LRAdfshvz0p7qrLbzMFhqIJahgCGxIfEEGUp8ve9lh+hmA0ouvfZmYqxb61o0wrG5ze1Dai4cHX
J3EHpERZ6ND/ghfHu7o9ov38FMd1QlgZdo3Sraa6VnvU5NL5QKSG9+l0LiUuHLaAcJJ1aQX/JQR9
1B6OAxOWzfM0HfSC5cBfaiZivtORM8BSON8+SOItWoOVkAXNL7Rd6Srj6zLUuyGBGV5HYRwgDzUS
X6cvHFC16C0N6sSEf9Dzo4msri12vmlJGeR2dZA2jdez9MRtoFtm0jhMX1EpOXqmh6CnzYi4dMwC
Mbr3ddv8WEMc01GMisJ2dEcZ02b7Pqtt3J8qTB2m3RyXhavkG2zLsOrPyx20szePnu6E8Jn3QGPN
0ZlXyZmhRvf8HFsycyVBuMrnTDCQT5YQJaF5muJiisBAhX5onNsmuE25SEET0v9gs31GEJEl2btK
qR/bI/98HX1HS5M0vduUuKjvD0FbeCwjN+3SjVFujqSyD2SoUB4lTqKV9k2svr71sWt8rNiINDNk
xjLB3ReD1PcIhdDpo92hMboDa/qrUKPLIi/5ZjRaG1cvNFcmxXzn3JQDPa+NQ9WVlTPQ3DMLUL87
SvaCHzgiuBEbErR0t0DbZvaQ5ZfdlSs2KkomCrArTdHUBxIlmhq3/bQqUvFrfPgc/rzx99nLLOJf
Hpi9YKXjuiDUu3hMdIXVbmoHjeek1T5uRBN6kMoS3DiMs1bd4TDcBu1E9waH0CeoYDgMcMSa0pQD
PlDxU+CPWKnu2XwzBQ5ZvT75ptZlAAq93vTs/bg+HSklqChyOjLErZA3O/Tw5oyoMuCH1ClnDzY8
A6spa8cz0wV+fs/fjVleSfGJw+v3tMAfeo66J7f3FyE/DEvfJKIvYZy2B5uNG2KlrDRcXz7FTlNA
pn1vh5lYw86p1yOKg+sBYlGeMOAZuIANIvBxvPggf7p1gfsiqJ3s9b0mrrVFtyhDr63NW55Wbgxf
bAoZ5CdHdGAYdiEAl23FDUbqw5QHQLl9Mee/hXXdy9kP6KoPrvxKmarLSMVoQ9dl0rGW8I6NmsdC
60PaofThEMP/euSSFLqSVuBGEZxRjTSUMttTyKnQF80dNUdi0M1zIpV9HZgzog/IXnibhkThMSEc
3cDXwSnAfu582tiX9UaBlnc91fHCRRcU5IC3fS6Xk+OwdmDuZlhR1Jjs1c8tqPULRDx9x27GtxXh
ZYt48be7+FWxctNcJLNJGCyl8ftKEcXeRn1AHJb4MAjwLXC8uAnFY9TW90dULvytLO0nWSCmRI9w
3fBRX/PyLws66/7ClDiVnIE1q9ifN0dhKmBHHLYPFZ9v00UnBvwfUoWGTkgL67cOaA8i0RyH9zF/
3ZwnxGutCyA8irXUvIM7+iVrUT+jzwJjpri30/ZjEk7rDDN1OG3UfTo9BpFzH6oZ7rDW4l4IfMRf
MQA2MZIMcH1Lm6eGOVoP6VrTOOj1XY1n57QAHYLzCZH6Fk+qkQiKLfBpjhChGUs9LFWSEAr7nf13
3U0HPjo0lNjCtW3ivocfmVtei3n6ZvjF0yRRqchwUtNqudT79uZSjq9BUyy/vzOQbEMHxQ3SsmSR
/upucHyGJJAhyH55NQDQk7IgEUAJhKe3R5x6o/GAPbRjXRX4UU4RDmptpkDnfOxftYjMMsliTAkZ
NTc14sDXlx9XttNjnFT20YGPBRfAazMRGV7aS2nCk3oqKkVYRZZ0pCJwBwhuRNBk1tehU6A8mtpw
pFajhFBjR2CiuCZM/ju8i+gp1qpN28yuGJAKPQNk02JTMYAgY6WCQXVyUC2Wb0JVh9bfX/YnBreW
plspi8dCQd77bYHTKflJuC9/bTGLiwbQrCH6Moug7fUHpq5hxbrgKceFkFZrL10DOEcxZCRpukAl
v7Qip4spFq0qsoOrWiZJkLlg52uVegv3+9sTmiL5vRMCoexIqJb47RqAt601lmuZlPzU9tT9Zbje
3mXXkK4sdUAPiTNLUwjZ3Yl11FvAhAh13Vczzu/U6hNGtmwpvsa/gPB20w/guMauA/0m+nKPPAdT
2V6u5IwEKG7/JMrcub1grUpAEdgPu0AJLyCy4gSgp9OHO54jPhEpIxKI1p2+x3MzMCGPfzCAUHwK
/cz18xLpRJXfTq8La4jGcTC4ElzNnGnkNZpy/o9IbijEaQEwMc/87NUj5hWwcGWscy1nlkQo5jOK
5DGWifST8sDLtA5CwO0J/GaOsik9hnAoabsvmz7nd7PGC5AtVRA7uEdea6H/X+oficWgHt2pXYBi
jppvgyDLwVYMNV4oJWeK0aK6HpKfINZ2k/jpVhopddm6YQUJFF/gqRHa02lCKKOyWVgfROsZ9dGF
1WNA1NMamvxSM3WPgdiXIWrtju1S5n9JsfwCAeTPROvaer4UqXVTgdT0trOvvqSS4pNvAogufSYl
k28/d+VFTbEv7BjgJxTQRRQuoTetKv0Y7QeatRruP6TFili/ctTecPooSM9VgsTRCKhfdvRuLBA2
cPdAAw4U5REzJ6GgO/LQECYVycRQBS+ieDD5P6v6kF8/YAhAPkNqigFeI8uiG5pIs/jil0FQg28P
g+gDIVMDBIn4eOaC8+jEMV4DXER1YyN7Bfhm3VVTpElpOW/TptIc6MDlq7mAuLLZWmZoGmARLt67
28zbResh63pqSNH7RPOC7TJjk39TVU9/BfUMfDwH7YvzW1TM+pzpK3M3BeVMkFMwcF0KNePF1xFQ
ifvgsx6alDp0oWoY/p/hPKHNnGZeHCyFNM0xMMJ6g78sF9cYaaqmplp8mO7GHJ6jVMg24PuEDpju
1xE8vSph8xRh9TrM94S61yYYL5Z5i3GLK646G67AwSKfdYSIx2ORH4+cx8aHc2B8dbMB06tw/T0r
NiMhkx5kpbFFM8gPzE0mhbi+WvLKZ3ZitpYKZk76BCha2b4qJK2NK3SaJoVZ2z4zWEsQHDvu7agM
8Ps+odvK7fJhhIwMcHslaPawKs+/9uFB3FUsio8aj4ABn8iF66/AVs+yV9kp7H8Cb+Pf0yrn7q7h
anuVyXv6mJnvjlGFfMK084vl3djaIWmNfwvczccjBsTMHts6jI/d3Jud+JrXz9w1x923IIvC5oc0
vZZWg0fsM8VFO7WmlG7RoInnK1UgM4gCkfkk6VBQSjzKG8+NeJVZLYx4Qkk99CUB/33SdEIZtrHG
2TGA01VuSe73/zImBh1KY3hfVbIhAKDi9DxtZpUYXPSSW0S0IE7xIOrQ/Xbni9/9oFW0hplG9+fO
jZQG1A9RCevbZ6Og0pqEEDydgyOaP7SyTwHs3/lqeUyhx4HiunegGYwu8iZwTpAHzgWOVtgi0ZM3
gInZXpM17fUowk6S8pA0naBbKi2IR7gROQOnjcg2LUC8iPRpfRmKkgHRAZz9UujecJgh4Gn2jdef
LM+grq6k59VfTzR2UIjq4b7PEigFdWk7/y8rR59YKNuCsp8Xx/4Vhirz1dM/AAp7GGRFjyhXq1fR
wA2vEZ4mpnGEQ8GHaBPG+gOhvj+xsgVYu0ct/izLogc9tnrssIxbcvy61g4zFL6ftG3L+zFhwK3y
kY5Pi5M1qoxFSf//3fQSfdjEfZMsg1lm8IzBbaVIuURtM6zMcj4ocAq0sPXeChuEqozfQEMnYjIy
k/LosxkuJmWsDdbAWwBglujG/C/7ELF5M7w9ToIUW/bAVrNGaiMKlpyPcg6fz2zcdsdgBmbOOYYS
1SyuIOJgr7jowu1MM3FqZOvNw/cQKCLW5+j6/sXsH3jmbNLFBS1CIcn76hU+dZsQ+poNDmNBsnXE
0XXmBsXJwUVfKO9nq023Y48D0Ve8u4lsu7cufhFYU25YFZBfyCKb9MM5Av/B0F5+gYHWdJmDYGw4
KaPjS78+GX72MifRYsjoBEsvYVqSTv0rI8RYw27HUT6r2KyC9SWZcIJl9qidc2mWOrYTezEI+Mh+
qTyzr16ARE+NHvs5f5YeWZqArEazcu59Qi6nhbK3O/Qq4GAu2jQXpU2vyuniYYCufc0xfslz7uhq
wuR9wChuUUr+0/t5S46brT72dWkhhdrmAlxNrP4Xn/84nrwb1039WV5d4CbIP3dtGm1w7Rhvkjqm
chru8Cq+0du/wdpdnrlgh3ho9o9107+B5t9eD8fT9KI2w8SsOAGsAJHF+Sv0ssdPwlgKbgw8h673
OMZoM/+v4VAVp1nhRTVpLd2zFCzG7eRwXVl/Gsvkc7mUHSGtDcJunNgGNXhYOVcxjU+jlSjjQI5d
NJjp8EsQ/+kq+TI5XpKqedZR1gZL9IrTM3wja/ASVndBi09SpnsKmZSWheklmdenLSFEaXY61f/s
wztMhPtcDdI/tod8J0tebJPvYdBTMEDJrMmpzr5o5ez9HZRo8h//RO5a2LVb7A1RBfLKQyY4fVMz
CSuMtGel5CoML2AfKa6Cg4GabDhFcsag6XyShotfdz1iVj5af2fUkG0D9sQdKyZ1KLwVD1X6of6/
W0RGbfuLA6PK5m/toZjea7gPJcm5UkZ2hfvNoMxiXdCKNpG9bH/lPoIw/HtAtZa+fCWUX4HJzJ+M
M/8zqHMD0cejy36SaYcAoYrrZN2nVG1gU+OKpLb8kSZQLbeK3QRX8P/0eO5ZAcmAqcYyIA33/m9c
uxGumd53ViypyMGGeWejoDvGB8B2epA6dGdLP0Q/I5I1aZS3K6i3TRnomrrdSZ7xxeXZ5ylqflzx
G/wOmEQ5lrsMkaVaHiZWfVrjiCD1681NkTJhWJRx4x/wsSmXg/9JWMBkTi/99gBJgZdl+A/LHOxh
vUF8ZlLMB0RqeQIRwRm+sEEFyUhoabMWKZxYgq0kZ0LuddSiK8VJfGSpQm6kN8YGOHxxIyE2mask
aStvLdOT27yxhHnPrxuNvajUAXJ+kstMhCrVQEDHimDxRcHo+l648Sd2CmUF9gya19+AsbNvh0Yn
ahcM9n4g6940kfufXmUZ1D6dHXWJW/YP22oSWtYmnDJhYE8+ay5vFQfQfGaw7Vtrn7QUh/fGv7ea
c9VpmijJERNodvlErBADEITIEokdl/RZElc941FkknPOgNlX0iyG5EBRvpdM4MiTbxcXV38HKigM
2TOAee0rg4MlBvjl+1WpVFe/WMQqUz0FR3+N0O/ElEdwdGrJlqy/kMsDiUYcQ/y2mmdSfELohZ8V
1+BGAZN56Bh/tqTHpLsiw0nR8jhLN+N3fcC3dwQA25u9Os0Fm2HswwgPxaxhRDjzsX1kmyE8XW4R
Aesm1i7E20K1tiXaygxOJYEGn5/kMkf1CYfH8rDuMHB5Hy3rMa/bGKkR4zOWmfg8U/TVubLkMDVC
DieKlpgrxf7GNsADiFm8l1pN0yTTCbeNta3KPUOPbs6lTJCaFUUpg0hX+OeLkQ+GFfyIB0CMfEK6
yszi6b4m9KOOELTmVKfie9FX6Re05RLCIsRSQ+JIsde6ma3CziQU7LwbwBUci/gTlxt/3Qu/g3tp
pA5losPkPuOTL910O4UXX/Lhqvbe8ualBXFp6gUI/QYA30Ik4Txm1Nuo7ZP31DZ4gm5CUNf9xdbw
VyMf2JyKsyV4+CDIBZ1tDXHa7aUsKhiFNwYxHUxQ1U+CajiVLgPHWGCcimr4tgmbSwXxMMeZB3j4
f5pKgvflpPDqKiGfgUaRDRgY4GudUHkyTqa+Vh0fn+Swo8CI+sMR4OrUYhEIx2F/edmZb5iustdW
I56BsMsjCDEqz5TmzFc1Yu4usbp3BT7WEZaD37rA7EEEGQt4R+N7D6wTpO0SQ438czwngQxAsvJ0
ki6IOgZU5LgUuOKe1EgJ8NqV4P0Pi3jXOREzbXbwr06bPy1i1vi8e/h2kVitn5BBmXj59VuDEIrw
YxtZ9yCwb2JavfRmbUm5CJcRvThFbhdR0wKPa0NbC4gJsoSfS/LKbECCxPs2pfLJpPLvc1stlnRi
AdoAn8X3YYpvcLA5nvyEDFAsPlgW1vbtvpFPdO4kqXYr4PsrLwLBLmOkyXP3Z2dWMQ69GEmzr9nr
3B6U6cX9d11jV2890+KxNbEfFYyuoifX8RLeGi4aoQpeOI5t4RBUb94EvTMA8WK1afhY/5QHBBFu
s/1K3rBXegeEFDSTALxHsuFKx24MXRzqc+A7A5ZtY8IlPygH/F2mdRVTfmQ4RQzHQrH4tKc9HfjZ
UBg7mCnCYEUcu3UVxMObeVULoDNCzm2aXC4XQRNswsPHfMySOfbjaRmiaCbrGhoPb/s2x7B8bbOr
FvEoP9XSnodHJ3JDFPIdL44nNRv2wHOfB/CCyqu+m0VQFjOSUsj35sn2sTVAvbtGfctA6JXDyyKR
dWXbJLfn5d/WAzFAoeD5iVYkvq6xRm6USuJaga6YpW8REQqdIaVM+8Ogi1Eo8xey4Gf7ggFZr6qo
PW/8Y+IOqaOdFF3bZAjE+29CVRPptfFfvCRFgwh2vaGVF+JLLCPrA0GYgn8CUFwJgBg7VEfL5hO2
EZIZypsZdoWHuWYqy+8M4BtjgNFVkB4BuYIu2Cqa0PPAqYsgwbsRxpCiAMGZZn5DvSyg0eSZ2uGX
tDglIGxI/V8oYWJPjMlGljKJNztM11fPrf3JHdL8v1OouFwwYBv5qdKED0N9W+hhKaSZ48UHiyr5
OIH/jOE9WssncZHmbN38/VnsWtj0krlXvnkdIMALjDznayhzybz20W5p5eaYv2bIVYBJoPaQpAzI
YcpBuFmd0f6/BWwetCHbleRkuf240xKkReAxViTf86G2HplR3aAdI040zBHU3X5Wey47fmEM+FAy
8tRGECDjJCSXrXkG7zfjEMsisvUQ477lRX8D/Jmq6wPgrtlcQ2JFOtq9d8iGDUCzTHaRTx1FreFH
4jz55aFKyZ8uX6dbeuMpZNizEL0a6l86YenH/2mfK0HeewRsDMHrUwXeiFf7P6LEzsJT7usjThpB
U+wMp5xOyVde7RGAn1jpw8XFrFhi4jBQskwHXvLSlDKqg+61+iS7bFuQvu2b5uZEnniKqAvbPsjE
sMn2c6YhatAApxbgt/QulFIB5Kvf6lO1sFpulmyOwTVTOn2CMK0HC8zjzRuEir3vz0RlUMOZbHk+
4PjtpYundCiRtflW3UEInf6NF+mwhYMtFfxWhhOj3GUXLUJ1BejrG17KDtsqStvMWQtwUR3Mm974
5ThmxNsEjMFAt/cex/Sx1fxPH6rwcRxwdp3qlakFE1i2ESCZ3sy+nfdBa6h7lKbw0iydTVraPIW3
INVRaIFbV71SE1eB7WE9zV8H80cVvUdyeH4I0IPEiPy7G6bb7m1Es0qzWMdPPucD+XYeTaCrDoj4
hlWPlOvB44x+i43w3Aber8bZJdw0QJk/0f/Nb3t/h3D2CauAOLDLri+IAkpGtRo+DgiGzcq+Ylme
EfPAPxBXZqdatahe4e+N8PxQ9DLR5gCnKa9kTBP4xxWVVTgeYojvOHcsyoS0ZK39SHxcLPoJCfxb
CTetQ0IisL2Ll9Nj+B2k+Clrd/1ktyinUJW1ob061aJoCd2TB+N+/4NZpPW/ZbG//SAgXj6J36Dq
0e/JOV3ao9tXCx98Fyfv0aCkospG1rv8NuM14M1QmgnUmCu8vvm6qlRquUOVcnehOtVJhXji7ScO
1UADGEfLGmsheza9rYDNWNKaxCeTx+I5GD1UepB5EwH4XUFfu9653d9goE7UGHdrtaRvwmxy1BYd
GzpJb3ndOI502zBPhRhely2QZlkgpvZikzHuoEm/nQyqsTnqZy6EjhAx7BtEV5voUtlnF4g9Rzfl
L+38gskJGRacLOvLDjot+laY/moglUUMCY3k7qoQ8J5ip6w7b7/oPPXbtCXaQAEFvppDps72KdCt
VUiem6MNCO0VYd5svV4Z1o4V6mStvkLuXQnHNriWVwoRrTF+RqNIemqGbyieSe8th2NHdUGBre7E
gLBzu3yYqukHw6jAYFR3BCPGsAhY0Z313cuSSwB0lIL/l0M73NZj26p2UOfLxMtls4kpxCbZ2csQ
IIjEeKY+wwVJnNsJzF1jaNM61jt+c3tomOAej5IuutQmQgoRuSl6TT1k3NQluOfJMbGYd31YV9DK
1NYQCVdscz5oRfaz18rEqS9MxDE3KhrjRdr4NRpn90rHF4u+BmcBg/gr9wxvJv+WXN7nD458qteB
dMzcFcbz27fIoeP3O4tNojWm/TWPvRbjgxAbbcBRyiqBI2PMdOOfGQvvoD/2lujeFKTVgd89GCcx
OvZ+QqXyNrqeX8hrehZpUCy1DNgXDV9hz1IoOEv7y1qqAfJQ+0kg2ma3aVV0VdMFQMdKfATzfJlR
JjYfbHKft3BCyb9o+HJS9Lf5ALwUdH5OJwFFD/dLLnowKvflENHw5SgIbd5sX/NcqnIYDsJ+yJBw
L9g0bGFCKPjuycEIjkBc0QC1awHWFeyc5hFsViIGrZbncTVT3z+/KJO5Smz7uSjWGdjW7P+fjy7B
AWgi6RiyEZTgFhpQDrv4xpT1Z1AUIny4j/foJU89cJcq+LHYhnUTUTFSBzNRdhuFxVdQG6Q5Al3H
X3zOWld+0pf7dW78/FVvza2ePddtXrDddjJjp2+ZfCZxFEYMFD6te6/pUT+WtwrMfQpx0UOV97sD
kTm4jBnEA0zfdBWiSBsVBdbjAJWfyaUYvZg9r+zqlQAoL0Ie09KnfQqxY1GcUwAD0cqmw/ylCQTp
g5zurb284ecp0IjWEH/eo5Gy8FY2WaFldb4vfKegyKa0SZjdVstgjBw0+psWKQxggXtazZGz9366
sr0c+WuRbywq0RD6396IHwPH8ffsQe+VXBJNe1IEjLKLNzqwYnzItqHOSkAU7J2336dH7OQnRkF4
cKUgE5zJhr+z2iCd+k/Jv0AQ05w3XrxMpdvFtN1L9ijZpwxYDOA/2Z2syfuDZ1v/EbXFGsZ5oyQh
JWpu1sol7FWP8EQ1VAj82PpAZJ/cuHZTXPOedbx8kggb5cSXbqu5sRkmH6rYLY2CL+VC63e79qXz
SXLsHcwPTr9hBSagGpCvAGJwwS7D3NpUFXlplMUOMSwomPIC7mdfD2xTc27T++NOFtW9046nTYbj
LvA3NywQyPVRjWYF6xeMDQXu4V+h1kosbUOgGPRq4S5u7Vo3P4r3sxjugIKIEtC6rAicCkfPtbGg
Gi7opqn1XwVXbS84KhskVpitVu3gxkJ2YiCLxltPgpQxq8b+dVCd6hTZE/bDjIkcaH/igyMgz/oE
Dy2EzWmy23XEpXWWTGzfHi1+73EEhcLCmqeweHDJLOqUijijt+cutDaak9be5rqmNe7fJ3XyrppM
lXhW6vjvxheMBCL9pOiJ234A/TkK1XoxLHkVr7iLMw5JAlxgfvrivXkExAGucyCT7jxXUdRiXHT9
gDXrgh9RWRyqkNehYZi00tANn3pfpNb/SJ+KDW/DPZtXawKrkYPPOPA137BDxVvDKa1Zmj//5cLT
iBG6Cfh/LdZsFwBNHgIqTkj1WMVQT8xZBWo++I+eo+GhDeqx5ugdrYnSslHBvZgn0vM4bIqKghYq
mxkIzPhZPPVOtkBHgB1S9nPA3a834mRqas5OnMNyucSeutHRMPMDNSt7/o9KHwWjpMjavVwW94wl
i+Jh16ahO7jFjV7eQc7Wlp82PvoqbXXbXiJ1k90ZN1Vf26VVtkHFBTz9T9uNSNe0Ix/28LbRjnjT
kv/Qqk4sMjtKwe8fvS0QN5iwy30nN9hSKRlTcaad8pulQ9qfs7mFUNHG1q90o4L5nqpt1qk08LCZ
qLYPIJh4gyRpuysXD6DxN317mjeRBxEfS9dWStRtGltANj9eICZYcf5eSRFLY6S+SYEnDITSaiad
vfDwsLDguuVgt30vxTuRWnlHG9zxSMOMW+doqny9q4xsk1bIQaX77oN4HVuCb5Zar/A84q4yXk8p
pHNzX7tYT/ff1Prc1/NS4mScfUpo2v/Ysqlx1OkZT0vZ6RFT68YlmR/1cOZJxwJom+leYVKEo+Lu
l/Ng9P29DWB/t0YQEgUmDzVhV+jGLFPZvKGSw7m624lGJI+BBX/m6PrBApaRw9esyWrCmJ0zah98
uEhZiCcZ0DJ0ltVHGhVftFo/zdisNxeuteVXgW99DdA+S/WRXdHEs4LD/gAmg4wxpAPGkPtehcdl
Q/am+Rnnb8VKIdHHTK6gO1F295W7LRZjJ//p/qDJRcWvhMfQhbaYh6hdUOI7RPe4Yf+3XiUa++/W
2JqIWAVBvpNU97BsKN99Fh56jVOEV/axPeUBBEmDqHVSeIc+qu/moPaJOFZI9F7ipYHH6cfRmm6/
KLiXUVByiS+PNwAF4Zv+6B1cndVNUMSZalP41qnDroFEF6hcOcVH5BmNUj2ruawKaCLwsjj2kpDk
ppM8OitAD3cmRdP08u+/SFurhLr7t0AlJFwtd+rpqlHDr3Lzw/ofjrYBxyiZkRyhtAWqUGiodPu9
qbj9mX/SVKuWdrcnEAtaGB61EUcVrHLy+MUXIj+dS1MAqlO960+0/G1ClySdiva8O1OWXk5wQrgN
3ykyo6HSbHuVk6l+6C7o7aiiU+DEulDufEshSKYJmiTwLraIXQaL4adIPbO4OMZFs0MQTBGAYTfr
XMvdq5Xlj6MxK7pSraQYSYpb0ZuNRDt1pnhUoO8q7m7fn4KHhvm2fZnI3YVfcp2q4Nck4+s9xOAK
RWR8GH4W2xqLvSBb0k1odCrIjv4W7ZvvM2qK4+FXwctdt/dD3yKRQkb9xtDHAge+3gBSdU5BnVRb
5cHLRvjH6Zx6bXSS+mJDgw4PROxHIDC7i2nDtGdrzfajRObzpbK1zuhC3oK8TYJyFaGBe/Cbgnvc
AIfLQ+c+Izt2SRign4NvfQj619/XZDM4clJJsqQZaARqswLSA9euF5R6vSgqJb2p2gM1DazcRMfz
SMHpu7qmWtCVGjUkMYwKPWC8OfO0BZpS0L04gug2Kcu2gAQFMgyutVQ1qEj6G8YXNk9GRa4sQGfa
PFZ2WE+T6L7VeLkRNcEl2umRGBc/kI1YKlUk8wzt9MvQ+f+i0jfRyEUXWGeOgOZAwJkK+SWDRcGF
UJPrl6+BpJQEhPNOx1ZVwZj0P9s2/6f+OcAntLgDasHvrgUT3/yAVxAiAJoMfgK8b/kwyDnuV7kh
arl8kX77jj6CrR+NE0qanevnu1jQha3j9p+2Jafux8uv+6Zbnun8jPm38ssHCaht5ztX8rVub2ZY
cH86XcR5JtFHWXXI6hb9MSQrwgRXuanmg6rjLr8DUuhmVuUygiuqbTUbgrVztGPemQd0aN+DeJNu
YJ5shO+SqGV/eNXmY3U/IW9yHRzNqSM28oCJB7dXEwhWHfCj6Eu1axKt9mdSaSuoigoro4mMrIe9
wJjPde5YBW3UYeDEJSk2gB1oqkkW0qjsbUgkBOyIpRD8Ox6H5THDE21vC6Tww9ozdqVs/ws7qAJw
5QJiAinAfqgwe2SpObNtAWvfByVbI9Ki90E6NLNDttG14CzXMbGi0Bm0Sg/pJ5qXvyGmU7MC341C
ZTFZi9qyUh6xDbfw3Fvyu/MeannJ3tLTZebZ3kumzflZR1zZmrJlWZQbWoH54apMd/FOlllkBuUv
zPlw8P6z/3F77vSG91ooRSd09cKCNfTDOGMRQ+15dHJ5kBv842fWcMRkUWegqVFrxrVZwK7lygOE
LYRKPgDkiuQpdoKo5h7Ks06L6k802h4r6veV5+TtPaUjF63f+1VMrAxj8fCUFaoC91CX8U2hztjr
lY5KUaR4H7/dU3HW4vV8G/tGihug7xnRduKnCGD0wEysvKJel6QpLD9uTz+OgBlG75DqdDK4gh8r
whPAe714oeBr+SvrBHI3Mp8hFDwFk1Wr4s4NLKQlMrxp8mcGb77gy3fobn42KObSoXAKPHPsaKLB
uiBAW+otrMJZFSDF2/a94fBrfCUaBzQG2fkW3hNaHN6ZpFzSCInBOa0FTCuW1XNu18qzzYiyUSrz
tYQKpNeFK8f89drFDzdRPXPw4Mm0zZ+nQgiAFXLZlemUYHjbkXiSKpLXCuwjNdYUjqDc26ngPKPK
NUdOt2a+oRhmWu0xbpWeZGnkOVp9gHXfpJvcDvDnfHN0hiFX8ce+UN9H485Gix5DGXD0ulfodfrK
JSwHqGSOeH8LndaLXWHXEpCSbP2kTF/tB45M86kpqoLvPh/32MXF0/SQlkNlkZIKYXp5Cze8caOZ
3ufrBByQsN2AkPEDo7ID8hgTkA2oHcspIwM/kvXtH+imDyo0J0ndMtlyuppms2X0YMLM3kk2LLkp
Gg4czkAKOTcXe9tAmm+YjT/Bf3LZtWro1/4C/A8Gh46DiiSVrVURYokdQVvFr05DFaDEsiqkmzY6
b9ppWv2Zlr6nhO4zfp/vVBhT57yxlsI1xQJMqCVZ0qO6NWp4TDyZOkGxoCJ/ZWHUz/vz6gTdnFD8
M6uNc/n6k/NjlMNg5M7Mxc875IqByh38Q+tSyvIzrv9wKAvOn21xfVy/Yc2RCPSrmyT5oU9tsJLz
s0tFcC7uvgNatYnQ7cGYTw/uPZFmgMbXzUJ1kOxKE/0zGYqgn0a/S8MOIzQ4WViARnnawGVddgYF
ND4uMWysFmvNw+S3L1H5+CY2V4hURsDAWt1sbA4+v4NRpLhYZnuEv5pEhpAkxK68mSPseCcGwIBh
QeM0j9HPbA9dQ7dWP0LuLkd69D8X40zL018zQTezI+o/JZ9otiAIkv22bKh1q0ygaGbAQR3bZS2y
BUl4s6DUOrLwc+LGcS+YnSAm6mzA+7XGDHArjcS9IXCYOaNnaKTwCOlPx361cgigrPGdqeYzG/lj
Mjp5JyGImraq39vCktA6NP5VbHpanBR9QaX0L+RmQz0Q0+Wp5XJOk9P3Q/TzfPx/qM6x8jcs+U+w
8T6VlcCI31lep6nIGdVxZxb0uLoe4A/M45Hcb+hfvSgNZAQVx6KTniHN+USZNf4AexpGmw9e3MA5
96j0ds/CYaJZ3XDraQiFpxG7wpmyc1tFx0dJd59U4BxAIeWk4xDVphUMmeprPM3qtWSST3Szrwj2
GgDcxo5BKAhhxvfa2VuA+TWNUCD/fMZB8zC9lWCH4LGsqV+wXxgvnKsNHa2xp9JyiUfLmerqoMVR
AldOWIPtxswqK2Td16zVasq3fa92qa5wquvht6LrDamoVUQMRx/OY6ZXy3TcbIjNnXrmYRR/wVy7
rGt7ZArFy++/34Doujjv2DVbABz8kGhx3IjFKJEyvNdxPOb4O7+jehTeoFuaHenz2b+OmqKHncFw
CJw0Rnya0wX9gQj2GAq0907hB01T1p6W3v1kmg8GrMWZY5RhVWjSJsplFMgmgFnkH/BhYbf4ewE9
RZXL4jq+Ij69yA0ZkSNWns7bHnY482qjQ3iQWRD/I75eT0jZ5tMOBR/uoqh4RQR9WrhUqAPeU7Ac
OKOlK4CXrdUhkQGbymxC+mqA8hxsSEK3oLaxjCeyB9geX1dqD9maBDmDdF6JVW3I8DsgGNGnYpXF
4c9bDRuz5gQhQab7mwtSq72e4XfhULL1agvzlkfYkgZP+cvwQ/ecljgxwtrdIYwLApYuWyLeFrxd
hVap6vtQ+cAZeNd7K2Apd3e9PbOhCyeCUWeVtvxbstBE5bj5Ts9PpyraFHNkYC4heto3Qdehfa1k
TAlOXt8/phQGbqNbfTTZyMfGsoiA9u9axIFxrxkaZrOa8F1+1QF+0pARntHIJpDwMRkK4A3D1uI8
xUOqi/HDbdbQLUhkSzZ9Nh0YP1AsRWjpgVVVRFtM8iYXcv5Fb+LuBQNAb+qpguZDf1p5qDsQWV1K
Zk4/kXnj9ho8iTXoqTMegh4WayTYDS2xbIV48pOs4NAHKeORaF1HoiuWqk5ehdUuLMZNa67AAMSk
bY44D//TiReD58AyNXyCW+AiJkYP2+b2fh4Bh8ZBKyBQ/dou1sZDkzwVGpSQORMTRl/s8hqHF5tA
VX/4Vu/WKrTIOwyMBjh4n4/AvFFYTuQ714AfjE56rsmbTqpSfFAIzm6kMqHAhfUMcuRsWmwCPnlO
x2drvquUhuj4bqdIWAVMPr/wR5N+wNuFLP6d8jev6Cj09YUGfDUktbL9X0kYBrhu9Tg4z0B2jqJu
WiiICarY61r7kqEntkLKuYPU65QfytWW+abS2HP3didKlcW4T9jEp6315H5+JEHs8toAAOKVePXT
H/1Xt6VOI/SwOjHJuUHaW0yttPXV+lT47I6yJrvTYZ3+395N2T2kE1JzYEt3KC7vyMMwXmqjQrcx
T7UgOC7meVY50ITdRabDgR9H1b084UnwAesi9tRFPgU3GDZk6Nx5hdn2WrugYAAR2BPEI8mVGgyu
wm8lTYb+AtfeQF932r/gySONr+MCE+PC/gJO3mgCSH69cLBB471+GMPqvyjTF7bzF75x6oP0caZC
76kNMmz7a1e4Lme5QzzlEhRpSBCkEFga5RF6HuiF6baxYuI8B70p/RNwNyOJMrY14dIlXzC/z2Rv
tHNkUQReqMt8e+mi/byUpQGANiYBi555NvtBp6j7E0xH4gN226dWy7+5SHfkc72mNS4m4jDtu6Gb
SFzxHpUW8rz8ShryauBwvdxFHEB3wrV4m4p7q7ON51vU6cqVtMio7CiVpKojQVGf5agUusT2tZYj
2yJTSI9OJ44zP7tCL8485VPwu+7Xh+x7qfcnsSg8+L0D+f/6uSIeCN7VdnhT8ep6ONPIHNuOEdY+
dfpnduyYQJ7SP2vWQp8/dr0cMEstF64vdzG7GT0kR4s112VmED8GKy+99Ye/r0JqhzUVdhyrRaPA
tUzKVRks4YaSpGazvBfh4aIef08yzE8JH8bCtA0TmfeLXFI5KF9mc8ZIwB8pVWk0MsDLVXlTe/aO
TLR1iROgVY2OJVme20OehVYpvB7xm21R7LHoI0WQ7HAnUuPU8OdHJmzdS9/O2aFRYTBw4+u5IVjb
i2AEEWOAZh2xE9dCLtUkEs9+bMNJbKZRIpmCCXU0HhQ8tOjexhpWfh+1PNWjJ1LaKgmKc+ed1yzA
uPflkm62+IHqR4UVDtCrEauanohCdGyyvc9vOXDh9FHzLhlPzlxfmv4t5OP4IRQq1N69BZaMrUmV
QG1l143Pe8M25FfMHfDntgavXbU7UiJbJ/gvNVS8nywpj//u3twcZsOhH9BrOIJQ2DEdQEZqX+Up
qXtqdFaBmhvdibpHJ7mT9WetudkORo37L4EG3Xxcovue89KANM5z0SCTC22X2ZQd3pffAfc9wa1D
kNHfinTll7ZOykl6OsiC2bOHaZpD/M1CqOI1lKEdJPLBrHW/D4PFM5zQIJKAwZqoywL1aidnJgrT
t80nXwNDCF/TdJ+TiiBg6sL9swuihtUCMvUCxB28blVOh6zYqVnSt2oIBJetO78bP/W+z/TPGdEd
JXA/pcUOd8JrF5/m/WDPdNuyp2jyG9R2z/pqTgSRNwtqTXBluc2kKqwWnRDHfLNOW6QcH5M8kXbq
60pMB48q+dJLpN0Cj0g/JHkzecUPew53+U7IGF2Z02Px/EKew0c0J64Cqj2YFaU/JTU/O44AHcFU
CGn/29wMZ0LWsGd+kT8By+ay5pm9AZc899cVhTdxRGab7iQjBw2beUVX4Z1RRHCgWpCq2AKtUDPc
bDTsFEpKXjU1fFUT8N0T1P5HerJ97Tvx/WCP+GQmCEJF/lFwtekvLCyds96jurOK2zlbj5MURNnE
7YAPcwmNTNyyLirayXoAHIMLMNpDfeBTn7m4pNhjeGseU8GfkkvwyiUa1IfqkJdU+pEeLrm9dov2
gDyDly7ESkrK5+xDC19UPIS84lL6kaO9KKYZjCNRTCLUpzR89E9szYyxQVyp4VK1Ix9w8nssYvPR
GbiRrX47tY3gqzgO/3eErNbyHQU3Z+0h9218vdwuOzmQhI/eT5NhkUf0fJnFYIE0/qB9ctxg5TvY
yU34YRVCDgiE4vcQseggDBYoAP7+WJDAQyRrElh5pzXBHzvAF1boi6+Yi8V+bjdTbYksF5/ncCWl
ClPrIK8wQnP5y1O7uiMaYctvMJEMhCC7uTYd7xipQGo+OtV3gskeim8Dei2dym9jVgE1KKKXJVHf
S3p7rOFhg0XiMjPZowoQuApJV1bWjJRNSvlBSdFBCIyVPFRlJL0PCMARQ0sIIuvwQbYNOSncZm2N
f8Fq1701s5V5i+9dnK/mBgbTH/WNp8fiYxEmB/HegTiQFZzpngY6lXoo74UvPOzEDKy5u24ZzdEb
cEiyyR4OcKUIm1dVn9MvvyiRmhv4XIWGt2JUocgGRDBK++J8TxFTkdCC7Dq2CdsHPFmG2KfZTKpm
DtqbCvfGUZy9zLIJftX6mRBfKeVQbi/GMfGzbBoWkAltOBTFbRgVYk+dVkrLTZ9B+IqSYhr9q7ZM
xOlvImQ/YhL4Wd/Dnn/bOQCwRmQllbdheWdrwiCnLGvBc/xCJZ8WAZzQmCXXYivk1y8wTJUD8wKG
5+yklznyWtq3T8gB2VPJJD6DDYt0HLl9xeyI9BnHgrFffv8cPjgzAs4uzlHfE7pNfzxzCQykuLXa
7bN2nGHr1HFXSeDcx/S7EigibcsIFxZ35hsBDciFAgjevW2VrpaADrHg9qC4V7QME/lzWvf0kp+Q
rFbttqhWbXySDaOU5FHT339/O/y+F3Hs573TNTpoLHg/tT1pbuksbXNQVc9vLBC94QH7sk8bzvZR
MrQGb1G5Ws8JqNit3UuhtdHkHyw3+mnPLhAVEMjXI7sNgIIE1OwZlHLi3+0sWRQ/7BdAfNzW7UKJ
U0CQmSczA0i7cDKJD/pTUqWBHl8JibJs7dBc6ijITKcHhXKi6Q8F4Jx/ta77X42t57Fh6ZcZchmV
XWjQLHgAw69snEyCa/VvSJlXEllp5/huqFBtOmWRrhn+9g1OE1NwylicNUednRzBDUWr/tsk3iB5
xSbts53FWQlGMavepFvSi79skJeWTwve7fV3HV6Ljuu6uQy7q4R0CQdzNb1X3yrAAovvuozFlilv
vgcgTNPX2q3MGNx8ge7srXh1wYTfn/eOBSuyEyyZuSmgbaSL6jbROafF5w8FkjjurURECWkhXhgx
MaFyavdd7NKsy17YZxq3NOdfNLU/ypSX3VDYZ9Wz5kLcrghAsmqaVrBlRtIeaIGQExm4+Z6D8VQg
wG9gfmks4LrlIxWs4fERvu11l0YqXVvhfAiQ0Kj5MccZFYjteMhlw5eYjF9RZGmWjQGZPZF6IVNC
jJCyyFr+Db2piCMxqbMWFLGZauovuUy8TC2r/zRy5qrXV3wfBMJSdFP+NTaXeTPPQAslVhAHyBw3
U8Xl66PrivnMMaNz78tVWltI0V7WKTU4Wu+aaILvLuB+igjzngcHNVs3TvgElSaICtJyT+HcZDFJ
/mHIcGipusSZLZWAjN7mtDqbovfT9qKEMN4XD4akk/IRiJ3rHZOWBAc0vWmeNnSbqIbEM+hOT4bR
p7qMVhE7lpMoq7PBLQyH/drXPz4l3tBlSa1BJdm/Sn69igsS78dHWvWTeMLDSuN9MnfGxQlJSUF9
C4wUhbEs0kPLOLsIUVswL+kDbUoazj55Ldr2/sI16rOhI46xRNkzliwekjtGtQaGndcMZPUVQmjn
8cHdFzvGED4nFKGlMvgXQ7uc8PTI0Mh+u/ypCr/v+6t3DhBntGm5fHV8yE3Zbqnkcd6wsZ33cTHR
XJSKpicSugi2YQZ/PUWdOy/r9GFenHDIel27G+62j17+uWeZYMlaizQMUpfPR6eQXplX8ZY05Z7u
EexaWavAfRCh+mF3YU4xUS9B3n11Ndqb2bYNktkwLWExfttOX1V/ijPGzxCbTr34FipZEoOB6jkt
AMVwwrMIZjD/7VE5owUafyBlKSkqDIEHxYWHnTEiTRv1ylgw3ug+6TzPeyz2LGVmGBaki0AdvC6F
bmrjMSiXY5YE8wR6+3NHL7jo+2EWMcB8LMrgSGoBvdyhGmX/+3ZR7bHu17zKBxf8idzygcM7UlpJ
CFLSvrhD/eMorYFQF4m7UeBEe2v/IRsLvOVJYR2M4jjFGQQH137ALPIFwtlt+PMmH9XKFHSDvwlL
jgVOza6MQYWSvvFkAIzEpXa4SKCApBWFw7Q8m2Ut/gO1+q+cR+EBZtvwf6uzlmM1tMqE/bK2+hEw
l/3Ix5ZuSKMGBov3Hbk5GxHGFDWKOvSR/UwFtzLBRCzZZS/mCb3IktLlD/F7iGzMjNHUu5jWcP4a
VTquEkSvZ5o171cYMW3Mf93E49tDt8Sdy6/kzxZ+nQmPKAmic8CyTU67YeTRa4SQ2NFNK58tOj5U
j3E+vUloO7KRXAb4bztnNRq5e+7eLpfGPnsRww7yHrdzO4eiyzGXu8HaUqtCaTy0zeSPP6bf6hMF
VPSVkrEF98u6SIjiH1pKs/2AXWtCnQdJtMFhvHYsPbSsjVdys8k54FvXGBAuPnROiI/yklqdV4A9
mHZG4TvfmfCePDENBdWbBzwP0RlTLsuYDI+cIXtA4ZUTGnu5nIAihg3MJTcrVIiSdK7JXkFOUmk2
TE5F9IHYWmGG87FMxC1wvzvM4reECWZNCCkqIgfrDvbvHz6MqCoRBo3La0xbelHwZFskNowBm4Bv
YWSUO8LwygN/wZSlB390qX8Htk7srevGf08GUP9CbAR+YVNBR0pA3Dxpd1ixdHZDV1r8F88FPYuS
OwnLd/U+sL30bbjbP7viLNbYjCpn5Pkv+k6Jy5ibwgsnOHr/D9hK0Yzt5RBmxM8SQq+2Fe5mCXYL
8ZiZuxtsCftN1ZGHCXstFeVaxULcwlmPPY2phSDQt+2Q8CiBoadRSs0d1TLJdAsolL9k3LkR7E4s
BBNbhTjiky0GxwZHD3hdB4VwdI8zcXCknYD+BToxKmehjqcJHoiHcrHMXNG5nrYZf/6cw203OjEQ
Vij9KQxn9CASmtrrZTh4rutjGn0+341pOWU3LMJ+la0HXqzgqCHhqEm5xDKxPUj/kHIwRjGEIuq1
9qDN+0ESnmqMYJh8HlLiPLJyvcMiiJV8xS3lPuRxBtlIQAemI3ELltrzGARxwim2B8m0NLf184EQ
UlYTB9Yc77IE8F2JmMOXQli5yzp4CM+A7gR9JxRkXEBRQkXGXLwIFOdh52ha42r0Qulxu2qFYZQJ
RsKBLzaxuX5Q96k9GBBsYDtjZxiQMBOtjExOtCatn5/yYfizdwDNiZTHyFPJ1OAfJ2UWcUPmfiXT
/d3Z/biH9OY8BUJzxDtpZYi2c71dd1glyqgKUt238gEdw3+lHvMUIlrHVplUI7rr0PpuLox2G2SY
zzvwHUnwOFTfOhjyJJuONsZqDTqLJhY9dC3iA0rU5fHKfM6Z0HAla4B6p890J/b8cuJBDluCi4vR
5dsKoTwYJmqmfX/pKDLu/Ko+1s7HsAa7zqCvaUcSs0We2KN0IRnUFgTKpBRFOomNDOQcEssAALLM
4juAt5ccYKoouS0sS+kxjvmYF5OtU8cfy8FA3q2SUMaUvGlWpHlfpnMX2LdxbhTnPgFxpmZuZzGe
5LN2/o17q+l3zM6NLP+YjHTNUCYIJi8olsJxE6GFUmVmSYDajOVHipbV6Bh6R23wo7I4BHEzIAAr
hDaBrOVENeQdbX6oSAQKyiMYX79JMafEEhzPgTJwqZ5O4WyDf2fAyz/piNOyyeBF5GpV1KEBsSaY
CUzzSj1E9dTAux6zB7w2c31EqEm8N4jo4wwGBHePyTVRMR4ISWFT+PA0tLy11nGuVR84Ge1e82ZX
NL1bk3KW0SS3oWo1MWXK/iSJEBelNOXoVRvMA4TeaNFRxj7AwahxKKtjaNHv0yJae89XuGohzZOA
B7+uy1jgnVj1KIp4rQV/k9BQ1NpEMxQ8utqJEl1cwBtG3CSvYxTLTVKfBXADoxyzHGqdKm8+Q83Z
WOVA5SCeQMo1CWgUhdppe65o5LQ7E6dDdAatQPRRtIS+0LkCnGdxrWzJaFf9LojgTGb6yrIzkstJ
b0ycYz4GVdw8ryqZY6lTSdDhICjsnHsfsH9Cm7UWNQkiPa4KsWiNZzrntmSxehWiUbFT6D2DRe6d
3YuwkuZyHDMUSuWporjfr9xFynsyLGrYhvRKtDiVidbW34SYrKvhsAwRpg3zLC4np6zDbmCFumIR
Wuz7m6ce34jendHs3YoNj17PcvIO4K5lL2bUTiz6ECwXd8FiBElK5MrXQTf3MsZxnunP1xLcinL1
8RGuZlasVxSCqwce8hf7WGQDB1oy/E24I/AVBYrtSO2JmexKfgYqmO8T7Bax4GFU+3T83p83xeBB
ykyl97BNL6F9sWjGcAxydfmAZwBITslPoUO/EEOmgdllOVqazAHnU/1JqGpCC/1J/m1gIc8Y0/m/
vMlR3HNH9HRSS7uH4yJ2RiQvenKpRz/B4Qdppzh3RTUZgz9+AfS66K8S6Bv+UhZyF1xBG+x4a75m
pFM8Eq3KH4mMNs3qH+X5IJFor/ojwIQnJXob3tNlNrNtwIIqI6+zLItM/8GEsH3tGPS01aojzEHg
pFP5fFLOyvIa1JGXjv1c+emWXahJXOv9jXYPyPOqAEhXfvaC3KKw/izrt/hMqD316EgEjp+trKWB
3M8Cs7XLozHs8VyG1BHiRnZnNKEKUv3whhJdxcGzOv0Pj7g3TVjRELyZn6NUxUxGTQj+p7YDu/be
1AQbcSXlgXqSx89goQhBfjKp974tgamHUnrtDaKYUQ+sp11o1wqm8AAVE1hLk9QOVhhiu6UxgUx6
DLdpwYCcxAsTEmt/Fhc8wjmD9DNFuizH3m12OhpWZa3dWs38xTuHrV5TT2XWqRp/mYrNuKWfqfiP
A6ywUNnndaulsfpnFH2SB3L2TiqnOtuseimmbKeOugffWof3I8Z/hMWT9I3lEUN1mmoIeSknaOf6
Z7jb8fnTs9bjlVzzdHqYeRLpmFGlq7JXrmt6p+PsnYMsGftcvCUM3P/MPKFZLX5xRIHqPA4E2bsu
dk9UW0yWnFbiyf8B5Xiv5++tcINYbdkU0kEIET6QkULp/R5EVO215iXiEYZ3Bg2/RPJNQZ9TT9XB
JRcXHQUh8tbnm4BxF9I2dyj9L8b539vBVrvly4eikMtZYbmRewaNDBnztvTK0wHpiu9a5+1c256A
XnnUAZ3ivSoDuga21Tfpva1K27nyM8yfDmeBpolJzUUw2IXtf91kI7vBWpaiqRat3HS8YEsJiohU
ypefEqhsWWCa8UqWGSM/9G6SGMce25m3TNpvNomYWex+emVDrGvIMbqd0HlRC8mc1hJrpww5/xn2
urwbQxLrfDttjMuoyhimJ9ntEt0xW781dRED8evBrvRvRWEzrUw+YwhlPMQM1SN8+8XDen0Yg9tF
gt5t01OMr9IdRNkUqlztSZ6OUuMq8sEbhT9E/D0mGqnoesfjTENgdS5ez9qCShNglyNk0T9TwfS1
Ebf6qE6YWDwcH3aSMy4uZHeFxIktWeYAVYW1GkIE2VUcqRw2tSyZYNxIcnfyOIzG7y8U3+zxzoeD
CrzXousnXPIuDMl6sbgEsp5OnGtfp5UHbQenBeGcc2QpVcf4CPPenQTR77b1mdlQyHrn+JpBt2CG
RC1FbFxks3Lwz7k58APIr1fBLxBQ6+i8tXt1ULFtVxaLeQWdVTzq55ssSQBWneumoOaXTnxTwDsZ
eVW9iU2ewennPDs3frhi6ROxP/wy0Wkvlra5ADwOWeKmMEWXFDNPAUQWaP/W5BLN7Ea5UnvLDwD8
TduBYI5/3V+MmbsMTsnLLRYSStWQsjCuIVAlXwzqN0/J6s7CgxMIargHwM3fj5UNrunStEx7zZHD
BFoGvVGGpirtpUFKe0z7XfzGg0CO6N5drAVpxghGv5vzEPM8K5zH4mCNCE4wu2vND6A1RLLd82ea
2mGvrw0RUnWM3XcYNRcyetx0uougqZof1G1pPwpUmpOx376+AIL26Jc2jjIZ+L3VILqlITpxi6tg
6pAL1DL9Y7vQ3cmeHmW+y8UrkidmUsi1saaQSKWhu0uCXezgwtV9TAZaPD1qZEl5hhSp/BkI2M+w
3ZfdoWT2H1p/bUoddRi+5hthjX6NhtNrewS3DkvS7fbnnUUR4IbGKQVyU7bkIxWzKx5OXjOGM44j
HTiCXsWKoxXv/D89yRBkVms36N4Tzjm+mUxrq9WVFyH4qEumblU/qIMoJBAUW/Dev+9NCPrAi1hg
8Ek0fsDAZNGfLrTAjvICCrSzZSbeVr/Z3fukiuV32KrzgvyBWrMCaBjhbAQYj/uYYMmDTs8jZ3lh
JBNSZ873xA1/MUa3yN0y+W71hiC8tC81GgphaK+qP2qdv6tnfsikNDp2SACVSVskQNUmBUAz6MyP
RTN/S4J3TaAT6cG3ciIReHcLQaxQfknjfyACIWNmgeR79GhG3mVriIYEmdrSx1QKN4juISResGaX
mjTzB5Qgl35gTi5e6O4dXjl70E5sWWxvu0qc7B6UMLtfQhT8odOHiUNvNLv2EoBnCy7ERxiUJMGe
iFk39n+RaxC5NnzWAQ0C61UWFfP+2ipOnEy1xlKsHt+jT545nST9My/wA1PfT2JUfHOY5EjCkWmO
ks+14xFmxHCcExnfNsw9/OF25Tv2TY9koDlpBYgd1AOb3LQxpgxfc8mFYkSSmXke2nIHB4q+Phph
tDCWpIMdwx6qmrfHgHvjpEgxKW+Td1ItoGLPDdUL9RbJsXOaiBe/Vd740WkgZKTgFkw0FiwNjC9g
2lq1CxCXGnmsTS3KtnAtaQVML7GL/AR5+hrBFywwM6nBOI2CzelQSxSUZ3tHUdliaj/hOX4+vuOD
vfhQ4pEjMrS62NYiwR/58mgVZgL0J/8Dm23SLs6TwEHq3hLNryHkmG+zJYrk6sBzJP7b9lvnniME
nDSX4EagZYH6q6X1O9VxbhG09XjN+gQHLDkaplBMQTSEN2r9FqxzxWELaQvhJM3N8B4vOsyN0sKt
RjyYaoR+3BZUIh9Xf7kq9V59usS7mIops/1c2ap9Dz1/IJRZo5QfKcIjL/fGi5fgSqdaNcqFaPvG
XpakFGitJjaUeW1ie8rSTrG3O0gkxwpg1iXvaBgAQ5nYJqruQQrhKdjHI2Rud6Iwjyr61JfUWtY8
YbL8FxZR+/jySm0YKDbPH3BXMt38vKYTz/gfUP5O7eLgmaOoTzVK/pDyR9i5NquRhpS1CC9xjPEt
jos6nm9JnH84RJ2TPxlq6E1r7sXNNOy6qF+0XGlWv9h/KCw3d31ks/SuugAX+skGDZtWK9lLkF+a
SgG0GvayQxb+ytH91jMAMOzBt8nJevRL/xocDOZF+riAIDyyzamegiacLg6twesTKpnvJbh9/7DY
Szigc+EE7bPP7om07u1QfxX8+TyKt1xX1K6IQydlC22K27Kp9I8QR9ctiSN5cHXQYIjLokXZ1CC9
AgXqGyAYDY7LSbnjVYXLk11I/ETjnMrMNQp1YWOQnT8eAa+a5jb6jbXb9y0fr4uPcBMtDb2idIAj
Jo/KWStbfuimZERc1FvT4XOsW7kueYQ4qwdzqcXcFSfQKAiKJUnYKT5nKIRPrSqMlWmmJ0d/1Uj4
UsdRdgeAFGLRVNLs1oXgFOXYrGG9/2OxeDwipDX/OiVudZkH/7q7UGrxwFNrbWpZyHjuwLT7GcNY
u4CsYu246P2T0GHol1Zy8T/shd2T5lzqXSFO10OQztIxlMsF2ChqGKCkRrAoctMvG86d13lmqfox
7J06tdsds3O82sVRO8zNuXheD9NGiAKnvybsy+/lB4dNnbh0QUy4WbdinbVEXnlU9WlUDyq1qFEx
Ko2Tz742FfkbawoB0XNRq4c64ovOfEBm92WZxG32LpZXMRxlNita46MP0qcf9TKP9XE8axygmB9S
SmaZ6ZZpEest30Ce8xK6ZYopl35Jwims1em6x0GEq9x4X82ZZCaYfdDRxlf/ykYaKjLf3Z96Z3fB
r14cBEgKcthgKPjHtpLCvI7KnFxnNZIFi3PcCjDUdPk5MuMShONt9vmRiU7spyvV4V4ln4Oxj5wc
W+JxxTiYYhKhjf018ODJhhNSArKH9tU49OAq/WVutk6oSpLlD8PLF31IPLeHFJdQP/3e93+kB3T4
bg1/X53JXB8TJ1ZHCqX8CIIkZT3LY22IA4b/riVrb1ecjE/VREOrz90pmaqGApB5Jg8/W4lpMpyV
KQFcS8jB+7qapZaBy5q+fI/fznAP+U0aw8a3m6da4ya24GokZkX/ZeO39+hfmfhUtLGiqm05lIu1
zENty8LHLX6LD1Eo+9BANZaraKBchEqByX+Q5uQbVmTcZPktgu7cMKQIjrvZ1A3VgMeNcVjDoIed
pTo47TtYHMVcASzKIG02QFTK6pDOzDcqoxydrv9b97GTk7R3Iv2W1FO6fsXEd9HSqHhATd1sXEEF
V19DvSzEmYapUPESmuBPPdAFeCC0n08uUJldFaWuAOUPy05cwk0r5x+/bEYnd329FH6XeOOk2A0k
xTw2FsH8c/ws3WgHVzn3x27SqylIPJEurWHSEtjxjVIh2WgsfecwiUWxcv5qg6XvSkEIaksUveIZ
Uo1ZIg7MhJYgvfUcDmmsonS9CdoVSSKDI7zwvKCJAZzga6byq1H+OAGpe7MXHvaAp89YcFSuWrUl
u2Zhtak8L3nseRazWqjbt1XcobcRptGv+V/JvDTPFipSUTaUgkOmEjXUKaZHZQzfl53Uz2r7uLHt
8SsfSIfhrEpbCFefhVvf24MORt/EdW9uOEig/qhktRrvd2ajivuVlrg/mLcrQwOBmsqDXeOPjhC4
abz7FTf+gursmxx7yH72fzT3i+f2xQ5Dqk76FihLIjuZX35YbQAOyH58siYwsHpiN4XuEraVm1Lh
QJ/My0aYPT9eEiGUusGS9MV5AY3H44M25SGuuPdvc/we4nQC+BL9z8jcSzjHuslbCpuBEPiStIMh
IacgMfkoIqcCp/dVf0pv/iFwlXA3ihhNOa92NW984SOZzj0zDxX4NXD6/OYB9AjNutorTeHL6b+n
gpxhB1rsvgBbBM3fbBYLaiJCtQMv3zRdcnzlcpn6IOTagh26/RxarXb1JwM/OWSWUmOVCw+EjSxU
YiggBzp7Qjr84PQJq1yHeEhX6nlFOVJMgFWu6hlzz2cgvOBYcRSnfgxuMB4gZqlJgqM5hLpUTe7j
Y1GJAoUTI4FyX3bn9OvDWW3LbUGqf8lAyKAiVYMsnFTR3/XebEFnaW/XHiKo/kxHDvSPN9x+Pti9
Jn2a0hNbLIe+abJIyh0fLXe5kkMfa/v7Ezp46WfR26eh8Sn2CXEaoXH6GA5uC7F5WvPc4VHc2xdV
V7zR25wf+MzNmZwLYABPah0YjIvFkQ9CF5fTOow9vRgc6v3lRrkkD3F4muCadhB9D/BZsdV53SXv
i1/POIYfnF+RmSGT0Q3k3IsbnbmSdCQZTUEDbdYAQ+BoABz17VHgngZr9zlCd74OZyExo5h/uBao
zfg1A8TFaI9RAcxXY5mdEUc3RJz1SYCwM/rlGbifIOpiytHUwrJ0wX4K7r3UZZ7ubloHiZ70ZFGe
StKE0K/qjo191mDbmsXTckifiSTxS6SMUGy+HUFQEURIcTXQ9XeBIHmPiIVi13g9a9P9+GPiD6Y1
4b9HXNEvjUZTbXhUaGYrWxM0N78anJgp0iz65G91vHx2pHbGQilEUTvwM4Yl4xV7lIAB76IlULHG
Ju326/jdTBBiS8eKuJGR8ew9tJMSTc9VVz478yzpjUq8jLY7zUZVBktO3y9fbALnOtcxDJ7cqt3P
wORWY18QA5q/f2dukL1ej0E02MWOg62YfVW2q0Mgp6G7r3uxVxDaJtGxK28/QZP2lGnoO/2fmAyG
AX6goy/LO0W/zQ/NOdTTqv42lXe54aecY+CCGsGI5nR5f6cYqtxVhW9TJB1AlnJEpT/vSTARkPr6
gt4sRRdzZ4mah68ew+PXyKK0pobc4BdBMKmxFkGV6mfRhgt1kJ73fU94pEdWl6oUzMtYFQtpEQo+
LrjKRWa+T/ZcitBr3b0fdw2/x+VbnRxbWf/tg+3+NceEZ70lKHKEwAHNMEvKF/nsEv20tmIv+bkl
UTmnWlRfJGwDn5uDRXOGbujekPHXYWTl65rEXuUjARXenNloRSS8mgJ9R8Rwzgq3dDamJeDULkH7
mkjfybsIgEiB/VW22NhWqRrYh8ORyOmJbY2A+UK6vKwxXbPn8vFTTBn64q1no5nr/vgj5LedF6se
fxTBHxZF9d59fJiubhhbKvfX7YrsPNUblZR3w0jJTCk/ggPpj6UkxcFK8raV4XlqsGvfZoDR5Jdg
vST1FwFXy9Kn3ojfM/lazAR0vJbyDQubh1c1wdSAeNb3hcXWEkPCffkkwDPAawVep0UjYLcF6jFJ
3TITVLZu87yZffFV31DQiu8GI10dHf0RUzEb6drdT1Op5z8VOQSu2l50aKWL1ow4HYavnhVovkif
993pAbNO3WfYP0pMtuL7N+HVSbDCyQ3qt0HgLP61eBzWdcy4UPlU6AJupo4RLymso9tsd2VWdnwV
JA7iNlHRXd22TaUXwrUZSvQpaMIsN4A8zTfXhgbmKlo+dolglKYcgmVTou1qsPXeBGzBefZSMK1Y
JAztveaOSmlrj42+mmhbLz2TB+s6OW+EGcRvwhFuxMjRDPGFQtaCBY28Ya9rO03VV9wswEPi+d6X
MHjfa4gc7Dvsmrkggm9AHIAL8dNzLUevFlCNfi6740p+g9+tc/0oCvrjroCbW0oKJ+TM/sYjReaQ
XvI9yDtG81MHo+b2yI9oYfNUWXlCWIdyUp7ps//sluI8e+Cn9jMYgr9LYubdD3tsaQ5DzIuR0yh8
xWSfNvt8zzuklsa2D8uV26czn3g/L55dkwM8UqrT5uNBojxvo5p01nzYtnNRYkenY+ACFozu4AVJ
j+RKSJeT2/xsF5qHEcKLsUAfFkQz+WlsxE+XUV/6wbJ2ipE5q2MhDHWuBO+rveqDCC9k1kaE7YXy
5lVkJW0c+UBxwVc7gG2pa6YaO11DPlW1L0e/m2/ICgLIKiJOPSK3UZXKVHeA5ANWgAdZuJP5SPvd
EBmCrOJmiuKthaRaXFtyc4ozMkKVhJXY6/Tu1ek1+HEtke1KBLsvtXch6PpLH1ZSpl/5auTU3h/R
hREVr2oXz6vL7dZcCON/yPwE7hPEqKqw+YNa6Xp9ONEAIKLuYCFy6XJo2YlxvYWTOdFSODrBu4Hp
/lhUtkNwUe+W9GI2c6n9zodueO8aY+439MSWK/FqXTNsUg90CSzjA3sVRgW/i9+b1y1edWeHFuXa
AYHoNgkb099QigpiKvqnSEOrN04KTfA+ViKPJPkKTVZcKMjC5I4Rzn02QlNwHPmMyS/XmqA+lApz
Zqf2fKFOITpcgBQr99/LAc45UCUPaJBuhNyViQH2lx8vt9z5+r1GEp1PEMfauPZTGIDnFDM/BapI
XhX/YmlzlVRbQBawzn8lO6NbbN2/ScCuHXsw3B7tItAPXOAfsx8FFGWhcwx68aL39VcvzK6Gn9zl
bA6VsmKkX8vNJBksfvhbHPG0q0Z4sXvocbGhrvAMrAJXkAXqapiR2hAT1t7VwjvsXFk2tLMFu+j0
h6jNzFASS4oUw5VrybflaxjxpQg+VUt9km6IFf94Lo49Dv6H3G0tecXpWENOIZ2lNhxZe/ueWIOI
WPnGMLmkGZCZ0QT84wqqX6exWFJVnBY4+9AMtuyunUxIhNze0gKVdO/EbQ3P8nP830RRlU25PdA3
A8pjtJWEUgfOS53b/djN4Gy7btyUPieSVddhHdrcgIzhtl3FUtvCb+VpfBa73Rc8RO3Vm30m9jAV
zknQTHAgGS7NfhYUbFgN0BU1okj2VvTPECyUWD0jRAF+GZzqWqwQfDPdQQrw4JRFRkYAFJvSfSxY
SwIu8HKZ1s3pVewNYoQk8mR/yz9geWs/YRPJny9V9LnvBO8DN3HtNNrdo+YuA6SAT7g9/kFkXFbv
RftDM+7Ol6Mr3Qwir4eJyGxZxHwAsThqd/xWZRTBAAGzoh1OUdtGpLzHGunvQIg/B6r0iXCIHAX5
+OFmhzHySfMGuAwTzzSS3dyzMemDnOouy8kaL89iTNHFR6neNfBaFP+42OKShTBMDeuAdl89Mrms
Q9qE8b/fNNQu+H3DkvmD8a7VFklKeY8hxn8NDmPVJ+U7D/65U3LJcyPysu+aNOnfDYcgtZl26RzV
YDFcGpNFSfG4N9wuWyIbQZBn7A33lY460Tp7PCNUWw8KuNdg0NYR1gggRrtFP+9thbNzJCTJwkMj
eSCucv6bd2ylXa92/hyTOlR/pX8gf/qdBCLbWDfqUYo7PCnqU1ZfxtYTpZjIjBC6E4DkXDKuVT8D
KI7yvGDx2TF3jySlsRoZcnF/1UWprGx+xm8s4mAhmmIquAO2hYBXFybM3X+DHLD2DW/SjjEaC/ho
6uNEHxMQlDe3IXniSMSMi2i4b/YqYuehI4zz9c8ueKVZQW34f1e2Kp5RGjEwZMqowwaL7bcJGSKp
qO+AcnQI02EmM6CIqzI/EDzLXp9R3phhJ5U6x7pPK3jcyT18OjtQN3a7nLPuFJFqFSCGIcjZX8pY
A5eQ5RTlj8F3+SNajvvbwUSZNCz8BtX6kE7oB9W7et9Ug+Z+pXhCM7h2gAMT/GxRbqikd4Dd0lrq
ckMVTQVpl3F8HcSIbIbAfrQOBFcm7MhhIL6W29RGW/wkg1typiSsHrm/NG0lqp+SAI2/3fPjMg3h
u3EgzZzUy7SmjxUNx6t5YhYdyGgSvHQo0jM9M6AHktCa2ZqzqEeYKyLPJld6HqK9pSg25tUyPLvK
Td931qVPuvJ/B6kjcg21PKgjARyXXotn9koHcMt0QN/XHVoR6dl2bCjA99M91INGGspWHBEuUJ6N
RR3zNfXh6Uj6c4zcb0NXhkguk1n1dQSjv6fZ6UKwFrgvxmNUwvXUuZ+zme8s7WT+oP2UrzlklWaT
Bd0bekxpmFVl7kv8C+slXMWK8cmAGK1XMp+i5wXL+babBGAKWETyIaRzHH6IBQthmSsXBrNLg78I
ERAP7Dr9oEx/ccftLTlzuhQf96kuXC9NlKZZ1SDBDTmOFj5P/Mdut0uyRUaQ0c7vL5oaCJOX/tdd
Gdy+JbLZthZV8x7uT9fkJmlJTUagbUJXNiLaUsHrU8A1JmnARneXmstjt4QVRBbJA4TCULGuEsee
HlGl9C2wTCebO8NIxuqPMJIqVnUkOkVzpWcXw16+Ptum7ysOrHiE7FWLHIFnSbfUXqk4r5p0eneA
l7M3v+ul2/ZyV62qIrfmNlJSWFvu/1ZSwanCvPh/oChw1eNSB8LFCMzW5QUGhbpibzCtsjJ72w1o
WS198j3SwwgdE0juF3y6rGAebbD+W+Tz7T4o8YJPDLHJ8L68MBiDRzNbgAU1Uw0v/k5FWZ7surXQ
VgTnniIrbZcsKebMCyG04/99dWeShbpp/wzOB1Kou0LW3T7Te5hulItyS6p7bwS6arEkIiWIGi6t
jkSPVvSEdOxAwEBPPKMiGw2mwU4TnOGsR31Hz2w/9qyI4ylj5kIq0MP/d8YHdXljpRyVemF3llqP
PfVap3GTWmKdJhP94QvMzaxizrFS/E+nycDjamIc1jl8D+XW2PpQg9ab73AmpuPxReQQqZV9KJBJ
4TOzGzERfOZo8RcURhV1UOIaR420CEmI6XFrbHzn74Rz2YwNnu9DtBPJX6+n+n7jKxFEmIWEoLaG
edN6fox98xnmU94os7dSJ5lD+PVZ2kh/fEASRklMwXSCtqqvd8GPMGOdL6zheZoVyUBR3wMzEybi
KH3LA8OF3zLZNOrvNWvxjivSjh7xxfurSWx2KlfAb715nwK6ULqM1gGNUNWpQA9AXSC0ktth5R1w
dliNtMRa6ufcz3ElOFQepLUGxQmovIFFbfZk/4+sDibeW/xButBm7ALD6s0s7V6xW6s8ybtPw5Sg
2RoYReZuadEDDob3crsygUgjztEdCjFZ6IOuTQHOriB2l04F2gAH57WIZlc4ClX/jqsI94UtH+k5
wzLUxjyjMRI4ZK0oUoW+ZBZGVkUy4uLr0eGcB7JcK4+K9cKltZAHyZBt4rSK3eEzvHK7GU/GwqLC
fRKJyzbL5mGu8xrRRH8OUOXVZrCwBHomA02Ym9pIqyYaMKRpKWoFgTFSJYEMVXRcycBTmw28UooB
cLdzHBHzwZj17re01p7a+Wi5p80rOL8AD1WndldEwq2QCi+NAhLM309SCwZzsYWtHa4ZIYeQAhqT
/vG4fkni1wG6aYXuV2ZWcuPzliM5OfXRxHkdD5orY3n2M85aV3JuezYZcTrhQ5KtIfMmUUkY8c5C
xK1pjbRy8/JH93htWva7FKShckntyBwt/Ykin0x3uQIOQlpKWS1wAEGbHjN4IurxZ0M/tduVdAHF
xpegLxGMgJ0RsdRq+fq/zg5ftS2troFiQoe2ztknE9fW6m2AStNbREDWTsYXU8Zt2XUsALEcPVbO
DGOm8k/wSccgXSmW1SPaS1wIXtwL53DxtQqfbdm+WL/MQO36o9nZAw7tTgE695UYTzTLmfTbLJil
Ak+Itw0PidH90dWwBbkCo6mSZDpTJrSY2Ea9i8Srek8+xLXJiPzNHKEt7ijdbNAgrnE6WLHY/a3O
bPU2rGP5OyTCP0DlrWFwswROHazAvJyqPGJL3HVVcwBcnQGglnPSJtbfh+nPrg1+m6/IbEdXIgfu
ZUkS0nrfCFPtgCRdH3Zj5TPhubyUjc2imKDu6rvM8pOxU+bLtjEtgrSvY9ExKmCwwlslgQZfyKPe
X2+S1njUNcn88W8/FDXxSLZ97BB6lMS8+MRRxblaXrb+IN9dzqpItWSLNCu8ikzXU+mvz275Yt97
7oaJ0kWGJA2WjzLlLHyfRtzmxx5Fi5FmLFrrvDkTCHH7gpiG7pNBAQFUSIZ6gtYvP2J2tvIWBpch
RjKZBrE96dmlhaKpnas/dRGEKcTl9OoUoEKaaSmcFrqfzDsfYsSKyzGkOQJ7xNlvt7nrtJszGBCh
GvxlNASpsyBbXpJc7Go3msH6IINQFTOSOZZaQYPFxlMWPA+wsKCb8oP/xmuCiuwbzxh5V9YAfscT
huXHUStNBGcN5Qkh7Y9nU5uXnrxsUSfJGHS3IkOw2dix72KZKucKd3ezoGoxKW4MVH7L9xZgFF/Y
oS/cvV3v9n6gMvgXI9ZqFsiJcJYmYXshYGYmkyVsnwipdmrCI+fHryTSqS5QYquUQ8KD1AwIGomX
DEFzSXnwoyeidMO6ltvgqLOxl4mLykyVvTvNgY0VvKa/XPGKrtZkwPtsR6ixfrweVLyEPNTznPLP
moOqNNgrbcvyxxrvXTq/fq9dPclq5YWhLKtuMU0jmkKRhxHa8SCSBWa5E2a9JovWcvlslOBuEa5m
+xu74p1i22LEYzhKIJeB0i3b2kJBBAfBXufAbfIaAuC03niqQZ+u6Tbw+C9Np6UT1rajZoM2jENC
h2ti/RP2nmuOgvs4niaR64OwIRI8JEoKjH3BixKXsLurlisDhOQsZYhV4+9suW6ncksBgKqj/K1n
3Ln7ggVUJj+2s04PuaTJavVHPlXhFoKBWoUq0N3YfJj4ZKL4JzLr62OI8iAuezDVhn/SHbc+mfaI
fg45SsNQNmeBeoh4HysCsdh4rxjzN2QHv1dhgZNyoLt3Hbqj3T9d5KdSK5W1GWHvyyYRONRKTTuL
UUAFMZrt3q68IrPyirMAywyMteqw2X98XZBZhs9bKRxhe8wpdd1Xf1wMX2emfvYzOfV3GOc+qlVJ
bom10AWBoMJzgYJcK8/U1fzOGMTl45j5qiH5Q/FKLIrdqW/oTGoVbLigN8Rhve1UWz2XiLm3Zz2q
rAVoFKRJ5qRsCuKIazhhX1DSHwAztYu4Dp0URHKtfGpCu3CcxFOR90NpGFugUe7WOit4CeAAcc/U
UYx0i/OvkoJ0Y/xrstRlbthZtBSXTfAlcrzS0F6u6b/A1UHBgrAE1TWgZCqmz7rRNCfHuc5dS8oJ
StzVXU41uKQD0vAhcR3wEaO7+NOc30LnvFKZLriJfwWiA+BIasv21s1kkZ1iAYyb/Ne9EC0jm/5G
s2qjONb/k7i3BB0PS7MUrNwcBZgnk5F8O5CEF/VhB85W4DpXa36mkO+OvhFtm6d52aWQmikAMXHj
gU+bf9SCdH0j42muLEtbSXipEVVWP7kG4F2+DkLczzxTX96sQEdv7q67e8AIHzko3sSM5ran7Usq
q4HcPTzDpATUnzZotngjmmDBB5SF/zFqaI5d5v6UyqlZQWSPPJP1rukLvKrS9NnBQYiRdQCTJC91
HW5oqPZ+rv+QftEIx43pQndBnUTody8CcZuTmNqlbBj8Lcqtts24/tDbYfm5Kd92qE/9ZD1uYdu8
OhLmxgrwoGfV8GgbOPYH6oHjxjmQkNsPuke5vDCB0TmfpBwNGYoiRT/+dPtYcTEdq3vBx8Th8zmG
+WS5czY0Myo58KtAXAxYCZLtp1LUBDlEXl7nn5mdciLOaDMQ0za1gK34ofnfg7LX9OxasnU6hDHz
aP3ij9P/QkNW4m2D6H6d9WLiy6ED5IoUAgHDbbP21L/5v6/Bqs1kJvuXjja8OvW0b+3rbfozhzL2
dTEcmQ/lrezFgm9NxBoETn2ZSEB4gdpXrY6dU8PAHzVL1Y3FlSH4z0y0QI3Y+pIkGZ7N1SmwE0u6
rOzjQCTq5BiWmq6FFBbIjQw2b/4U1a3CWrtne351dVNcc0n7Svg7Ka6kgnlJf6TYV40wFPgvo9LZ
ywpJE3ZiMoV96T3dRK5a8WakQN/jrEskXr0yghQ9sOFDo/8lhB0Reni8CgZasiSVqwI9Ww9/GqN0
Syl1QslO895k06zzNumMucqlTp9ih2IWNmKocky1owkpG7KD/XARPn3d7iQZRt86LUSiw6owFk70
KYKo2cYyDFpCQh/eQgOeC/X/yuduG93bxS8QF1TEqBvEMYHi3oRLAO2kdOj2vzTeUSTlMFaq0YTg
fd/HRiQwtWjDCj11aryB7RFM1PjVLm7LcL5+1wj0l04Aoz2LGTN6maWK2eWN2iocr4IsyTGVy6DU
AGqY+da7UC7CnZJEE1D2mubd0cnc8Nx9q/XVnZnbRZ25RmLpoz3VqSootWTY4G86tB1IRjWMdFVM
JOrvpyHX1nrO4ho3U8uchU0uU23amX1IUNgC7iXGyQg+aQ1mQqRhBWVq8TQraaXPGreJ/3rb5D7u
P2D/VemRpKTjJPJCYW5l04y1kPOeGDGpC1G4PFLoNUPrav+Z5c6TtcJGmU7BG+bStPK+3mBW7bli
qM+r+NU7y6Dv4c0HccjucNovxrcMTvXQiSgrCHQl/6M3cqriAIxccQpjk/JsLwNymvHDxBKlYlP9
5X8gVVuVSBZ3IQ697F89fXhCNWRNWVoWuh2q+wJCPNCzqykdjuVlC+LmoylqnT4B9CM5IjHwC9mY
0qSFX+xbGS1ur9mDr7T8nFGI3PMDrv5bEFPlNh1cgTFxzqOWp7CsKANiDaI2Rlz+uhVNxwH+eyyb
jjlmGelDwXTKticqxs+aFW7wy737lAsiZ4hL8xfGZt+MpkjtUsW+nS4DC1fr0hMSZx/EYUh1bdV9
oI+obKUTg9fb3chGNEOfeiyLlk+Dm6dpL3QYpFXfolTWGv1d4m+nfcFymhjc3fJhNg5Yu0CSn+KE
JsUoIWnSgW9zxDKmZSapF9Lk3qP9hrBTGqhvoeIWkSo/MXCeKzHvEwnjuFuyezCgxs721uKIazxF
xV3i8GIx2QO3mTvQUaB02ChSFLuHyu2bcQGt5oZSr2yxb4tuWp7Gp0c0Z5BAHYQTwDHQZlSA158M
dEzEsuEiJGonlBavtlo9ktTPgNy9qvO3AMGtdiwbHa2nhnWPsoxkG3hIiQ3Iv2wJYRCbQxfgNJxB
U2Lb7AMEgmJXIglrM0+LJVuoysNG8Gu7ZOLXgm2Vorfsc5+QjPpRxBc8KmgL9fh0qebYxf3rntDX
Pbpg3+sFdfYlxZN5mD/HYsTZ8AsQKL709SS6C/iLygKyqHfqJL4SJJ+B5NNkIKUtvRrmeaMI3Mbd
3rWt64kyebAMoxGTlsRPfk05tvSwZGOIauE2RJFgkzJbayA7UYFH2CZQcqPxDp01VdTswPb2mYrR
prRMjQZR9wr9xnsVObbwQ3aC2EEWI7kdCQU5gh+lCR3FfXAcRY5ziFG1GrRzYHWlTN6smPdUISjv
HYNb0wZVI7LUIZq0BueZBlQ4xzjnVhvVjJofC92mqf/xyjxhaw+dcFbeeIIw6Jv1MdYkTHsNNk1u
empeuxnVXDWQ8z/R3RtKCERaO9pytoG9f0ZjvpH6NxRWZ+WgYJMP6rlXuhPLcbC4CT1L2VS4FaIo
/xjS3v/tyodOOe5mx+QFRSQlmxc0/MZWhTqoD1yS8ea5ZSCf6egg5kidi83FnvgYX1/zM2FBlcO5
y5r0TfvgOZCPTI3OkzI++QsAQqoKWXpyCiOq8V1cV7hWp3wO5NTCFamW5BOyWjHFrF+n/JXVoCU2
dzl4GdZzZfma+5mFOLjNpdFEigkOX/+TXh7Oh84Mva6PswGMnPKP5JPiNjN5AXrLK5VRlllX9Clh
6rie9XePufRlcblVLpt9ehDQLjWS0Xf1wh3oYOmPjEwhjiUiv6WrO+FVv6ulTXvW+z13ElEDK4I1
mDxVl7Ag9KmuqYXK2XG2LTFzkKjkZuOmxJEAftXLX1EuSPJf+LDgd1skzXatnG25u8qbFqMW/Vqq
C21afjNSfQVnjLFNwJ5TNt/cvWlsYWM2hVPTY8r928F2NyiastcrZue3L8mjYUCkK5xk/BGtHHa+
kStxik/7f81ByelbJfUPOgHHL4y3zp1znnnLxuFBxj53o8Nm9ZtMY/ls3zZ0aLiNsk4ksvNzFmSx
/KBb1/AOe8g0cW9M//+vSKVVJZTQVopmOWyuX2Pah2BI5/ht8YZcbk0zjCo5MY6nWx1RiS7X1se9
fiZOEakIDSNbclzOyuHfJ5oCahSgZg/l8MGsyP5dbgBCXXpr/XMMyZua6b6j97gTC6X4UqRIq5cz
tv+l5uoKvVkpiv/skLS3jhXd9j9QZXLk57RTOelj5wGTVbUlSSUnTuM5wOaYphqnkrwtPSCsE/u/
AL6e4xM3hoATTNH/xxcNo6C2SNcZuVDVgBVOhF9qmOGOGxgXOA5Mzjhpq4BfxxHzz86Mt+3j1Wlq
KYRuGjH+rGIP/fkxnBYBS4F3NvDQdX4NAKxd00uxadpVOig1sRMtPo3r4BfxgweMAPZoOqWJ7QCO
iqptOjR2z567NpIgeQDc+bMmx3vF6F9FxqYWQ/XYq/Am2fv4qR2Xr80S1GWhEn+2Aps1U/4QavdL
IoKb78f5/U4pVDe2hItFlHVe59MBch25AiCiUkrMah2L8E/f4lA4YqNhxf9BJV2WN8KFIoxWkBk9
pe9fG/PTZO+wjdeHWhM92UMvY4XvwaQG+SlfcNez4eK6avO7wXke+Xgl93srDjYKk/MN7lqj7jc0
TYt+hvN4ZM3BKajXeswRRZXWowpMkXkqTof2BqUd4r2boLQu53bhTHBdpCt21KpSd7YlBD587/GQ
HH2LYEbMdK1NGoW2l06LfJY5QNou++4HXf1FmZWtBHrMMOpEi4v2OXMQDOyrrRuOQDJWoAYA03HV
qCjXznlKlA3E7HJEj6N6KXmaDfnYA9mDBYDYRWydSsdXq1AyUBdUs05qhiBLAH1bQWVACJT1m9vO
syS8j/7lBvDL19KYQEOlRt1/iwzBXx3gCNxoPOVCyGm2h6dMpEtF9Yzw1C4UFXqZx8hxJwpcu6yD
CLZvGMixgiWThGvNSOLDm5aCJoeNKKiQEIu+OIw+sC3PJFlaDYTCNFIGSc1lpIycR5JKa3/eP/JT
iJSklWwRO4Lh/Rpvzl+YXaNyXntEvZ4ve1+kKCf27AbjtkuUBHRMUPJFs7g86qIZf6t1tnsDpCMG
Q/Ph/wtHDWqE9Vj36cV2rul/uF2YdQe2gw7/rVp04Y0VvvzfnrSS6+0o5WYo6llGXe/LSM/BRLpQ
XG2JjuvFDxpopDM2iNS/CBRGhrJ5wncdcYPI04Qx1fT0eCjx+sT74HUPjep0bw4AWgSgo64YQ+is
FfXLZ5NwsiXpQCRoc4pg+S9OY8/SRB5EhuiFdaOcSYT+LdaNAdyN8EgEvLlw1qFBZ4QfAisV37cl
lL1SRz25GZXXr9kdiQNkIdaabgYA6WWVXDSz+baiAKOowfEEuSlC6XMbA/uHsCzwHvB8UDDz5mPe
EOFlPOuiPBpStt6INUk1fu16+Qo5rdg/EMjjmavCeak9/Er50cjLtubU77t5xRUci6huYVk0/DdT
rA3+C5Hq4A5KMpR2ihUIFf/B5jxJm2CGgn4vKiqfafmlgtwUdDMCxDl3S8kkymGD5SvhG4G+ANP6
RIwTdB/QDNS13mUg5uF7ZcqYs9z1GJ8xIISMkjaRWnZonay9uD1DvhoqT/J3zlm4bC0xHXx073kP
RGbCZW6thIbfCf8GHetWerlEBY3tNzdyD98DsRrotVu1nmFBD4UoECaP3OvGgRIKPCAb8V3/RHJB
HiEfmGyeYYrZUMyuStRpu3hV1qvgReD0KG35SgmiPXjioTXoM24xiZeuF8k/jIOJ3g1aSkaG0uCQ
LjA3gs9GbzmEdk9T9KaX1+zfBWZMJZTTtyZGjAMNFbD6mZT1XE4aqm0+L6dqKRZ4eR/+NPzRNbG2
o1I8QtP1RjOGvmuR0TV17jghDaG6moYWjJ0QB43pGjaMhvPHZHYM18HGbSTcx5ZtlOSztb/Sk1L9
g75KIgWwUf3JzO7kgmzZo5I2/LSr3f+eMiAL6opPFCdWpI7E4K17cBfM5g30siY193xWKJ5RIv3r
+BVLtDNu0d1eVxmPfaPFzD15n5Zafqgb1DM8dlgG50jsfm3FL5R5vy/IdQfGIRJ+w/zxKVapMWiM
VnFrQ/o1naZSH48+QbNEm3sk6fqzUDi6OAO1IM9TUlHzpbWOoiLhw0M6aSnMyFv0mKurvQOgL2Mv
zKdfQxpueMw9pb/RbhL4ev+3bm5zcvQ/X3KyqWoJIKtEyGcDPg+BQhxYt4r7ka9F7Z9HxhH9jVX4
Voif3tYQsjFmRy/x2gpjnQKoRIK/A5sXQVSIA35h7dcH4qCpYeIG/+S4BLUQiOcVZLLvMSdaxt0d
rmqoZrLZOu1m3vvkSedN/T/x7loUthNhfSvxUy0YFuHUJxj8OUl+pwBupAh6ZJwh3HHTdzGetANY
QDNcFL9hCS3O1KgTq99ZJnCnjFRVAtQRkx44FJGOEjoIf6Xf9lT1igJC3nGYCWEYMsnIMNALCVYc
vuXYQHNh7MeX2f7p4DT0RazpAzFyDnKcCjoqjCzcfB9VZg9hpmc346FBVGmJclXJnY1UW4j60U8p
KSA0/To4BwOt1APwLPPSN9rcFC1BZnN/7w7JhFSpveeoHeoIBgMX1BO59BzViISGjYDyVot6B0Y8
/vE1oXfADIXAPk/zhGM7Q8LX9Cbp9x+N0RsFSi7BgZ3j0zfpxQww7qhPJJB7J0vxLNzfhIxx+4XE
tcoCQGiaLfaneBJ6Bhb5Lc5MIvf8R2mWsQuZwWR1w1sS7H2wMn6n9mpdefNpox3gGPwRXDL0/hnb
9wXgCG/TT0pztPa0NEEoA9k7x8zBVupOPlRoYDs5VSkkQ+c8NHExPInGNpWg8p84c8jqizDTrStO
hs7tJu9vztvioiOvkcKqF2riCdRNwYZprTmumhifG9ciIf7d7MTvLZEC0KbcWDGDdn3oyBYd+y7U
thbYV/UeLMsz4u/ckcm0bCwZtVR663DaO4EylBH73tI0jD/Dy+3T5Z8+qpLBegydgXPMPo2GphOx
VsYjswh8DyvSkdiINdEVQFI4ZdBodujyg9e/yOdOozxbsqiIBKwLNQxxiTriQSUjB5tEN/bIT2No
zMxAs/BQYJFHQEKydRx3DTKWjCoPDMNyz/8QK9raSUVu2r9puW+vZX0yDweGj0nAJxK2Z22PbyKM
ppcyplr8FatPOfYn/Jn8su409kGUhDy8PCuMOqqmChUa2tKcsKZM59my0PXTcl0X/N2kTxoJyWeM
54apjgq5cAWDqtmXHkPhi+BmUumuOLHfg9kdnVqc71JbIGuBUfHAa2nIdxCizEruAtxLYfq30yBJ
g3H/OYrx+dXTDLLrXYsFXPzi41hCtM5264HTmI/mj0cZ1CDjUe/w40Nwm9hgkgO4+b/C8IXB7Yhe
4cn/hMB4JCLXXLzBq0xWvot/2Bo7DHtV6gmYg+vVhrrj5DWtcKAUk4qwwm+So+C9q6YG07yAYNOc
ooO646hlfCcG3aJ8rDqa3dIaRbqdANSh6deLn3jcI1QO6S+hf54Y74bKftap9jheF9YAfR7PJqKq
3jYJCxSkcwMHNu/gkr6nCgO2gLb7+meOVR0Yn4f1/EgOLX4ljIfrOR1T4/GslIsCxgbvDzB8+3JX
fAyQaiIDLiswBiCewp2lgbqb11juWLW89eafgsmIv4BlPJEXGuZKH5JgXxKxx4bl0YRB4RLD1bpF
NFIHGVOkW0kYt2v8uVQ2DIuBOQcSjttImIRUNiCGqTUk3FoIL3+2nekp5bg2BkAUUbyqKYHSSyPt
QZ1hJDKh+4DXBzXpGAQIK/9Ug68NjQOMFQLL2GZj78D3U73/9zmsLMAdO0IqsD9LkoqOdWgDH7OM
sfcpzgH6fCfuOYeUaMGFiaL14KLGZdFMvoaI1hD6Z04EeAQZlZF+Wt9ZTMWhZCpEd2cY08XZyLq5
YegYQQvFglOzu5p8aibP74+LqSq7ATrFg0C9EPOMw1Bj2lgBGHH17XFT4DDO5mwWTj+uhqYU65IF
RY9tA6+7JENN5rCwViiepgbI1iVbrCWTPFYHAm9aopzwEXukwxcpuE9vEmzKTZUC9wu6EahCW6At
VY/qRTWqw1zz4Nr+SrUREDLzKgxNOo8KBGVuBGh0bF7FSzlXm6w+8HKx/wSufNHCe0MXh/vRmMa5
3EU9PIY5PxYfa/xP8K4HeUXh29KGmjsU+Y4qXrzmKnOcb6bBwLHpI9XisYEtRBvxxrleOz0v3mI/
QsO755ffyBasqWCZL2o2yPrVepa8lcJ8HZQPeyuOi+MQP/h/FP6JhJBSAvHtvDhj+j1doi6EFUOd
4bZgUvxmHqN5EOIdqGIM7Us6hEYS/ZXK39c2+9+2MIRLNBDfFZuc+Wkv3y8aMDIblVRlFyK/8VAp
xfmU95saY9/+Idqu6a2ZAY6ex+3Q38HWmYES1GeSerov5sM0kuaDcLYHW5yJ3OlaE5PeoSyoCCx0
5R6BiCPdHJMAxqNeDhEERHx0LCHMtDmeZQ/9w7nrWQwW95BwKPKMhHHNwVOyCWc9xY1uYhXVdOxE
R8CZpFryTtoie41hTVQnLuMUSeWsZqKzJ9GqIp4cR28WhaGkJlJeSdleLNbc06FjviY+G9PVZMwL
VyyydiabPO5ujoOHnz32A5yJj+ytXPhrJOSySMC9Q8f0LiCVKHve83duU8hoOvoXwWXY83wEtf9d
/iMBEcmqHxYbARN9f5Dp2zPZChpfd31FtKVsE72bykN68SUIUQ0jyxP93S28H9hYacO9xj8OkA++
FmpDySynpiagS2EQbprFmYshCidUBKWW25cX+6IETKTRWdhRcXuNnK/7wkVTd08y2YExzJNRZX8r
CmxOriU3tUc20xe5VpwbXM7VMsfu5IiJXtYYMb07VWrG5SOg1sL/bZn2YoAElt+ps8gvXNy2OCNI
R6D1Gr60YphDPgRDmJ3Z3aznUOkuIvd1bhOgH+vgAGfgh2T6kn6E2uHxyonoNN2Z9UvzMmFL//eY
8szdySJdpvWBP+vxeET50L6XYx04A96VHjmCRXeLaijc9zEobqAb/TeKZJtGOSxD9igW7Vmwz5UZ
P9/P4uFJigptjpGveROxFlIyedOaHInR6w11AqGuMDyhFN9lTI5lq/GOzs1rxAywO/XrSk9sUxMa
TbJPA57xRzhn9+J7OmElwaWOUM7yGoZaQU4vX3+Wb71OU5FdyY9jUJGkt3k9cQhiDDGD7lmy86e4
9jqShS+FL4pqhR7mRioJHBe9aMj7oFRoEmc/jf2mTaB8NHFjYlo2Bga89ITKK+iENzftk3Khjd4R
WF1wjRM5ZUBcp8cQ+ufHY+0i+fCbyAgmqop8l6lzeJ6dgPeuZYoYBLWxujbMQNZBJ3BlIxsTT+hN
NTUnLA9jGFQqS57OtTlnKgwYFTGo5Y8+sj2GM4Z9vMas+GH0paZHhMy1q6/0KLcN41SE7dUxItgR
szgqkL+yPr8AHObVy70aF/l7ZtGcwMH5S1SVXQAntweMffDk2lLUqg/uz+7ZJGF9pSUQS6NACclb
JoXyeZ9gz2smj+kxYbOMk+V+kVRR2CA2fainfoSv422+oOlns6rkgppMlpv4rRopjeGC/g7CalYO
v+XdK4D9Pbb3ZYcx5U+NSegCKiwwabgZCHkDLiZG5yie7a7SJXqylpr/hnwHcYT1OY8U+8NCyst8
TTklKUx2pV/IEsfKumUgI/CplgK3Zk4FE/qCwsCApzTLND6Fib0qJH6bknEeS+RzdKN/r1rmZN8L
4dK+5RmdgeD1dqoVzUHjtX5/F90tkKDDj7o9PwRO0wMb3XtWtdnq+u7Bdl9bB6XEUwMYnJFzV4be
YhPQ26KZ6oEJj5ERnnl71XCT29ku9TRpNeeowsIIKaf5SNmWIp0xVFdvtXe/2N2qKbQsNl9NP9x/
/XG6uzKe3CQ6TPHWs38ah0+wCe6GoQmRnUDWpjqG9YBFTGcxcRzJIlh85H2ZvZHhKE6DLfYHvvBL
Gw3V4RsZioaRLjbp2Rd3YIsFBTjCWiIezB4JYjYPpeQ+fdO/o9WIjkujrdMib4umoRT+bEJd5DW4
JeJ8CGgXrNpiodJVGO9HjSZzXryWqfOfm0fbWDL6X6CXFpqOi7u0btMUbBAbFbyKzDn9QgWSwqDY
b6mwOYT+p6wIYtYvushhz/4PvJjK3c7+LS3kQ9b9eNBQZ6iZmVZI9kAfQvrSNdjzGQBq/GgnslZw
kyfL9UUwIcofzxi80MKxWDPGkyidKF3iqcDfkW5KOcY5R+Zsp7oQJNvN7/BHdpACPYK1MWU7Rkw0
GwdIMMhHO2/77iKEbD1cQKl49JU4u1yuPTWVXK+MUijOyn2Qj5NyOTDsL01KkcxhkjC4LVLJStVB
Bx3cpqGce/iv6yTAio/roFyP+qubVbMvvEgk2UZwURVP5FbUo6CbiD48lkpcR2FFtFiF6XibF67H
09W0Y0n/l+BFdNYTibv/a92AurMR7FhxmhzsLied5wbWHmiq9u77RvYVcZBOCe0LVkg3xwaCNTbC
NH/H0R5OV4i8CIRgq4V7OhV2WwxJA0idtxxKGvA9tqXOPwXNkILcpwBltx9IPe4zL2okSxUXj/lI
g9TueRooIO9G0Q1PA8QW/I4J4ZHe0hVlMcPeUXy9BGMUH71DrIGll2d9ETudVLp/QvGjx8TFf4fu
qLEeBkq3PjYRdH8ew2/Kl+5+Wdz1UNg9rLlhw20My2C4nBGH4GGDjar/O8ugGAAXbkK8/TD74ayI
uxpl//4Fcz3Ta4YwccvtOHK9sdTbvbUa1QXvc292gnIeA5umy8hCBgyiQgfQ/nqRd/xLMb+cl+4R
KqgrluPzMYFFZxeFj4S56oIm0GneqRpl7+Jht3I5OzVRRJPZt/e3jig1e66FD56tg8up0sg2OhgJ
uEEMH0TAFaKNtKFJhb53Ht7aAvn/yJAiPksOydpmeWJP6Q0YwhDZzxtPfWaIs30ePY96zcI7gElr
ywzASIfvcsFxzx5hmWl+HtOrTgE9wznBxwqe1V5McE8BrMbqnXJKWkbZWB7PlvNbVg+6YSc+sPqk
G+bHaVW59zmQ1E32OjV+mo9jG5GU0xIXn4LfnIWtAxO1x2cVJYR68RADbLzQ8+KY1VYf+sB4MuVJ
f3d1V7jxAIC6yYVWG78G4b2wSEZO5OibJk2CgRQC2zLHoftLVPMCwwnct1SrPcKGT2EoCldRXKX8
u9ulsYcjf9JKkGX9x0svtQ391EaiiNskEYUF5d2zYqcevmwcpikgx8RKsjFoOfIumXvt22ZPddqa
LpJeCFzKoTDDK5ee3OuH/iwSxCQUiIkuOcai57eoTKRZJsihF0StpZDPe57DKFCv5DaMGqgxDAxV
qVBhvaw2rOjpaaHarU9zxnDX5FVl8curPRyvLOXrr/wdQPoGpuxwCfahxVrSVo/ATmDkCfy9RICN
RYWzwUzAITXMX71W60eefEHVjj+hLynaWF5ReqSVTwZEpi+MvrcvWxHMHN2NCv8jLx7tCjBD+5G1
Y8QUU+jJ6wI3rLGi71NlNyZPKmI6iSAlfbOVaIGUifLvoPJkgOEaWb6vvXrVdsw5xQGioC3BcgHe
y8ZmF/AtpfCDEo+fWHuBgvISezVvsPSLlqGzFCp++d3XbZCa09lRAjeQDMo8zog3TYW8MDUmXDml
csl68f8Xj47UMu7a4f49bZDnJ31z+MYpAGapPHQG+ixkduPlq1Z6L5G84oZJ0ugYnyUIzbtWfOKa
ODK3P+Zb0XOl3FdQZuI1CpDQzFSa6xTN4pMuysf+YOBIrzIbiLOsCudZLGCP/dLfNmYuFIA7OwkS
hRZQkH9hZgLnGaUK271JkQvHiOKRfO5kW6GsKjxiqE4hZAKfZSAo18uHJvgHNNDZq4pWlSYfpHhD
SVxBUB3aff4FoS3uB4lZ3NEUJr3T+Of0qJGzxc0abKipyfgR/ZjauTguPsDzHT72fUBRX6IoWi22
dHvoHa7KwkaSLscOuLRAMHqF5ip8PQzEMPUfnRes1MgYbPhn1o4ZMkCERbhcQ0vTDCH5e7Z1a1jd
4ChBRbNtz7NH8C+dmvPXEEZokb2y0HWySr6gFIYjifsT2JFkKBYcw4WiwzO7yG00UjLZjGWU9a0b
2bT/GS5+wopLrRuSlUuUQk7GQEV5kfGN3m4NIuzqU3wQ8Yyt8P5bJJUHdKA92JELbuzSXa7ST556
TXWYpLaQYIXQMcVRfs6gLz2YHhjuxI5zXGSJRNXOz/meswtEsj8DdXh3Tl43jckvI7S31vNcAAZL
eQPG1mhxYqBaLPkhw+8ZlllHJ6Do8NDIuOIuYH1HJxm+KgTp33kZWg9i4ir50tb5XrtzKv8Qz+9s
C/ODjFzZ7miYn9sNL+vqYTNS8/476IuTT2RfUus8UvlUEUDhNYd9FAynHM1DaRzpqRT9Jj9IG8jp
XpH/pk1+ajsd/4I3RBGzauLz2jJdW5JPSG7NNyQzqnnlnN1HrlzhnX9xsoobWji2fMLQIqTKnlrC
R14eWT5ifqprg0UTjf39TGY7Qp0AZoa6Cz/Aqmx03jnwzOFpZ5Yo68IAcB+Kvq2q7LIEYqXt8h9j
c1C5YMMOxrOi9NWC7con5l7f4+tJ0C6im0tzRIpHsEbPQdFE8xB/BrpLLGnzq8K0cetB/yiVvOPZ
lM6w3lDdd6dpOQw95aYPlALN/ek3+vL1SZmDfjqXuk0G8GZFYrtr7jecanIXEA7+C5V1rlNlABMh
/F29jovGwy1VNYLhjM0BA+NUQPkfEevgTUo1VKnZW1O7ERWzc0LFlSukFv+eh6wBmoygxj3sAgUV
ZDzMagghd/MyNYMZh9cGtYLIpOkjQsVpioIVwcGP7R5c9znTwb/JHVXngo+4rIH2AetwIu61gkEg
8GTSu9LEwzVB13lC9Crw6UtDiA9IVakNUqiDRQ5hsAlCCGUftSp7az8IibhJzImtjCFDFkXraOg7
aiMAZ2EPHbNRrd2Dbv5mKZGuII2+SXZw+/iy7h6jXCeekCDQ71CoQvqkaQepdwiQgwK7ditElvTn
QmMJQ5ZwjbchIZz8o7YR+DeTkc01Eo4R/MapMkhBJ5sng+HnqhzgewizqCIpTVPLqQUlD03/0xJz
AxZW1Ii2j8v5poFLXfTLjundnK2YbfhZhkKLimTVX57CrfL8fZQwkAJTPNuYLtXmVmqbfw8iC0QJ
ywfzO++ClMjEfkEBtuQEZLVyS3xSvSwlGkD40d1NTR0cPZ2URRgY4SR2Nf2K2i9/Qu+QIqwneGq1
YIifbN5JJ+FcanK6Fx2YEfhERpfE3nRk4AOpGU7KJX1BVkZXhgviFItWfvOVvvGZ8BfQ1NyTwhK4
F6g9qxJAOEoZXJDGMXNyN2dVm2Z6jyOz6t72Fulf+omtH8V02Vk1p4gfOGqJ7NFvHVqSTCnDCPP9
Z3vmUcpjOcfIwixHX2XfirTuAd23OhKD6Szs+9pF+kWA8EhMdl1/WvI+VgpMybLJZpFJn+qC75P8
BbrYngxcvGh5WdWI5FBNPOSUoXJyZx1FgNGqm+64QPQqEbqyNeOLXuosGR1wr4+yTZEcNqB7FccE
eVObity8O7tHvFBmWaXGdaR+UthG8Aw5cxo9gFvqeGcbbZB3PYbN98Grko3q+2Xtgn08WJFyIp4M
U5hgWRnrRfJwd/5dFJS227PQv7W59CIYI+bQcbN2HBrv7TlF2398cPz2qs1ZNlNI7GFghWUAplTL
PaJtVyKSeBFihbTISr7M/0pQbmQS7dMRrs8ik0LyIpbweF8Jl/7BgBDM6AGZTsHIDYwMj2o8y+d+
B74iu4KQMj4W+duXZdzUw/2PmrWrKe5M0sDZcOtPjDimTQAmdLuZ+KHizrEA9ijoVOV1oJDy+JA2
ZKXisWBsrFU9ided8CRMFM8hw1oRAC1wri5czdiM8slVfMKsvmV9OltB3vgJ9bMwQS+VHr3ZyfFa
jbiXRGhMEOFQlsINIagzHrMRdBRFC+psS3cP60+03pGnrI9fXAIo6fphDwbXvGuNf4f/hAYHb36j
VmGCBxJUBxpkqDPPwQkZV23N84hMII28zN9wLNLIyC+F6lpU+28Qx4DSwpZXiuXdR5ClUmDZWTEV
vFfzHTxES4biF7c40/MueJ/awc6K0oWECnbscNLrXvo1jRRCH5xlh4TJn69oK5hlbfZ7VCi+QBn1
5+urhOyBUOey3WWtwUdE/qtRyDuOb2ZZIROF16hj5P9zKVGuCzagwrm2JqgWodZE7ZzPaWy24QDZ
Oip75VK/d+V3dtcp8mIKLwvTp6WVFBDl8fvhTvqE1ETgFsPeYGk59biaKnI8cIlbA2PO0FMecSgr
W6H/KVM2ksCdaS6bFaqfWi9zIS6JzeHO8O8g7bf058Mo7ha8NwR92s0qSSa7uOPeIuFSzkRJc++i
WwbgzXfl0soZi5ZiwPU0P0VlURiqCtAtkWcW+S3GhyeU9UJgzZHKlQHG7LIvP1Y10Q0Zlcu74HmO
lWjCKDQg0QQ0x1cDUdPVBrzurglADxR3Xwx2FSU/ameQMlIO+ZwmoREeHVvdEYIXwbAm0Uf2rham
uasVvNidFSHghy185zZY4VBtVY50QY0Z3q/YX5K3k27nYxBl+TjKe1Zicl/e5QQeWQ/rsr9oVOz2
JUVHSseXQb6BPSQMQjmThIPhAZ3N+kxDeINWoWEmgd4Z9r9WbLPWLlw0cvrYxNyWZ1cpiSa9UZKG
2Fp4FG9gI2citW6vrf0iKSQia817yF7pKu1hirvg+Y/2iKhel6/yxj4m0emzlYbc+gLe2Bifik6P
dlf3elEUC5QfFBjXpN8mSZgGky52/mgXd8t1Y6iXLxFRcM4Akgd5Bnlr8/cp5HUesUGvyD3MZA+K
Exj/Znn85PPrI9bgGU7WEcKp19BW4ysdxsokCaRbLKRWo5ZYqm52++Am5Le2Nk1xMMEQmyluv+Js
xyx68apAk5iMmFSdktmfHvC19BnbtV0Fkjp2cDTsR1WCkcfQ8+N5wAO/96nZyQ6hAy13qGhRO/PM
aSKOwJJTEiywCJSxd/7nTcKjjGASlCgkFTBWZY+UCk3U74Y6EdGL7WDWITPDb/6F4Z5pKxV7wG+P
kduo//Ef0Q3plbFVJcPcsrIuR+hX0nvlc5VhYGhZBarRr3CPb5hV9W0MZhO6jeaRp6VrmoFIBfEn
vU62LBWzHyKQlvNyudUKn15nYVHcNoUKvcsZapEbAl8EzXVada5RBfifkuzmJeuchl/f5L2wNOCg
/RX8o9dvxiwoOw2GcfmZ1CJ1HcJ0PsJA8y8IPWpY391jveUtMLR5fSvhnVrvqs2PI9GaiJgZIYbs
d3YGox38djCNedAJEEd2+zFTnxjrE6Sacdmu4WP0rHiq3wDR3jgZsoNvyuJr7+zGekisWcfGTc+m
YnscPw8FBemqr4J3lziakTfpX4UNFvwYXT24sb6XO1T+3tJtLvQmdUIwNvtu1fh7AVJr4yMUOnEd
Dd8W9IW7Lem9PaqJ1uT1/61dt5E12cu0ggMOLKz40gQ5qPoUgXitqwjdd0PIOh57wkY/ioilnsWN
nj4VoUwUrKMwr63IYiEoFd0AawXIuBHoFasCB3hU3EooMeOiE0DhmDeyjFdPicI/9K1YPDzVfmuJ
2pJhs+rpmeKuPjw1+WDrKZLXsXNbYZvXnEsB2He3KMbP0J42AqT/KLon/qtMGuR3ce/S52H3ySAg
+aAHuttLa81j2LHa4+jEN+RvCmlvpcZgHC20Qo+rtA9mT8wi41PmQeq98H6XueZ8gAWjoAlTSTlR
987xtWOfzls/YhonieI3G1WCUqJkCvuVmV3wUoDwVeqgS8Sr1PJc64XiNjxk8epO77yUAgq1mR9g
es3P/7LgHRyun3FFrbcOIeL+XL9354KU1xpw7Biy4XKZz5Q5vPo/Z2wf0iE+F8hdMsi4Uz2h24Fz
TKMRlRB50b8+w/qa4PCjIqYRIJKrNHfkUbo+JUZHHdqaaau5yHGWxB6vGB6Sr9x8X7204ys805SR
QcWzVWJONN0MkdUWDUDncHMqlacp5MWuOpilWvypjrK3Qkyqo3c9VBjtozk4NY26TUB43mWWK6EI
OtaJQ2i2LPPebio9ZQbpSXh/RUGic2aeTjc2KEXzlYNECLjR33V+4/EQ3HROC8Z4PAEKBE5bk0Sd
4RslKM8QTAT85mI/r60T+yYROw65grGn0fbyD+EdDRoD/5P/8CI6oBFo3f4L1tS0Q5F9WhMSEC03
ZhPkKR9FOTn3oRdg8nj2A7A+EuDmQ0JZy/yBSaCZfZbUalR/2voILipWmoE5cfIccWKGwK7Fbasj
7+nMgiJHPf04edwGRw6XF1x73ZByNoKippjkKJtz07HNl2/mYVIfjxuuGtE5ypftOa4VgGagjQiI
dTcG355FnJrF1MfSX/HQUDfjq1ff/EaMVTwcDmDyk70tPCHSdRcDUOuGzCNJOtFR22oRkfDa+qqR
C/yl/P35FiM+mXNM6FpK4bqwk8VzRMiRgJDMUDnmmBLlaD4RLYOb8Fng3P3fRdUv8+KBVqH80vUN
21k86KXt8fLc/kLJQNNJES1pkKrwGcG9KbptgGSwRdPjhJ2NPiXgd6wHxV4qkzHzF2vzjEBEFXel
Tu/EbzrOI+6nA0hA/fsvI8FL7OpXNfHOTllGpbF6Is+6ecje9CTyE6IXXTaB+luQUQhAsfHUM8cm
vTBGfe4yxtBU4fcUPzqQru4UmF4YaMCX766kNHKaRg559iy3t6a2MPrlPS9AcTQcGMhgiz30N4AM
/QYa3TckgR1hTZa5igOVwSz0akq6h43ZiC1gI7d2YFsXHJwusofFukoxTldgKPoOeTMLHr6XBEV4
WhZqdImPP0gtMxnKfI4X9NmLEKUKTK65hFlQ/3gIoTGU72tj3C9bU5vszjLwVKh4AoTMD8vJ6fiT
U01I0t06l5i3smu4c96F9LtOMNOm0/fKtW2E/+ZWzE9Zg2Khb67bHsFSRsuZEp+NrqpIg6i2GfjG
xDJMPWc1MKimJ46GaSS6vXOmLmUcjRsZiBW6NvMcHkR4Dxp8h1Xn4celf18bwavZlUyoWHuITASD
xE3HsGsZ4J//35gOqO0pLKwL58hxtTWbXtjZUuVNIci4fuwp/uscXDu8Aw+1X0O3Bju2mbsosehC
trZsZOVVftJ4zohXejUHPjFsSfissR52lWBImGcZWrLNYQ4yRzyH0qIApAbkJpi72ndmMLrGztrX
ZCVdt8wDpzTWPrutyrrIiN2AjUsP8TzeznsXHuVdhyrpwxklutWEPOCuW3XcQFgDyO8lpZ7CRU1z
4Xa5R4nO5720u/AFgfcbhkbvejBzFqptDbEjT3xafacGME3gJbMh8SAf49VSek77Oc+uv4qwRiUs
ibOc8gc0bOzbdskW0CQCDDNezHqgY2KTzjOlv381SEdZzqcWTvBfU0eFXnaRu1QZPq1QGVROS0VC
1GoCuz3V7gis5HdfI1ib6I6zJZWdU4lrSElxuuzCoHpbWsaaGsPpJ0NJBC1djpgX/yqY3yvcj//F
6U4wemRlJ6QBGMZUFU28BTnUzr9WBds0wHylzj5BDffD7J+jZwuQpLDcGpX/SFoTIbDLDRchOxMZ
mcpLb9D7t2oLascTUvf948s27sUkjJXYtwBhHF3UtWQSwXFN0U38Boy60Hh2i2XEpVunBVPMakm4
SJsu8PIrHXENe/atqAfxmx5FhGMp49HNGsgBhbH04pM0FEeMiM4dxAamFQN7SeQntzoKvLE7JXH7
oHpulY6Lh7foy5uKpKlzxV5nQd+NHi2Z0YsXrow+yKgQ0e86ODsGyjMz3vpDxQq9zNJtbpMc9X9k
C5SZVlsch+D9lM8e0U5A3YlqZOYUhys+iR5V1+J8c6hmEQrzq82JHD/+0ER7o632NPzbf4SzOtUm
0KTLatB+BRoD21UEIRGAYWTqG7tB1GMdm9RA8+/kIh3eljyUphUI3sx/DSPeBmIcwnIOK+X9ZS2K
8bPvmOWrLUDSNSY3AXSOVwg7G52PSLCoF69DIKANwakJttYpO0BezlbKCj9ysK16ZhuziUhlfrYa
kN7dCmUjsIESfN7vn4w/9tN2nCTXkWvRmLTar3ONyIufY1NjAYjQaJ7MAzG9NS0Pq/8muzpP2E76
Fd0R4Ll4FvOCjXt1NcqNmSLvX3YwDyqMCJ0WJEU4MmnYaDAerBKKOucT/vGCvcG9ooQXTqMIhMek
E0+fU/Jk2pVn3UsS9I4L4lryiEqcxVNf0xb8n5W9FlZMTD2eqgkA1STPmb7/3+DK0eq25qYKhWnW
jYUGChHxlnve3nrJXZFc0SlpK3VEQkl42JOfYyF3ogObN7a6KP9V0esE0xByKWlWSWIk68pkvvfJ
m0kY0//CkwvGbd1IA5gS0BZSA2hzKa8SIay73jLqlmL41gDhFEGXiv84QWOFvLZXiFzgt6vHCg+Q
6sL0TIS8rLdGULJ+va0zCf62IVetFMuRH0pnC8hf4/gSe9iiWNs+KPmKwDEz7rPIJhZ/YFPHFbEl
dBXE+m5qGl4NCNnKwcLSa69ZioSgc1GhxO88FgDmWMdmvMmYPOAQaQDp7oe6Jf6p8hN0YcrjpmaA
j1+WN1UElU9AUW3MO7Dq46uQU7j+/ZWYQlQ0xrGBL0OCD8NqCLJSwhJpa0wvMuAq0J9yO3Bqilvn
3Cfkhn6MlhGVkS2eJ2z1CjPz8lFLOgfo3BNOtiCq0jlAe1Y8BP71GibVQyAbqE/W7bYr8riG0rpb
mbj4YADnAxEi+N6TkoZzBU+doeTAsE9+bgJXDuedmvr0amHpxdHxa8ucB9MsVtAPMXLyqVULiBK7
7qQLphmyvMFQnf0/u6TozY6XgwKOIeDgEOBUNZDsxpFh4JF/IHNy2uaYmc/ilvbpZ7X5wXc6hgWS
HOQRXb9Dfh2ilzP3LtnBXBx8bkDl2963OxWuGoOlLlnQhQd4DaziKStRukzkC948JLpNQjxWvqX1
+TSp+oOO4mUo8ngrL1lokVzJrtN4CB2NaqG70LqqEsiyFe24WwjTACOX+zx3RyOpuIkcpcVhkicL
/HGO9T8uh/PAKgc1e/8qFKUgTZms+x+YUzKaDWEWBdf77A66KjC3OgwV7ajtUObOJnEZopS8DPYq
OnCzSoFmv5BiCqlJWZDrTR1gXuSpTPp7/lljpPkKOYXxTIFwT1mnV1RJ1efOwcU7Xc+oy+8lwajA
YjiR2sZp/uFmZ2RlYkTuc5HWfqNq2CiFrjYEIZ7VndtoELFjwhWbXlSkcI6D60miwWDKbmC+Dsv9
gBd0N1usy9vJB5mIN9YgxXeiWqAnGDcVlvxvdM/EaXV47iAp/qd43iPFnvNed+1ONQ/bUgFi1vWJ
KUatVcxZ/9YlJ/zxnzpoPh3RKTIanXywWIM9WIuDqbXgxUb9Kh+5ecLgpB0I8/1TxqOZD7BAOAmL
h3WOh6fRAF2XN1OaVGFZ2W+xLZtkR1Hs5XCukWpD1dQ1AcOyoSzu3pPyba6or3OdvkOUwLszF4bj
zmvsQoa+PgeLwid39HKwRCbnRsOmmjUWPqd5407pPWObqgTKkYsXlzZRjQmh58rGXIjfeTW6OzN0
eDQEH/ySWkvtWf/3Wqfpd3K30buZjiYHE8rgwH1e3iEPOBN3r4OqRH2H7wHjOlK4Qy5XhNdQEM3P
SZDQo2fnRytmj8yr/RVf7rOFBQodPUZXzdpQb5HT9JH8nc7dogQC+zTKU50/fF+hkAzAAnIdoUSA
qukmO+cUnQIHfsXzomeIUKcHNsAyu9LcHy8zm2dHlyQQbpbNPhAsN8wm0/z5CfPf4ffoCvT0B24l
lUu5koNeh+x8JBgArNYCaUlbGF+wafEAQuwKcoiYBl1jrsTAEXyPBUcdM08mfLaagEZcvqyJb2h4
4RBMbSXIKiGAqmL4Ne9WAstCenro9+gk/vF8yVPlyxn351AexwLRlEnCIkOBYmVNaHvqLRRoviYV
3Pxw48rNCBJxpHoMl9LS5j8d4EmWzco+Bg9StzoShT4MwCUq+FO2dgzO7fiIYtlRigBc0uTUO9/0
1w+0vGoxLgrmYpaRMsZUjQJ+zlY9jwhXnP9MpYLgwhWQogD+LwNHhI2qug8koZ3kBfF9Og8qmtJC
qBW/fZLuU3fsfnINKp09XYylCt6GyadXP+T8bZAje/zp94uCc5Qg8T7tPnIoV2+w5n1CdyIkBJD0
90AsmAC5TSgVS2deO2QSUP9tlXbw0uhlOLBF0SS+7xbmXqhx33fIZJFNeVO0/mm2N1RQ1upsGJCb
zyKbweobGJ7fKRZqc9JITNh5MJJdZqfrd5j1gatbS9wRnLZiaNCv7SNII4q/+ZcUhn7d2SEzK5dk
QA1h7vMAS+VHbmrmVi3SlRJn2LFYhwLbHjkEPlWlUjCESG23SmH7rPyr+56c76KZZruZvAimdVlW
TutAHkoya3jV9ihgAgO7TrgSn8PYel5EVtO/nN3+sk6yjueyVQHm9zPTT+Sq5c6F1clhivdmBPy+
+wf/CDazraJO5FSYccuX5JTSE1kRxKfumwEDUC0cnbgcVWeqFuXmh1rhOUu+TKgfKzFmW9RCzt8S
okIPCNruoOR/n6yifqBUPXdUt+/yzRkQAZnjLFUq68Hru1qkH4FUZP1vmirVyRLZEVehVv/hjWdg
AhCstLhn7ke9Xusn7+c+HqVzvv/Y/YtvWwK7gfmonUvNHaVfWBDGiqphUzpL7muwW7JWF/Vjw52W
q1vN2+5l7n2GsSL74HKYWHhjojKWBnoMC3MDaDNQJ+PZVL6c5gN19r6h85YCXAvjk6fUsvLAKUnq
bumQ0eaaT+RvWG83gDIhAI1gU8dha8bgdHqbKxJnF6/KOr0lBE9LtsYBpGc32Gq0xHC9lszwNWVQ
/DtkeEHvG7TW465MC4kJ6Mdbp3n3li0D4+sykW4vs5GtLO7qZcdmSOtdCIGyqvbXb5XbXQL4nb4y
BRqTcOdxHWcZTP4y0bxUirQaq21hGvjsjOTQx90BE7unbNU97W20ysEYBClAyjf8x6z+2s1NVRCB
pLf0w8mhfhzg55d1KL4C1A2JOJKFEP7CgMRMDoL0DrR3+KOFINX71b0kjhNNOyJP2COmCz7Rdcky
flNudvC7jGqJvp4KzQcG2fW4Q72MNMgQj2zF3JdjG2xCJJ4NoWgQ7m7eBwV5kcIilGXxmiGZD/B7
rV/TEa9sJXvIExNuogfEO6iF7dylw5vi76NnHMW/z2+nF7OhL6vm0vEnbBRisu7a1anifXohdDeu
iznMdZVooJ6vrWGW7a+gZ5OCq8+dr/rGQfWQztfK1Vc1co62ckumeZKF1rlQjvtR6rPwliIs85Rw
pbOw6Z8YVWKBS2ynkBNMNU7DWf86RFgIDs+SOYpRPIG7Mitn696o3cHN7X1DQGBBmfW/w0LhCIdQ
+DvCfYgt+nTIoWeUzKDGL10ZY69VskFQSZ27Fadx6vW7xTq2owEhR0NByRNzQ7Dvqi5w87fI1YnV
gAXmLFAlbFT2JsSmxn4P/i0DnGp2DxbGzzh7cZmsirtClgYjUnRRlxegltmupzMSAaCtxpVAn3ee
uExP3mnDrDu6LdKKlaqD6xlrMHTnqSJcs7K5Le4LtS/bXQpohA+mcH1xMK3Rp6xJdLIlCaK1PYT0
squmjJ+mCqtlpde6W7Oa7WDAS7Z4oHJt1z5ZPQjzB4qhuDxV4TxRNULIXMbjKEqLmCKAe0IFuL0z
HFIS74z5niwsTtRQYIvEDbe1zgHuQQpjt1n+iMDZBro7eNnu6bLJjeo2tcgOWHeImb3vE7ddJuPi
5UlRliOquhS6jFP+Eni3pdLM8sV05WMdlruR1J22o2XGFGCuDTsPf89nHrJmPDWFkXrCYrHw943Q
8PVOEYfZhzMw4N5kc9cTy0YgNXzmIepdMMDXDwVZaxWP+SNFdMJ5RyuhBb5T8076wc1gYTkhDifx
qgNcy+Msdt40ooUmb8Z9ULkrRLfceB6a1SZI9iv8TFhMsR2AfMEUYnxAxmFXivjW4wVQtI0vv3Lb
aQ7qH3JJ3Gsxlds1ym8TMhvHD2rB3d/D6tTr0Ny8EXZQ0y4pbRo9xpn4i1/m+0H/q8Jjg9z885io
sAGuV58K6ZsNSKf9O7SKInELEIdlUwjSy40kBBtT7hxgekvrhAUZdRHWfRc7uZc8WfM+5qrnSQLh
wGecSZGE1qFw8eJ/7E5taGgmPez9AFpSCkl7KsSq5SWudYZwKafP9WmjwMdUhrvXxFmAjoD4B2lK
NtjCYvynP+Z+48fpfCCvPfOcYfahUmjEuWYiC2PcmYU3R2A2EozlMUnbuWnZUHzXKcF4Ej7OrpKq
qQrLkfRwKRRO4G9HJY8/vDmOHQEBeOwGhcrfCUg+EHEPs48+G/obDF8tvCNEY1O/gcj5kVG9FPDJ
sb39hEAaPitjsOO91j6VykrWnVH1B3ZZ9KH/HVeZt8+sMSWImkaBp+jn8kFOgt97FIr51yzD/Pzv
6eAGg+sl6ED3bY99AhjMOjI9CbE/G7FcexaCWdbFrtjIFEVI7+mU5HztYKhP6PbhHu8N+/ryjG+x
x/hFWrt4+nHpcbjdoX+NNR/38FHx8BQSrImVKKeTP+w57TIddobafy6eKrv2MldK9uHvsRE0wam+
ipQktznxXBhmNj96ftqYA9SViVM5bLvKr1f0wO5SWEE49ULygNGAgGG7rnzrT7YZS0w6GSG2ODdo
NRWbwQoCVZx9h3TQzu9aLQg6r+8ysvqk4zo+HfsHTQtdjpOhPoEq6SXoRPeCYmnZ6kqI1csHPZbk
5ESXnAbudTOiugjOmf0Fan7dJxxHdP2/OuIN2uXBfHbnemtz0E3MCOx/t4er75ZZ19Bw5vCD7KFP
Pqh/MNQlXrBppzGSY1zo3QJHUlscWa3WeEQ/chkUzoI+WRC2vnftjtLcOv0kP0fpxVORH+YO04+C
vav56VINnZzwNT4PGMdtiUd5leN9Sfi5cmpRGsy+8t+2obPp3NoMDqGWwuplsBPmp7GQlpL1GXAg
lhkxLSm4F4C+74iJ+xK0TfsEX9WD76iHhjng+E5RhOkzc88AgzdxZv5vNJIs2cIrMrqRARJTN1IZ
gk9s7EGDWkQzv6dk45fwlYVW9rkDk94Ji9m9yYziY6+ysl5nO7PRRBFBHPZWPhr3LSt9wB/ohxkD
04+sMrdUWvQheYNzzoP9KbQM2lAPleiz+hfr5kCffNDBpH6T/ZA8JUKH86L+kz66VoRoEs4U48Hi
sLXLd4q75nuo2++PK70b+33ILkFspfb722HaqevRIY6lzNL9kCNYRGPWMwCkY8sMdqGEIwqpTiFl
OGPqbLH0wXAiDZkNEgeAuNiuIuQlhxnKwRtSl74aLwJM0fVq21uq+WFfT95d0gpA9G8q0rbfryaA
0/DHZH+QLRieHE5cWnClo5jqlnhyA+T8VDrx0EzlTnUWPMsvgecjPqkYUHIkYrvLYQreaJd0S3Wd
Q8zo3DM1EI+u0x6fw5ggKeN9JNf9IfSYorparFsRbIdKJRUnkTdYi+LlMv5v1A278QJsJz/Z44mJ
i1tFWCwa5rts69Cw+LV1jaT1ggI5b1/q7LvoNGKr1aWwz3/n5EdN6okixtu8ykm9tx3C0CiFE6ji
pEJeDdhG9PPsFN+kdCMl6bk7G7IyLMTm8O+EOxUu7I5DnwRpwf7lWJGiQR+vjBtK33tmVRExNlzA
5s1ULleSSqhciM066q5XcYrkDe2nClVrcL0k0tDhTb0gEM6N4jRX/VyTdOFnlC9kzVhGPtPB3cwi
qG5YaA42jJjmXsA1KTnfCC1V126DRT7RUq+CJycQ68QmcDc5P9GMKh5TRDr5FTciDGvikDAxDg6s
1R8OmfFyCB8dai4NNI8Ph/pjtFdc0aDzFq6GGW641IJuoH6D24Rc52jkm33DaW9ohRQCJHW5mO8f
H6WCLZOn7ZHp66qZGBk10q9gYF7CiPvTzTDeZFms/oOvjdT39c6e7bz14aIiw8ORbbsLyEJyzh4V
+95FRS+fXOnv16OxpkHZAyQB2btJROkN41ZloWQqTyk50XgouuKBc4xgs6wfuTCCSOvdEM8Oz5ZY
HocBZubr927eJO7EfFzsg53gEa6Ax2SmQK0wroAeg50Z8JYLMVYBPvxIIQ5UDWsleRjzvAxTQ01r
2LBpv23xTc1GMuBxwHFNIrBSfzfBZ8bNHUT25WtPmWhde9oeGvyg1DNWaTL+9bvHe9c8F3FKOjpR
WlkiYZl9BuilAs3i4AY3zJyKKm0TMFWnUGhLRiaqCCiF0SDpjOigwG/hkNiG6f4Uztuz4fdCyBv2
pSIKW6dNgRx5mTAzOg0KGXEgh33ZkkRy9S1vIYEZiW8k3WYBo6LU6yCQp6CF6yhseTpBH52dzDps
yekbQzfUeHTG8B5WrAPU1obXVIjjs4otI1FqG5BiHh7uXyH84rBr57WYfJmkoLZOkZgvze0nNPXU
g3PD3++etU455Mf/Y9hVivAkuzevAQgwf02DuGyA7YT/bj0tTaOquo/76Qc048ru+Xmy9aL7hUWh
kPT8HD6AkfdNnkRefd7R6gw4zdTMNGp7cK8u1xMxa0XfkTewGZF3mo1RpnD0fLtI8MgRYVYjW+MH
8Lqu+gNLdUAWfH6K7g7H3YpOjPtNRxWZyVxB5Mi0LwQbKz11a3g51jUFwaxi/R7cTWOG/NbkoAdE
y8s9AO1o6lV8TrcGzuoAuGJuPINUB1sEJfNWC87edm4neBdogVpoyoy4EtbxeT1RvxReQxOYN98r
Uk+RDvjRU/GPjflj7OISGhFEWqQq7NSEFvOxEUq8x4EdH9ZMo9geVBflvpmFiXaDjacTPnKQ/EI2
7FqG2ar2EGPHkd+WaR9S5O723IddGw4kBRV3scvbzGGK2hobzn03nb6OA2XcSVW7O/v6Zyw46wGb
VnNnPaARjRVAHjgSi8dLK3EfTZq3mZ/btxu1bXa+ULWhovij3QiA5r/YVbv/yUup2ljiZFtGhT+r
4p93yuRxNIaq0Qc4LXLyl91uwBaNd9fJ9lwuhqIPpdw3fkf1jaD4/xUohBFckPK1tw5augjBBIiB
eZJQxMROrsYdn3nUEu7x2CDEyjGz/bJ3WeVqgSku4/r1ubxAfu/Dq9z6OjZGaZyVkS2J44WgYRhL
47v7qRrKYUiWiSDHgu+cfEdymoqlQtclpbFqDAsqC5gNBANGGIL9dpT8XVnwRGYjiblg7iVafTOr
emmaP129ERS9DMNfiV/7BBeCo+JB053uf8y5m4uK16a3o6ItZiU3F/pu3CPJ7+PNQr7mGRRXVFk9
uxxGpciKNO2y9CKPI+8ZvqQlX+eKb8dI7kEz9VeZrcnbAbd6x8d8yGWEkDtoCZg+RTocJXblDokw
7slCFQM+VlopOV7fbbgGrtqaK1RhhiSe0eWHuzN0Wc/Ii7hIvlnDVrS6Qx0HwdrJehXXLn8/H6ef
IyVHlIjew/eTzb2NXlDHPt/tAmWgByA1WK7t64vupGtTMCHVqCzI44O11HyIG0fXxUigkLHOJBAB
kYdgykpt0qKtZsl7X4z5fW6VVh8A+NJ3OB9ycPiBjsfEQnrvvOFAf3X8wfXR3TK4gxC5FbdSo+PG
214moIzXOGK0Ek7qAh4YvLhwQXrGNPRdcNvsEuuoiXDj0NpUBfpzlcAYnVGcER6vSK1Cr8V6RRsp
KSNLuFi6YN86lAjOzRL6Xbhvm2lIC8r+IPZE/KHtz2RQhffgnbp10bcEGd+FOKLYFO3jtn+dV7RW
8Ipheoj4OhIQNDDnfejV8lPxA3sUJi+/0gom5HtU0f6R9p0rbrU3nPFkFdGnxCaTNDNHPJIi2N0X
zc+D9XBqNdC2Xd9Xs32O6WQOsWmLuQITXWpLc1CvnqdxPnskwJG4yMjF022vROn6xdAWpGvIlZqM
K4GeepPS6yhFqMfreMAUL4B7OcQ2UZlwlHflt5JdRPPCMz4oaP7jmR4mm5BnVPTosb6UJeM+xUi3
kOjo9DOt4WQwYRk/CUzbZ9hBrxHu3eZRnLdDePNHclCnh5Mmg/vGyzkv/UG2eivd7tMWIMnlfrAh
75LN1UQe6b/co3l/4oYWy7OkyWr2JUtQW8a/9eh7BaznmSKf9DNQhQL6RT5jSPbuVQE8oDCOyxT3
TKZqb6RWTDslDjUn2PJW56JuyC6Sdw1jDC+L7S26AThO4y/Ke5Su80geuMi8GZ4ehyp0QuUyu6wG
mCW+r/Kkd/6bNsdrA58icXCgDHZIKMCGW7fXJd6v/i9wFh58yTGf+++iAkEPP8KG3NkswYIoDX3V
lAqkkj5Pjd0IOlP9Wb2FdtSatCfeWHnfFAOVbf2R8RZiRjrcSeWCVKhPqjVoQHXlKnTeT0idaI59
LWaSL3q3SCpjv7oq90yRiuhPnWe3jEUP/lNFFcd3/btlZqPMvMf0pzjJscEf3PZ2J55+EGRIs2X0
NCVUHsKvgu0mwZZqT/81CIF+7paiSm9PByCWParWPrhu0BtInPoY9waFlTzitXEDocHseBVfbWdS
+gr9ma6CObEpYG9mQRjJXgXS/pogfzibuz0kcKWXgFb3Ac7nFDbLLsOGSL5IH02Z41+QjE43/xw9
sAHsmUFly37w6vu/PF+3WjozDT60SNlDwyOV1mg30So+/qUPMMg5AyUTIwqSgYjm8HNI9gZjimRJ
fpe9BInK7Af3f0mJptrlpsWhrFR7oc6uECUNgzxFa/Wfg7JOrLlOR2vwzHEvMdIqDpvyvZ0AfT5n
HHNIlM/zbsaLx6RRLEBhNp0UIgZCFJHa9SksSdkksVj6458p6Y3ZFpYzz8xlIhrT08QyYHeEluTW
dqQzcOxh2jBuCQqBcL36K11S2OW/IBCOh8y7X6lRwcAxE2k2wMMfrtb6IB1dx5AT1x3UvtPNBdrt
FugTDYhaKdG5XiRdneG8sjqczusTveCDIAravdUybcJN0TWWQTdsgUWVH0v7nH0Cr/kPDeT5WC1e
9UDwNoIjYNwpBEeBAx5Efq8UfSjbXkSajHAbA0Lxa2GL9hY7yKjh96NHZf7kUDTj4TSapPkpB0hX
KPL6nhOgjSoKOBrCKG94QQ6TOiBXRScE/gef/iYdiDKIxBCinaxFMgrdkx2IK0FIanCY1vxK3ljd
Q3e8vuDUvIiJBzVviTXq6L5FJU9ZawSIzj6l3JPsXBT3IqUZ6vet9v8OySeO+rBA2+9ue23X4qWA
BfKAZ9jdpEbNpzon+rjDQbFRP4+86GVwu7F97rrtzMENN4q657JSt1NuuDHrU+wdbBIUKbQsqBAL
MFJZmLRyJ97uD7KJQpX137Eyxg2r5Pq0n5yU2jgGNXYll3CX9w3orXLZ2r+a99P0a9FwHLnBdH4k
sr3fBYMdlrE3/LYFBAJ23NUE6Fy04AwHxmlAXwi2lyoQtADEpel5ZVsn7Q2zmWdTj4FVRO6mSUXw
jxD7FuIIX6UKjjqeSsLUIyNBO+1WGW6BRMfVfiD+dxtvmrTAXp+2FWvW7/4Jyy8ZLn6/9x1OSpgc
shPZpzvzC084rKZHNWO2Vj4qYC7H4rHsA8mN1M13qvYrMnL9gjZh3FwIreWVKuL4a4mt8x+Xxeva
XzrFhISNKsMuKMyw0XiF2J3FTLJoZN9hmbC7CR6VHPx2HrXSZUImca8wU5sufoPbk0BEddtM+L4R
0UQ5wBb99gxTgE6DJG4hErnh1xQxSeSojXeDkZxDo/rjEUeSPMUZ6NmTckvdyM9gAhCsKcQ7tTFh
jGIxGv2JpouY84R1Yc4iqUVyQ5LPf3BRNY8pKRPKCILNIbm77Ah1b07/aKw1x73STSa2O1HWEWxO
p1uevIpA+Rrb8eRot/mGVMrkEB0z9iIg09eL5dxAkmAH2lGQ5WBcHo1CUm8JdRYXG1XANXltNGPf
DTN/EOFc64RQ7qhEnwkGUC76B2qpgBx0QaudsJxYLed06+GxBtWNboAWUsebWC3dF6l6yR6EGzeL
n11cRC7Bx0DQDo8hFeSm5mEXY0ceHmpspXSGbTzc+s6ABHjFaRrbixiQVjFTxk54kbX/Ie/rDQdV
3fYj4OC6Mikh+B2s7z8HjyCy4WC8JhHkQyH15Auty+zopkaLEE+P+G58PGF/oz1C9CpccAl+wqqx
5NaYI1qhoIIVzBIRzKS3flcZve57RaQUeTx7mlZ3KeQ8pThDkwtMtGOixoCPYDWE3N25M6Lfd37a
8zTNeW7RacqmBUnAsvhCfSx/KduHx4zOzC1ieILPbczLCLYBkBfiMEhIxZfN/gh9pvCOKDzsMkSa
/q/zoOufrrx8WBF4YVapf6DtXs20PaynPTjHNDc/qJNghLR4S4XRPuqKy86/OUse2a71/8ciqr95
ZhEM9910bFPXPapQJR75QfG3ZayZSQnL7F6fdRKnnVtBea4YehnctNmKOpj3NVZWbpxBLZa+gREA
dX6KnjxMSsa1uJ8uKujZUx0A/5AMndJbUD0PD+tXXDZ43H2l9VDb393NKay9gXuPXLwyqjYfxqFs
rT95VykiS/8GVttavQ5pqCMkEp2WttOOHD8rewktZLfSm2Akh40b0AFlMWZodTy1h+ufw366za7e
lQ5W/TQ9efkb4RMpyb5xRlKW6sdfzvvkZXJFaxWM1V44m2BRK2zeM0fzv8Lqn6hoSpg+a6NdS+Q8
7tNMSDe85fs+YPmcwUK/XV9SBM1pCVrzmjGvBwNZv0x2ZETHk9PKT2htplzd6vW/7csmq8CTIOaj
XltdXDVV/r4tn734VkxdQ0sWk0LpBoBazcadn7/S3LzIA74s0uxd9T9DnYCreUEMMJLRplIiDXNi
0JGczTl2599Oc2105k9zdnXJ3PGx6DeJDIYf7CWP0T8EK+3E3azBZPyI2EWBdrns9OW8v5Rr5k5a
APKe2EfVrqLeM4ZTUmX/iuUrtiVfpWPwxySFsckILWDc42oKgQZ6YowrnjeLWvPga8aDSKhmfX7J
WuUMo+sYOQbCp4P/9l7an6K3xGp0fFEXvN+JUrms95mvgSr/Q3dGVk5RriWQz7Pl5OaJWhB30H1L
odgD8lMg+KIxX8D2SN2zKSmtDyThioqiSRpAoTQNt7pzWReTa9jjDMLhA+s40odmOND8kDq8s6vv
0TfwElBn9MpwXz205Mp02DMaYvMcdOIvKoW8cs2QhCVg+t9JFBWwCqzdYGYTDjToKgla9vnhHP1Q
rHWcI3oExVtFIdu4gHRz+siwJdeAHuQgh0x+YgC0MM/C2Gkq4cUlhSRdTPdVh65rmWlabLgTuXQ0
ELvijmQcQ4kjaG2jwrft/RQf9e/ubDtpbN9X92cCTcFMtWG3uoqPF/t/h8iF8YcPon3tijSGazrQ
WU+zvNKeRFXPisChmYq6uB9XGSj10b2cb6nMpYa8FUqG5Fq8O45mBZrG14vze4Bzq0jcy83hR8tZ
pkVP6lhvAUKqxocgzAs3WKfVrYygcsfHV4GrPKNDOg4mbFegz/yST2Pwz8n63tIMrE80f9LMoBok
O+Dctyk90ctgMHIkfsG6m8pti6MfTUI+XRTXrfNKLQrydZZuV7AmE0UBKRWlRflWh0f6PAmkPrdT
rvIj4PG2c6Swo5LEb48xKSy+c5RCXfUAe+uQupEvj77n/2WxQtd6H3sv2PZghzbesBg2XVbeSt47
BJwqoCWbEmKfRL6Lw/pf2X+CmZZqiBqU4TTVtiGrgU8H6dpvWm/kK2H1biL5VUtvVQfpEj63ZLR4
diBFRzL8F9mibIeazRCsb8CgY9MyjOOYegXTEuoITv78ayPc1GqaYY8kReMsbpx8z2ejZLhv3RKX
6romcgHQ7t6Vm7EIPmuFiqeHgIrSSQEVFzn0yKnTt9YW6rwlV2LtVbPj+K7DHg7N/qRMsSDaW3mz
Sv9iEcVYVUOPj2MbS8KRXIBOMnJHs4rzq34sJr2asAl0+UApmSvwgZPcAZSyRWVtgMzmKukPnHX+
G7soxuMw82vw9ykId7RWswAQK3YwcTwlOCUsVuCYQgslcvh/2IpcJ9On17WSZGBUXzgKne2xJEym
07q9vglPs8TqB97vgJ7mv2yH1qpE+pZa2Jn9oUdXqbeCWQkhZWZiWmNpCH5dhk6SeVwX/GXxIKv9
zI42BISvTV0G0/W0EA7gS4avP7LwlUAtW6NuF6TqhBaqActqS5vki7oJegh2MohUqCV40iuSPuOn
dbBTmPpwfiRV0rm6vrEbde43ruEkGwH2NqzP8G5nnysgrdhzEEqOlGXjH1rF2tJMSaf5qVzKBjbW
ghPTdZk7hmOHUW9WBYsV9z69iTGfIQGQ8AaoqfEj0eemexslBLvGlCvLtitCsI+tcmuj0IaPLyLq
Rz9D25akF37CvCSvbX9ZZdwSSSlag5D9ONaATGkjC6HCNs590EtX03Mtohp9caPq0bXu/z6UZ76b
CBAb+h7l9qT7wZNrkfQkfpB5O9cvdEh4dUe5bkwwg3qze0kUGXo1wD6NnV6/cSTD+zrEcns14rRa
wQ9yW2y0OV3vz1YBeYtqtWqbQksglDYN9j4fZNLBY7RG0mtJ1dNDE7DUP7JUP6vcaleR5yNcyLqv
tHHIJLsWd5+2CN6LwCdgXx2la8jNGA/mf1LsDQX+vF8OlKYkW+6X33/oC7vk9+u8Q1ZNC28fCers
WPWp+IRXO8Hn6NBs7LfJj3DWXpdqZ4GnBPZ02qP5NcEftggPJ8t1PZ9zDJddYxA0eeIj5c31mvuU
HtWfzPBloOoFO0FUDVTloJVVQMiCCb/kNLnueGdPkbbqouiB1wIRc5WaVbwawwkL6xc940W7H3dx
X0FjFPC2Ep9pHfwwahXHCsODh7birliTqmEK59siZ6UI060sf8l81bjzWoc/o7JR3jJWNx9LqA6P
gCMhezB+v+uQDbIGJLf+2rys9eBrmZp5THLGouQ9Ynm7Rr41JR4GsM42IjwDRgmo+w1cbryVf4CS
DE4/v1ub62xYFHf1OQqlC4rcCipCNve3C80zqgnVnZwNvXJsF+a3IUAB4CqOmOtD1s8VMZZN9kVF
wV2VG+PaX/DZCzlDHQTTmJKwNOxSH95xXCR4CNEosq8qT3DKLEcLDUgAu9fpl73H08qRNVKUu2fW
+PIUiGbDezXGnJ+OfLXlrD+OgA6B+5c+yaAzVrwsgB13IhCveRklRu+mdqvs0n15azmxYuGS+Jxk
lJ04dC0bKtuOa8w8R2m5Or5npmH06UuFco1wlGlzquNWgMtEdVKC315W0OWI7MXauiNWmTmtbqJK
HpPV1eYFCon/ZkLOoc4CBUxbd/3Zxm8GApeTfpqdvBYXdbZibAfCk26Ef4vq5B0L1vRmPkQc50w0
3idQrc+5LMTic8XilTsOrL8RsMmBSTuE6iBcbvX7jdF8SjNp6mH9qzt2MRl6MRZIdbnxbwfcd2VM
NRu5qoqaqXZYw7Cocb9EeXWYqfAF/uovXUyx33GxB/sIliL7HZo/UUIN8wyiFlZLkBdxiUV/zGvH
s+fkzuG7fYMWX7eIMqQZBORZls0fuQM1zkxKNATZLeQSWNVZyfo4XChVv1xvinocrPrLGRVOh5DG
KjMA6MP0TqkyPPS87JQa1ep4qXv2SVaY0nHCN3jzFLTfX4cvMs5lEPIyEypSa23TPqIP5nf/xvfR
zV/bPUqRYzojYLg8jShtQ56rGILV5JTSbaCYA/w6S7mlZtK4IJG/5bjgFlq03N2MmIH1nOYR2fBy
Zs4Y2HaoSss1rCCEjHVd0lS2YEILJfYJICZJJO2p/Dd7jIl2/Tlrev0tvMfVf0bvtP0xlJqxqHms
CqLamqS0E1gTCcEXzzVmxuRo5nqBBmR0bYpBQWika2r+cuuQTH+8yB0WbnCXLHcPfaUZeugvB1hc
zJNXdXaduLthRVsKqu/0FfOwGE08Zu1HiCCy/MfcdDKSOnRSAoVPtTtofH9Wx4DjPZIcF6+nCgFE
muZlVIDdbvXR4hSTeSo8dJR9annpr4vfnneUCU04mubAOYFL65Aqj3axbeTMCjFWevNLdMiGF2/C
PnHSv2Xq7OCSrNjRGHrkL3gFLLFM6NQ3yaf2e85NhmCfg8Eai3wsjJfKfdzvK7/WhSXf7PpVqJI1
LOMGFO7igMnUxnvC9c9NtZ0m20Evdj8DaxcNGMGZaL3rBecD9RYp6F5SLPgRo8dDHZfVZj2uHp8T
Ud3ErxMXkbQlh4RHpIsPzs9Dvge1AdQcsh2v+POgK6S5c2sRw79ZPaakGJK7zkvUxPF8yEu6+QY4
NELtZEeczqGQeKaAPTqgcYhbuJ4JdCzZ5TmtXlUn9sp+Nn1HYrLdo/KxkTWDi21L0vU48dn3idmG
TxSu+8ZIox7VGCTBtGZ/2LADMoY8qNhfDfSYSpVqTR46jt29A1i3q5iBMHKwiG8Oiq0lRz5TVBwb
kTcrvnKSy+NwAj6gNiXiVEk8E2uYFHFtTAdxtzV6l6Nk6jySaejG9DJei4ue73VgdbnYL2hr65i6
9+h6OqLTLoW2qfkfYNKc8SRw6XloqnY2dPXklD31uE9HkaFT7S9jfjMqzrtilwcRN2kgl2URHpgp
8HFPlzFv/ov8ZFHcKe8MI6l4gInweOe+jpH2yncCo/7unnxjv2UIRmdg62mhB6TfWdOSpdYAnlcQ
qWx79m8jREaa6GWAAbRhUoT+NoqhjRQA/2naZp6h+/+r29wVBVBvP3+v9CuIY0IjgcGKM+bjbGY/
Gj1B/HQ+KXYbH3VUQzXwLAFwfRloJB2zLbrJnL4MpoeSmJ59VRRU0V2yIhBVgsGJXD/cioLQQ1gR
xdvzUkOozftE5KBKMKsOdEholdOk9mcZ/ot6BAggWBehsXsQL3z7QpeX2MFkXnMcR4fp619GKiqP
Ox55aPf2cbiQMSPKoEQrHnJ3+opKN/UyroZVo4ALAnB8NfkBW1D6MW6atj/SGWFq53UQJHfXx8J0
1v3XjTVXg3qTk0s54vadW0hukU+Jd9AsIom42TzFaf2AG3ulaiYZN+V1m2Sri5BEzVTggVBMfvyJ
KgiwK0flto9gd8OB+1dYSPotGOhGd1LIvcjLCIi3qEn+NAmQQNhMraNwloF9d/jQTlj/VtuZRpu/
37dEUTPUyIWoyYqgOW2/TU9qYOVZRunYV5jBdPlj9j2aSCdb44JA5rOjJuJpZGmoOY+mIbu/6SnK
warHE6ubLCHIlbGSIrDRTRy165a9HO0gKo8HEtyt5mriOZBuHLsIeTk0iFuhFcmHojVukpN8dynH
ZL8478KPb9JFE7S4lRTv0uWmuQqYugID6sQMZs29ULkDyfirOqPxI6TdHfFoFn7+F1u1qsKbp9pj
Vq8sCreC/BprPS4BazCe6jAbBSsK1PqrLrIMo4tceLQvQZg2GFTihThcF5Rr3Lx5i+CfcnPw53PI
OUeAVg1QCOs3ZHQRT6QIOdj0djc2f3xw6RGkrsfDXpH9aapvhGTsiKzkIRiC6ESyveBIBNYVrZu0
b1gid20/MAtw7/hIoy0vyrXz9itxrnC0bMUJ48JrVQwdBLiJp/jd4cg30jzDbHcGOv45zbwXY8Hr
yO3UyUNuDDacuyxKVJysdizqp77d02ORwotH7zQc2yV6tRomhdLxbnz7xf4uTtdMx//nybigcJlv
S6efWmyFIJF3Fd4ecguw1IWUp/CDplUnrrIOz273Bn7Wf9qumFvRg6rpgTp9HRHbhx27yfsUQUZF
f1S6CuhEyxDqfOOEpxBVw6S+wqMyirtGPA1GhE+kfpZzJ5c5z/+VDSKwoKTuAmLrehfPw5JJfI/5
oRWi3FfM/qDS89HnofPSacMwejguiPFBRa8v7xd13pC9u1yAIjHIiFvgEtsOmQOeNNcS6ENCXmCM
lSILSJPfKcClChPIFkONFhoh1E7ZuLKec677Sji49H3REypvSz5lzk+05NEXw7y7sub8GZz6T7gR
6EdYAQGl2s+0GwkO3BfhMslBPF562hgzNh+GG53neWWiEY3ghMOo9yGj4CMyJBJYjJesfyGQlZ5E
20p9zzhzp10dGmqipoIASskTcAEqYu+uswsdY1nC73Z+R14dEP6yKf5hwo9WmRDU/oTZo8uLPIU6
27n2HevWivns0EIgUf12zqYR7An3AfWB4VM4FooUpsq+GUMlT5FLPCgvS+++pZoQ8q1AXhFBeOCb
icGj1vf+Idh1bAqigjaHKN9jqHJGC8aHa/6zP0Wde/sncPVHeTaeFDpw9sqwP/Q/9QlF4f2+2oPk
SndpR1QKLMJI7YaLVfca9Q6/2Q5zcyPsdA+TkweWjXkwCSfJKQGwXeN6kTCDCrn5fmUzO+vM77E2
TWFXqmZHFzQtyxjNUrpF6doC598U9/XP+aQe+o3SdWO+eJeULjcmxRBZJHl+EgNj4ngMN7BuBp+u
Fp8Ru8nf/G5tjC0OJSxRr7TZTwzgcshSRkw8MOhprZR/6nG62uLDNV2eq+tSKDE+TtidQE6ZkRtJ
yRtcTz7EWhBnlAPE6vywEBVsbPHrAHJtVRXsoVbx8lql2tdBWLoqUg+0I+rCGydMLsbWj8ST2kN2
JyzvhkqX09DxJFxBlsUmEilw0RFoMn48el5oJXQXg8MMGYt6barMwZcK03dZKPQEFmhcWSGGGOU9
r4jWfRUXXyMYDgJx2odV4wXcOIDsqcXlzA1qphLApEDrCoJzO/RFL+ZkLMenSjE7KelAe16XuDcv
+urT8jz4yVddNYA/veRYqKyKyA8hxWgeiYeJk7/rMtQ27gbLY0hjRh8SBauykcGeYOqhIw2ymeZo
gmYnRWLm8xFZq2iwVdzdqICU0g9EAdcnDQq7BSiBU9SFJROyEeNzRt9ijM7WTHUcHMwEYFFlH/KF
pFKGfJr4AB8hJyBTm5tODwSMR+ALrXs9kqCPGcETs1HdHhegye9w/jdK6T/NtBAZd93xJ15z/JxY
MDgRPSAgyH7nhsOk7oIROofqKsWS4qkQ6moLTXTzF7WNlXWDLpC5MzXlIVX5IDP9ju3tvkV2ujoy
xiXAZyQ8KeQgo4Jl+lW3IQbvH8LHgxBuhSF4y4XFs11aeYjBqyWijEHEsSSEOrfasN374lZhqnPj
qIs/vhrMv1BXs5oENmg/7/sVo5dbuVnLftifY2d74I2tDHf5bp4I0r/Z07LvBwdLdufFuPmcTU2E
TW/WmnjHvp7660fXGaehgCfFxMSwf+sqf8wJmupNskKCEzywkwuwJytJP4iWf4PNe7hwZk3q1put
noeEPU4e/y4BoqxRc/Zk0ttpJfPwHCig9eCa1yEl2an+aqYlnBh+t6CDpO/dclXV2pz/OcK8Kx+b
BahClnBl3tdY3qpv+kG7z0Pjb50k8zOucwPKzjHlBthxASXWyExqtXBvEGdv25aechklbVX+i9qD
vCJg9dav0DUIxw3cpShlvWA0UN+V/0DbKQ82vfULodX6izAP6xxMj08qiM1GpxV9ByChJb1o7Od3
tM91K4DiU6oQ7gH4yXVLU8+qbOqggRkvC0SLG1Pqrs6av+PIqxD5pQhRutJvFntwJaSa+kb6VtJN
gqOrFur/SQ5gNjHi8S1MFwYukmhuHO0+W4W5JOu/7VkT2NF57zCNOWuvsdDL8fYs4mAdLcxd2lfe
vpqpLyvwyM99SmYNP8XZAMUWgUwH73rcZVghU2dGPFhMVnY++M1baPQ1kJg6MrDbbRC7V/OIOqJ8
e1GSZ5Af1mCyyID3AMElrXmGaWoNCT3g5hH9wb5zlzl4j5trVGVyMduBjrS9MwbafvNdX9ZpxMdw
PPl2afIwiZ7XRc3ndf5VwBrF7Z6hkdEo/pFy1QbSAOF7I+68ZWEn8kguTRf0pJCSVcORX/3GAUni
AgbEXbe8TulJ28uTxBi2PpdQaztHqhZ6m9NwHQQnm/oW3x1Lwo1xJ3x3no1cPH2RSp1yLU9tK9da
khEX07Ov8Y0AJFG/Xd+ZVWKWtdOT7tbUctlDV4geErX2iArF8U2C4lpSSiEaxH5EpwTcZkbXTSwV
9AYN1AsRgFhM9tCiAjulU7ruBHXUP5r56FkygAsOPyrcbmZxyiymrdpKAVkcaTNwKE1aAfqrwQQN
0symZ9AoukZ/OdxPdpGiLqdo5p1QCoGZzj25HNsnlItpP/T6aJ6h+XvI3AEnITkE755xstz3M4H1
g4g+RBr2SxvDbYHt040A9zujDu+KWl8z7s0bQhVk/oNVZTG6uUxShUto/YjRyD/fmJbSIGnQO4Me
KeKiTaOnLXJ8nqQ9xNqvylu76zoKWDErnJJlOHiWPw7V93/TLPV0aCCuKHNlMZW6ZoPFZPLW9X0m
HLu4W9yUpOYXsrriw1vlnXt5eIv0dXxmImNTKN17SeL6+SiTySTYb5RpN75SKyJOKQazJWq/b8tZ
cWSo3cLAMaX16zvkyyuJ8O4Y9DMBwDIlqM+se4jKVdgLbf+s+z3g/F/VElkaP8a9QvrDYZ5WgML/
w6fRYfKu0JQaqhV0/RA7GgjHt7ZdMu541M5amffZcvUqd7hxGlmPdj82zc/a/nXaZeMuWcpUn/WG
anuN7qIzNkwg1FrljwYPArLGPExtGPSvRirZ5YQwIsMDbnf3wJAyPvm5brvWlUcWpp4CJNB9hbyJ
IXN43pc1/8gSW/quGOXnH7Wzv25nM1IsY1HTOLqlNXMzCCulest4Z6uSCFD6wUH09+aggmEfITst
2/eGhRYobo5aC0Tv5qSSPcpZgXwmVFaRYh1TUD8fboC2sNNmIcY43IokNXWveApeATgolVSAcEjU
dcuUsopNmPsdlkenx7nbb+S4Q4CNYkleyNt/JMddt+IWWdFhtoO9uiCP97sHCuHENaIcdA95TtrW
7C9Ht4NiTiwo9rwADfovbrRg9n/5n9iDC0ISaWX1gw+2WzV36nzdxhVcbyzjn+HM7BI07YP+WejL
UowowhBdEZ7gm2bKYAsEoApWf4ZlEzIt0YLKskTFzADWFirftT3yKFShQ5ay982b8YGTVaQ8Kiml
5C6yoFft3Xjke41CCTmqqVhiDR3RzHq9YDqCMGp0w2JaO9luXgH1LeSF0DFPoB235nKCbZWaPiUY
tv+9Ii9IX6Ax8hT5LP4dw4+dt7WaWjltUEiyt79bcbJk1ayDo0g4iOAENEOnBZ+G/JvxJr6gNgVW
p69w20V937oaYSiun6DVAID7sr9GP0HmWyTylNkMT28vFwL1YWFOqSTTH6B7j5mz+PmulWIN9W/L
1PSh9gEz2Lv7DAfm1TOjOkWQjisRYFIDb+eESW4tRnf/Da2BKTJ56tyij6SDzwRb3Ivrf7x6mlQg
avNNcClbpvqIeseDCJq9wtCC5NA/emwKom6jHQlcTufBwE7gdCvKhmeeND0nkSX2rkNMiohEM8Ej
Nt+1N3jV/FS2Nbb6HMk/Yo7HO7HHKx3x1QvQJic3kilvr2o4fdc9zXyb5rpIZmaBn1cv0bQYkrjH
tDfI07SokJMqb4ZfwwL56TdfT3sZxY1v+LZ9jd2kJaXt6X/bGQ0LBTdhyhSNvZH4bMIyyCjCbJb8
pcYRaJk6m7XwXQxdFrRFy2ZM+l8K5mVci6S3FPwfzOEek+3PcAr5O+1WMfa+pQ0MQiLw9ceNKU5E
xz/FSzHgj4PW16IptzgP1J8/dpe6G7JUbzYZGWDBmS1x4Ct2121Di/jZqLU0Za5E7ANlI7au/pNg
9frLe4o55yh3L8e5OZX2NrRdoHFJ1fmd9WVTZq1jZqY5IwpeMC//Q8BD7k6+TrJySBKYW3Enl0Pf
lUJdIZ3CvU1oI3whVuI2WmuhYJl1vPWpLQUBfCA3rLYhumlCeTlg5+AlEKUSuWH/uFyp9rexJBuW
vgYtRIL69tethUh8brNvZ7jYMxssRQc2MlQhRaOcD7EVj3XsbC2e9saX8nGFBlGE6EVwWVUU+bwz
VkQoPMbyyfJSrtd9ToNEoRhnAOM+4s4wS8RRRp6WGS+qbjAy+fEvSUw2uLp1wBX8trzOCGltueLB
jBblwd8UaYu9fHMxFhe4iGHH/R3FuhnE8scKvgkLq3SvIHXxhMYUtKE2UFOTKLAROnp43IkXCO8v
CSJHlhKNDW0McI9QVk0aHtfObsUjETEFkD9biV9f/2hl05bRhxp/8WCHLnjUDLyd88HKqr+0ENl1
LAI8241+oPLELkyVQIilPV932muLeIGpwt/181hgo08cTNWKjlAoznLjRxXEjnSYCTJLjl+Fj8dM
LICjplSK9xu3iW4V8MbbnbDT/7bKGMs/Y39jrnm3WxVvEXPw+iXOUAXY+kNuCggjCiRBEGqrrHY9
xEk27iqSOSzysQYXXM4E+MxGE3aTD8oiR7t6fBfh/dLPr8Osp9qS15kDHzxAOo3wk4FNoRnaM/CV
4bV54O6UPJi8XtizKlgQl/m+6UbdR+3j89/lwutxlWs/jb/dHv67U4BNWCMySlw+KaRYnZ0PjfDb
04P93x/mdv8jbdVg1LflKHzILMzGVBNyBO2Lk5uQqN0i3EYRdztBH3LjZqJ3Gm0Yk/DtBLgSmVCm
EdSASuI5FeWByWRKy5NaEmX7Vv3jECM33sP032HoiR+qMbyU5OMFoGdYfR0hRig063KSirlumy0J
y0cVN8u9osLH/QMWdv65cJENUb1NGCPWUr4kTz5i81TFoFoIL9wKRFzPAyG9X/Vv09RAbZKoXEqY
pZSRL4Vpp/IvAxQ+DcS3ADn+NNokKv4Trcchgh6vZ7LXgf4KkGV5stcCb+6zG+PJEPVs5k0bSpe8
e7lyMY9bxc9c4fE/iu2/7QFVq9hKdIlxTP8kLSVUADzYwQ5OtTJNFUs5YYNR99ObADOYN+MqINMz
ho3/hyzV7uDYf/EdBxYx0VlZka6FXdGZMm50snmP7QqLdWXzgY8Jq0/d6UwoHW+JbHWftGGU8IdA
32Jb6o/BzN/Cfqysy9rReg6SB0s7F6jtyTCny1jguBbXEcSgfSU6XZn9VY7cMUbUeujXFquaOR/S
KPceXaKQvSl3riPZj7uEXVB2aVw9kiuhqH8IkVoz5KS4+HLIJYiDvOiqATqSrN3c/3NYnghIxcEp
LeTr+IlyCqxGCDHf+i4SlvkcH+Yi+7SR7dF9GJl2622MMcfH8U4StV/NoewUKDmCx4huiquYLjJs
E3SN5ctlLbrHH79WDz3udQyCloyc/ozIQ/oUmxsH7fyrmjLNizjteeiKaBA3qnR0YNunGn2389RB
LdE03d0THEqSgGNHwKveC8PxTjxcPlG7/HO2swDdsRNVDNK6ZiTfIlIhtSkpbL51LKnbUfaivk9u
JRz6jmDegm01j7AEwuYP6iMuJsvviGZWruYbtCPH8w+USk4nsm0TPRyVgcFRYLDzzkeWAHBaE766
yx9xUPeAWzUia/opWEkUaGv7PmPv1sYbJEmzWWLBVeoKXVIuj2umdxgpGUO/pjzYRQNdLdcHpznk
2hzCsfVliG34KQJb1ap6f/48u3NhsEj31fPoJJIW/XEVU8/m7vWhpoH1PdaOHZGHuTHl9vS8Z7Aw
x7+Zdt6jQHAJId8xaEgmnmmdxqHUZJtnd5a07GeuYTeedSaXjA/420lWeNL6NIOERxSzgxYY5HHB
KdNvLMcGcN9I6icFV0LyT7c5wh1MKqMMpx+t8SCx+gDTUsPmBTyPINOu2ER1wLE+lGBg6Vghi6xp
O+h2gSFfOhHOYlZMmcvqEvhn+MP3OIgLKIlSAaWJtsdH19idAiOEfTlt0HsWz/Eote/mHewpCdfM
VouoVCEhh1j0QFesJenLaVDixX9S0u2N+NLvXpUH+giK13SavyIi8nmZdV3JWggT5yquFh+DXoNG
KJOFz5m6V4qjT06mwloSznzBP/PZ1TPKniVPqGHSxWvUhPrQT/U+zneGJcTQAM0rDGqPSGGdoJTO
qSCdotDxNH1igEH+U6ApozXaXz2BVNhCYnZHWqGvcch7fYQuSj0ytCnf/n8DLe7sUBJq1o4o0QVh
6TJD3MgmWf4LpQ/p0Cwnc3LhEjFWlkc5ZbkZgaj7ltFDst90g6APgF+DmLMCUB/jP61SpLJz13vV
+IqKIlEdb3oTZtrumlkFZCpAGrr2OABISV27bw1sWFXTL2TTxcJ9ccyYtfgmzpawdmoYNR51LM1d
T8qhMK0ZmN1i8dQNSmFoTUUnQHyNsMKN+CYq6o3KgZDpTsPCayzDImCH2cCpYXXqGa9zJX6u78t2
xWErvfkSq5XyCCvGpWbQYBmBJcMxHAwDEXos0YVsPR58czLxxHtVddulE9YMFyNvfHKd3qi1TelJ
cqVKGlKklFaPpm/l2YLT5pTa/kDa44Kd94x0k4gtBDd9srpjziyck8WvPyt3mNBEOQPsgpnJJsn9
gVdxJgp+5O5tN6vdO9J0rFJJsIt88iEjtacvR5wRYUkUJfT/+7vRFpOi+LzfhCtEDvwJgURiAAIl
IXOGxofDPiULWTrjnIKClAM2zSDKjATHJHchiSpxgI2xB5TOuYBQFZhq+KxPBzIa53mwZ9L2DWWu
i7c2Knl4j6Wav/w1KLctO36U7c+mS9cvECQ1+1qHN0x0VkkS75JHNgCg1fm4eslKVQwpN6jKW1IU
woXJxuW3La9YKA8or//7HL8A5dxE9my7iqitijeOvZgFNajEtgzwtdCUGIfptC4feLC1DoRY7MMj
dg55YMui4+0zG3FpJtOxCVginuWKe9SWHAeC8udR9YP0XRvxwS2DW4oP6lBIGsgb2y1kQsbQHmYn
QtbUngi11c341LRUWMjo4CXG0GiLaEnJql3wwoFLwHuM6QYQL3eVF7n/oyv3Jw/X4H3ofkMbXp4t
/YL2meItFkHN6m728QpFQcRzUbYR/2+wcSOBKJb2ZjlpDQSxu/Y+Cb8xLuS0oZkCC7Q3CqEUiin4
adYUACyAVqvPmBkG/qR/e0329AhEP+KWkJBjiouVfwaOHBZmzloMdzA5iYL9z8YhcBqblQGrtDyV
s/Bhr21Nwdp39qw+ziSVhyo4I9jwvqwHXGRPEOJn3VvWER5ykYTV9NCVhEFMKPcAggIci62Kbhgj
KYN0tfjNVf+n8RApl67y2XAen+KqJ6HOE3QmLOAwgNmUrnJ5IB7mUqKwfAOYPACeVPh36fAhnsiI
WAEZuUymACOdDDiJFciKWvaxTjXf/0+ty8mQLWnKVEVOqMsVnYbir9+mB5Din2+6EleKNyHEYsoW
eYIvb+88x/+j0DX+6ULBK5RJkqJqDIlTuzL+XwSF3LP+cl01Y5Mp0vLeZ5NsCN1b30rp7pJzd25u
fEiVWXqv4vg8++VReGSXMf2TLTYODSYfAcgKoVgaN3Q5jKGChXcctyIgthArhm12f1Vna7e9+wTP
EX1YHV9NPh+5U6tF/VN8WrUF8jBBckqJMdb7IlwKYPWIQLPUkLfuBRLS9VcvaaeUbxfZnvBGz0M6
wpv8D8WeGZXQCxw6heD+a27l7c3UmLhL8akBT/Z0zaYQ1tGAu5DGBlDK4OiZmbArFvR5FtV5TAku
8PhbOXscUH6J7RQ08iVZBRlD1jAs1f74xYS72s3DhLxLoY+RgPJdoEq/y3dlnoLuNqRm+REdeNBC
qWz0NH8bMvA3TL2bokEDXpMxLTDunNwfdLkRrf9FUVuxszqqekXiOCPaXz4YyzUI6vUy4bcsfjr5
cDz7h3auH+HFyp4UG8UKX/K+woCjaGinYcf0ZArC7SJQxOi9j0LgDPRzlzvDXiEiJj/+7337mx19
VTnrNrP1q9CD1yB1FtXiw8HNu9tu+S7X3nDT/Dx1+R/yGQ0TzSWThM48AsgJTpzdb6dq8cSXFoYi
F3dWLon6M0QgIB3DNpm0D7JOQcVumtfjdBdgFtRFtxuNOw3m+VEIjgfYKuB+/eK35RNb65FF0vA1
zqHT1E0Wk6yHXiNGF/luoZxH8x+FVWpYAtC1GI8n/JrQgS6vsjAXrUdVTE1WZMwnhDcj6rUVJCE8
aTe/NjzZ+Qy4zH8Qf0jIaUr/quc7F+bL5dhEWJDwJYb94q6Yg1izdlXMTIQv2YRyn17wHqM5DWBQ
nmbr/Axz7JHigsm+J0sdRFkEImycOZA9Bx7/tEsaC+2GO61x88ciCil4xNOmsRaFJW9ra+YZS71U
uV8nMDhr03JYUb9veQIaW9OImEvgI7OHjlzXudCsRLEqk73QmJBv+m+9optBCWpOPadyjk7fPUzH
MBXqQVheBuUkn6W1HKMohQEZsZQ+llEt73gI/ycpUdh5GZ9ByvtnDzX/ekB9sLjSDRhivrd61c7a
bB/sXYDydmYnpnP/7BIgEI+Ull5S7nR9HkOT5Upzyd7blqJalRVohHCe6g8DZ3h2DEgDdbNkOEve
YfQw924cOYRdoxhAkyPSnlOWUlgwYkioHuXBKfj2lwgFSg2F5XYIOceNiK3AVRvgxCWIuyk8xYDz
5V9C1HNBd2srPp/hGwsurkUuBd8jBtCDceypNe0dxsMkix1FSMhk6qnahkLVcoO8zD/zFKB0H7vv
3GoCX9yXo348vy3rKh/vs4h5wAHu9Ps0319NL58xoxoNo/6ApNt0ZG8DVpy2nTty/J1kac0hFQ08
++3ldKv6oUeBtWS6EAUV/W/phf/V9i6/YyBC3b4Kr5XbcX9nWn1dXanNzLzUzyyngSdMLWnIDyYH
HSaS+VoYn5eEDFAsTOQOfVabalPnRvR5MD5zq65QZAo3cvOajXed8HGevKBNzM8WtG+Ehicf6Qnm
B0UK+uPJzD0bYqsOCaISoHYvd7249+KXEt8LUkslhG1zg8rFduszQoSU9A7EX19U7T81oevN03DG
WUO5jb3wU67KqzZAUT2uWGiB829vepMkqufSahN4b69vSNE28kwMS/Nd10aTYy61xxSmTc3rKMnX
pbfpmgidU40mc7a6sr8VTTs9GoVa39PWDmF24s/TXGgmve+8zDUYpIKoQeja/M537FBObacFlDfM
t15jozbTFpX3/il71HuxIwXvYkquPGhQ6MxJJ6lyoE3IQuPn96Xuyb5HEkwOWCXhfh+CSOicx03y
W1iH6D6/uHkiMI08Iq8CfMGSTJTEF0OmbwoG5zKiDO/oc8mkzfnuUa2NlC1qaTuO+7RC6NW6rKOT
tTqNpescaSOw/tX0b1MXniwipEe+dIG4XDTItyBXN/lyERz4uU0hnH1hs+xQ20UWpkUMaNosG/aI
BoK4p9QF6cFc4y5zho6GH/btwSakjRaaO2EEGyk+PaKIAd9qiD72B7y0mqJnTnRKfRBwVoFWiVTx
LO1y1Hn7m6ZC2aCIscsLWFj9eHUIg0DDWVQ53oZw5jCSbCgboSR/SJNPXnFVUPf17Yr/4mUhZGbB
3/Wl2Z5MxOtXT9JdqamB5BDGwrODHcw2RQ+mq7vfbokRIJNqWc/3PgQsrl4BlCzf5Xb+RVOkBEak
7y5ycu0xsjtuWYg70wbQZt7942Um2ptuxJX6J2k4wBrBu/lH14p3pe1npDdMmzskr/FuagVm57ug
yrq2Ublgn8RgmIdvLkc379iIIavQM1Bknzg0qTvQxkZwUSxafYSuGeGyjTwqJRxhL36JQqL/w3sZ
689xTqVzwG9jlJb4r+XYcIHwOzkhHn00leq02C0pW/R9PQg+ztNpKPJ0E1P1zXv2qggE+e8hvoI1
44gg50MhF38eLFy30AZkapDFRfigEtbent1KK103SUrbHFqpwX7+V9+adOkYjuXlcTQVVb+YQ+kP
JsmffArJrWue3A7IULzWqTw28rTi0SgLLOJ5S+lbOld6+9kS0RQ+kM14v3SEmCkszO7v7kCk2zAg
WnBvQ+7bjPM39M124llE1BHhNs7da+1AAUnlBFt2ZZp68HuEfepBhcECOrK4Hl1fur3lto0WSdXS
QhQWunGQd7sNTHfch3hpmMaVX9cQY6VIGgKc/BvUBZpi+wjFL6tKaA5KpciAt/RvZL1R9EH+J2oz
WkMKaOwX/CSbsfYU9UB1rahX8C89gyjBAMqrFlIYVLsUsdoNbNgwbHj9Y0mlyvD0vWijyAHOhKli
PtZXdCUFyYvioHQr+WwfBrYv/zUUQRHhqnRds+n93IivVpXNxxuBLo+bP051/JfU4cWCE1QJfZnf
iOajPyW2fGmiBIoHYFfmcQqepahNJfzqn6jaElE9F0Kr7gAkQ5APnHMBHb3NsC1j3D07qiSWJ7ms
RjC6FAhB22g2rc/Abs6UH1Vxwm/X+xDMo/7GoFfFUyHDGIQZr7PPS03B0ziRVm/gCi09UtAqtHzH
+3G2ftwo/CU+LS7lCysuf2sz0Of3hjYdrWe7pNHQ4vgJDQsCj+fQCJIoyNLigrFLO/BTbEOMXskz
rHOWZYC+vKS6zfRdxi9iA+pVjo7iU11zpv/ZJtzOiMSQDWh0JAeDfP0+isS9d0LMkwNdf/7/RXVE
qydbB0B9cHFMA2WcEoQGicds4unJywDYJ4YtgCnp2bQ/3LptUpQIFCoDU++seuu30qoaIR1K/YKV
UYpAIntMTLr7NllXBriMnhnj08OjcYePCN3AZ1HZG69ml7ZRoER70F2t8VloEfkCNSK7HkVq2AgZ
yznZlpS+QPuElK9bfSVziGi/c3cyXL+D9+9c0/6vlX2oma1efvXdz0HMROrNiNvzkv61N29WqmSH
A1og92DT+3W5r2BWtykeVkZuFwZAsm9syo4UPQ1XlkHsSATswmxDiZgDTNps3vv5wfa8n4O9Mqlb
kU7xoQYyaSoueHADj2N6s+gUYOkfvccN56ypLzSKNo8PEAUQdxzqaWjDFj+ZAZYSLLvamy/09Ssv
hjrUrJb6+kc5B7pz87O7XQD2cXmUU9cKvoAAk/cABp0hePCZ0tCZLBb2UYc2VUD+xs7xKjj9Kj/G
Z+uoMBQPXYvmZ0XsuUNqJ/0sfYDF1nduZDDgKHGDm5D+n8pfD6l0BplHQ/xWn04GJypEv16ufYbp
1oePdwVLpJNdlsPpsBJ6ccmP7mvNQWd3dzOambL3B5DrW7H5vn/UUQPtlkxnLKgzG1XfrJX7OcWK
NByOqWYoByUgHBDxahcgx8vnmHgAGdaBu44mShxF3MihpMjEfWvT5I8hznpypLxkfhuAb654YxgR
uhcCnw/FtGpwbwMsL7bvVMtOgXb6qh75x1qxp3rxDuAk5EbGOYEIHT8+fIhFdnXkOS2ayCRQchxN
lYm71hHr25jOGeswxzwNomTvqTXkId4BOs1EQYij0fBTociP8lnYmUn1t1EijRQFNs+QFGub+rby
SbFEpj93/acn7nwzGogNcEVXkddlEe+ERipDr0EjqFGmfzUBe+SUGVhIBu2Ojre9X6ZW32dcPVH2
gUhQeQZePt5D4dkicOsisVyRKYPR/uqeRrdhh4LkN8UxPG18Kos/BpG/iX6wtF4zSEP5RU9W8i5R
8+hQ5POk/oFAbO+2rGuK0uJa3L0L1g4ryu9NwxdKEPCtdGboxO/4M9GNM0birCOa2tZ6thQfFDtT
a5xKtC8AgQvUoS2Af/T0ssV3z2zB/ZuVxoNCQbSaTdQAiVrT4yzWk6ux9Cdo8GMx6F9jtRp+xG4M
fNnN3tbzY34Y/JpWNtgXqM4un5+akFokAd353CHNIQVxbH4Vl77LcC+l679GxpNJBFN0dAoPFImp
xsa/w3iF8a3oo939z/EIC404tz1n6QnRKDFdNOap3G56OTQzUUfQCg7UuREbzYin12wGwBmtC14i
r6kLFR2YGE/sL1aQsihgsdnvDnaRmkhOZ2cwEweqM5Znbmk/+xovHn+77wBjGDRvOx27YC9OISGP
k3ot9yYDdJYkklS8D88IH8wHPaE8GU6Qr90NOrjNWYJ9fAANRus86u51OovgAa3PRvQG68d/D7A0
XcuGAR8k4x8CmbKU4MprYrD7Fjq89IEqSl5Op0RN1KHS1sMDw4LnIss7fyBXgFE5d+7xfuK9Xtgq
i9XvQs/4ffa4Z8Fc6BWu3G75gM5N8UrzKPbvZcLrYmHU0meAg8JEfK5K4gT0Vji4edJH659BmsDO
Xm7Ga2KWW+HF7KaGpC4EImrvpezzQUJM4jCdQuwbT/HBHi7/vxsfJT0NkujiaPtP77EUW66cgeZZ
rObS0MwXFbb0Nwrj7CbKkFR8envmnda5uBO2QI42yEWrwxKKDx/QyJxkA9S3sL0524wl3kRXGph3
QwUH6he9GDg2gJ/kAfGxnuxp7L1BZTvUuS/wRMxHsrnnaY1R2lh4zMfUsFGA2QNNpAt8XWHDZ0L5
V9131vFN7YS+eL0zSA6s2pzdoD7uIzfxFmNJLhZPy5LYjgC/SOVDxuRngVm/KzCJlJ+i3HjSy8pM
vrO3W9ulPlgfQ0kmCOpB1BnzTk2Fh0q7yMKnJBeAQpoxhxW7ObBqJ9WXjBxYClD7zWatVDYjTG79
AHuKkNqJe9Kpnyg3IedEiW1pwYmZeqEA8Ok6cgakmx81wHuL6NRWXWZMgO+SHW0Py9Xu9T8pwTG7
NsYWddYlnHj05pMi2gmOot7e6oP+DLZDFPkIjxILr9JZnmIRPs+HMqtjc1AX+Ckx/DB1dS2AFCi4
TmweVrkBN8/91ptqyIfq/AtKh9ZbS3J1aQYUYTyrZH4Lffd7XbMc6W5GUH/mk0txxVhn2pu24NvI
TdWTQnqDtyHHDObUjf+xbcCF4DrMJKw2taMJZW+UC/6kkcFW7TFglS3gBe334exe4GNfm81fr/PR
pv4RQjp1Gytbi7+QiZWqyAywL3iRFo7OKIWQfu2bIH8qQj9sIV4tCzmqAUooMMDw3u7Z14eZVYvv
+X3SYAXWO/Eq4EPmyQQJeJCeScJY+nn+nRiipL+/p2lSITfYRlhr/AbX/BcoMIq8uCGWF/Q3bs0x
eziMe+ovfhnzFSEaTaZ1L2y+rMeDNrQlGh009sQorcU7MbQ7FCHsTC9DoD8xNlrfRzddZdveGFHO
1rGC2vpVBszTl4lJL+0ivzF3LWqGnNsTlfFS7VFWFGkxAmLCrgPUS5lQX8K5qSJQrvZ4FUDgRquL
ziSyMbmbHFfDnkeIVnhqGPTF6VttZwADM3H5wVa4zYLtuEpDEczjpq220CqJDEcz9WFUP9apCOAf
bTfnwndXWNUfh2fqnGOA2ZSvuIYTMcw2EhdMpEA4sciip+ACD2z+Aw250AYkHBFb6lYCn+WqggNv
GqBjmDrwnOpkEm/YtjmewE3v29bkGEzVBeHjj9kxM/UO55WVDN9i7B7ovmUWcN91EArFbbLTgjwZ
27Os3KE/PVIguGcY5miqKgelNJ9pzziu4Nw6h4ueGgbwTkeLIeL9SCBBf4HrEbGvvP/+wbe/ZXng
CBgw9exBx8AtHKlFPmUyPgOazGZ2xgeqbBK52zYNaNrrYhIXIDBGsol9TEU/R3XByr4sZ2vdJeCf
Y460zoey2pYWYexseslY4RgmijaIMhHYCJ8mMle8gt3W2Yr/Yft2mdzrziScVMTmdN7PVgSJgSqr
Hdm69uCT9APfFUXz2n5xt1LswPU2dbPm/DqZM5DNGP8I9AXmKNjAQw5H+0IZoh/VX3oCutNpgQm5
X47llBLML7uR8oW53drR8JXNqW1jFbI8HnBUYMRMlW2VEt2rjkxn1syIMtvEN6T47KZ3kQQtCZBG
qZEOO99a+ECbMRWLQjuQ6WJq/R8zRZ9Z/HHz1htC/tOHjQafntC9YKN3NI3dWsvC061oCCow/rwF
KYiCbtZA4EwU956vDXpiXW71SEJi+KZvKoxBWa2P0dQMziMMf8m4/YYHqQJgCrMLphFaERo9F0GH
weqY0aefqJaNssaAPAorLJfmWeg3H40y4DszxXbadCxHvgSdRcFKjb0980B0zdwXrT+A7f5gBRGD
/Vi5xk6c51Xyc19h3mYnU1bUvmMLZzDZsbsOkCxy48XUPRjOFt2IZE5ifgWsE/E3H+svfJZjUtNK
M/UhICQ7XzwLigyjCo12iLL+QZRvWchpxPim0LF4oEX834eXOKdLOjKJhsBtflNmQXwhwQS3hIr9
Y2qdm1YgIHkj6C7YhDPIJjQXAFpokJltA4mDjNdbi47IhZG8rM45S2ZgfQQQq0KeZZlOk3LbeSdN
mH04sX8H6si2Ep0YbOSRK7LlzNNWW4pB9p8iX9ryU1z85Xg0UOKlCBQM6M3z+z4o8aGsEfre/+lx
CwyWDMFT/d2HCp2V1Is/1skeN5dQaXyWV3f2Ol0e+4reQNGNjTCis8WcOGTIqNhPaqi/14Sgs1nU
19D88FjX6eKyOwFq5L8XO2sJQf6S24IfvLGDIcmUZLgP4njw875YcQZHTOP3uikq4R8qGDVq9PF2
DJrUrtI7xyqazqtiViMBUM1Db13EvZ5YKtEGqj7T/Rat+lLvngXUTmy6U3LqZg9XNfVLwzHCqWd6
io+mMVmiJ0IDA6OMtRIiTYsZ+d1JeLKVhehhGJQ/dJRgWx/cPWwLurtFlOaFAFxHXPnu44pTMcCI
sZP3AlJjrJffZU6kS9mdwUnwQ6oJLChccEiSdUpa8B+L8aDKgKlYLjaGkfCV+RLkTe+j0pFsLHMb
htvSTIxCdOG7N26ALt9vrl1g89Q62IU4bQUGLsVF1Nz6eLfFbd7L/oBqx+62lkwggBwbVeKNF6vU
8xboXnCNQrF6EiMBCEzHQNg9cO4LLHnyS/CLBi6xwXSyBe4mFtRGc+Hu4XO1A0zRgrP80UuE8wfy
jjWxuvWeTpYcxnKcjHR7y2SPrmZ9Sx1hLnb1+kuyVIEUcnmv3sR6XzMnNWExvN4ocDvWvA5fALrT
XzjZEOhYa+rW/dvDAx1bxoS/no4ASKEBrX9FKZwfRcIQys7ZHi2TGzDW6xIWAgqNFsA0/UBsCZWE
4Bvq/7rAaVHpG2rnDzc8od7pjN7w0Kq42lxTlv6KlemutBFZWYJRR2Qne9ACo56qcnc2hhPa+yzJ
ujgeYhgxZtSm5CrrealWMjEmFYhd/T/bGctjxVAjyy3AV8phS6ii/dp1KqKDgt4Lh+aCxT+WYlHn
GIhQbv07r3BEJvHI0wFH2/7HLauY+CMUmfmqAgiQ/ri+11rMLRTmpgm7E2Y7LW+BtTpM3o4Hztqa
Z6PnygsYyf2cRPamwWFH8B8bNl4D4vdmVKANxr2/ocQ68//wVdB7J9rz9x7nJcUuORFOvkGf5YkX
iy3Fi64RV/wTqKc6Q8Z1ZV2EXZiX/bu6sz0R4IRIP+JFz5SNB8H1DZcglnsCACuDc4GpQUM0cfwv
OqPJs2C1u74TSs5mSf1ys5jT7tA6wVcPcXcMe4gfT67oGiAEx5Alyi+lq4Orf1YwQVm3VhOdj5GO
fqXSiPWS31WnMuY+gIXYthE58Zg3pGYeK+BJu0GucbD+stkgISlAH7Ai6zCH15m0xOZEPeBAs8fO
B36cb4AMmB8gWJ+tqC5llH6VDPqmhB2vG+Es2IslNkPQSm1gtmVNs3qriuQ/5YK9rK31iSEqIk1m
82rdGHARz9sDY06109jAug3lu33nL7oG/cqKS7Bfl3+KqSOMoLWUCtG9mdTuttm6VBh+ESNQEkmZ
MH9xV9aeWeP++fCjaU2duk6zDewOLLIcvRAI4xAlLxQwGAr9sRpN3/hN5ws3NR1sjmuua0yUB7Im
CybIyOjypkQDLAxHUzGs+m2c7iYBN1jqBa1uaLd/97UCPqqJRi+27dNcF95SUL9eZkgCEx74k93v
TsSjWvr6xzAIsOeKMwswtVjkBpny4fwuw91ft3IV3XQjiFn4JIeidEqTfv2zLUgZU3QY2xaPhDgE
80t0oJ+6sFA+kaRmYpMnX77ucFqHKxpmkJcHEwcZ1ngF1aRMcmeJMwaH6pGpzAGRzjO8pFSVAzJN
wLYpyYmwywZcl3nlq7zGyp7ZEqPM+bv6c7FG9KTT80Fi7GD9zBmHRrZWvSgiwUCg4la0Y9k8ORCp
rxqEJSPyY0zuIOHsYTJvTgHKTXe6IoPS8o/lmCSrkVed2yEWDr2JrTV877Jx7SQv47aw/L9hB5gR
LrLk9ie3BbSnfLUzoTkjGqgPpFTDSNsVn/eFwEpH2n9mZ1ACJ8rhNa4VWoYbGvI6a/DcAWIPRetG
fdm35Me+uj7hrZ4D1qfAOeWAz+iktaYFaj+rdOrQ36jmfiJMpY36y8VlJsRJ0OyU0MNQNo8ArgPa
tTTuW/0TCyDYLH28bYdDMQMa7CqDSzS09mS9KME1+b/z2qixdGSIf+eNe3ecbFrvMAOd8mi8lVK4
2GLIWLRC+ai853TZSMObnpjuqElD0kboalFjVncdwL+3+sNQehSTAAHP0LLoHHdbeM4gcDmBMrdG
38ywTzu6b6cXQgGYK2g4Ioc9ovU29+ijUds6QBH6jeq48Kn/XJ3fZ+rwgGowL1rxLTcCwoQT+Apw
679e/eG7HpAoW0GM2CKFXBZmPy0MitVUrOcNd75T2v7RqVYnBEzj9wNoyGq9hZXLHLX6pkFE/ywi
zKX5tHBzt0CeOzwJvEtlP5eWhnG2AT3VbcS4JFQuRgcWpiV3KQz5bzpzjo37RvI2rfDOwUgWqKcG
eTfDFpLaiWa1Ihon0IFVOnJ7tTO4OheMEpSIr9SjECVV8oZ7DszIOHnJczvMJchlwWMq3hEj4Dmc
xXg5TS4FJmUO8eWiKOsxGYidM7dn/auUVZo5hIzD+2Xo5FXW69aJ3ojMKJ6n6zuAwhURno3HcTBe
S0NFVMUzezifJs1PxRv7hNJj++WVwwykt3ef/d2pbaWZsTCLbLeUW+BF5itmMFvr3om1JycxCK8K
h19kgDbuiOSKZp3yP1eo3IVTAJULP4Za5XmK80UuCL5wmRTOBqbbb3Tq+EnWZXnEikNgdqUc1rl0
J9tkN3uJB2aI3Wo+Zx/r8HM1HPeeLVzB+mxCEX0hIB3gPcuyH9RlFYtwTKMkRV1oWbVtrxDldLu1
+kQcp/mqV+gr/xSIsUNkWrwVS4KEQA0HbuMwlAkp79WA/J8abAkII4lbmwcuODS0Fd12OOKx0UeO
a4yxoYBeTbxWPGwy4mGZWtVRZXTGdHNr1/hLT9LeNEMLChxYA4byHHRLxBHYKZkdxeXTwdGctMHW
anbZP8qFtjk+Jar8F+fLPRDnGNpR3HwC78o06JXvmL0O+B45K6Ap0y/4QcEMZD5KaPe47hfvu/N7
X2Z03a4OSzVyFlJomPLSmzIhdmQvHUn8bePDeOVjCRN7+EN9VpP6PbRSjU0KMCjJiLyk5kaBH0Gd
YCQUDLcZMccA6iyn3kYs7spF2vYg/zUeR6fvsfhrfVZtbCSUpbx70X84EOH3lpK6yPUe30wRKXbV
4SEj/03SAfIrDR7FcbF3asRARa0occCDcm4QCee62l6HUkBQF/mJyPEAD94o7YxzNhisYfIL5Mb1
u68IvMC6Vm1KykPfqFoAi34+tjLhjUT3+ZzKj3Cabb5GDt8dZTDuxrPCaDwYMg18Yxt/lZKKnnrp
baFjlP/k4dWWuENdKct8IxAct3jdXnZ7capeeKoUIpgEtF5LIlKeVnxUvT5SpjQ5pCJoSSY8MncW
xetFRgI8HvhlItBAoJIwrD1hqM2BanW5shWeoafPX6a4dSZX3DA9gffOz0w4O6m6eDr9nPcynH2K
8XdocIW43a+9cR4YrAYMJkPsWs4gwmnb4+Ccxb1+mSTLDuqZ/gnHP0mjajE9fJDuZvfWuBrIPZ1s
nC+HGFubbC67exSuG17LOgnZF/WliiwYOEhCWhsgQJmiSs7MX1m+qt+jvThh3mG9Zvi8wTm0U01M
5Edw2wEL2V3MKFfjTmgG6i6qxisk3labSo8hVTI05fPXURigwub0bDWr1ij3Frq0PYAkV95rpv5d
pVu9EUipx2qi9KhJJRinIp4u3dbIHKQEDH4LulB3VoHkIU1NI3rrx2yQTFOz8RjGYJ5wzQi1YPjC
bZcs+5Qe0c1JpXLd+mUVAmKrrWoubEmZ1U92PUYePoWtN0xancnws0x6DD1YtZU9uIBfBgKG9ZX+
saTgSFhz5GZ2tmMINCb0vEOTc5RixMDYbKV3/FDqOAYWNJufbEr9knMU3bKBEXGt0uZmhOm3Oe6K
9khuKzVPbOHjnTmLhlYQbwRWOma4fh0bnfr7Fyq4pl0FTFSkJpfOs9xdmUTe4CS0M+MKTTeRNQ0i
DpjPpjuKL4CyfJwQOkS0+QNYI2aSjGsRyEvEoxqxSWq8DMkDFAd2MQzYR7NtSHJUwH7D3gOLqY61
buqnoWbNO6t/V8FWrPxY8AQugIL1qNnKvOJjgrbdrMrB50PWgCDuDBjSoRp53Eknj7SW2RGtmaS/
mQlJAUGQv4bMxvyHbfwvsL7xlz0srnxGWIuTevHISUVq/nPtFpkc2/qv/C39wTSpyoJl+axI6xel
lAZFznseFNfR921LJhaEme8GeGxO9//2kRzp3ZO3ouNCLbh2rageho/MsJm7tonp/9B46k3pZisd
+wlYudEGHzYNsjbcmLgOaxkFiY7Ev2NVlqM1S5WRD546Mur00BRWCH/kYOwxovDxuz8ZDeF9Nm7w
v4Yk6lD2LX3IFOykXQaAQqSb0Ht1GoIECdAFx/OqSwm/U9nbCE+5jDW2VEKZIWfEmhCkowwfPY7H
bh/grrYbx3SxjD0rugxgx8ItijweCljQMzRIRdA4fyzkE1WagGBSR3CeOyVweP4tRiIuFQiymQbG
EpPCkNm1qz9LL19TN6HuuAntN1nWzfrWlFBsmrOk05n1BuBloL9+m9Smn1mg2mll6tOzasQ5fAH7
1sdXOUjaWUEZgcz8+AqXOAu4sen5ZN0dOxNCN93/WQBUo97CZN2b4joHflVOBo31WCDs2lPVK+IS
7Vb7wC2+kQLTy06hD4yq8ArM0csSkwNZwHgJSfghsT64MKQqGA2aLvYJJPqBMMOgJuLq2jMCMdii
051r2z0bl2wxF7q2LhYbVOvNYD1TinKLP3hyg7VBbipG6D+NvkL14+ZBHXuDTgcAIngrH8+lAGya
1Evw5E1EjHMl18iYQRmrLBI7jOGK6SKAXO8JYvVu0hlqlHhgVdD7wR5Vxvq7JkweCjahqtwpN0Qa
IZBvo+fUKXZbKm12HkJWXwVEsM0ekEcfafYoo58h++qggFP3pcMmRNsbRIbJJEy0PpG1twUO/vTL
7MQ0QHEbu4JXxc4HJPZCNhv0mO2pVz/QjM8r1JDg1PDZVGrlDLnJIjhP4gpTLLKS8cKX4fToD7IG
CHfMPbMHG+QiOno1yp4kVRle05Nqqy0yfP6jR0hj4mRsgI7gy9OCdQB25iweBW8ekzpiXXDq/In+
UViuW4yJkCvVqtDzQbyoTU4R17cad2hnRkz2CW9mxao+1aRLRZUuBaF4/8kyyonWLMr9IFW1DBQG
7rtrz3mFQu0Hwq9fNjzcjCI/bphGAoAlDe9Knbe1QUO5cwq/buooV++IaszYjMcbMz+FN1IiZQbQ
OoydaNeTT4cC4ANsQ2s1UHQogt+qOrMhtqTwwRiMV7Pp4GUY7XekBrWYLXTgzuYreJlgQj+vXMdc
b/2/Bt1Y20Jgov8X94vVA8HoCkbBY2HAzKsJ+WDULNs+Du8vl7DNu45F4gmbvp8qZXeIKCjFjpbV
MRm+kznWiTEp/DjdceEpKpTKkEajaGnst2oZdVqnDxmoXc8fkIbXnTSTd4HaXDHO7XtIGJQByr19
cndj1Xp+HC1jRnvFAoOcWi89ik9OxVXNRnW30snGxgeqfxkqdvYnVBHPsmoHuI+HA9fNUcgMz38H
UiozSea6Uk3v8D0kj8MLIAbgNdZUY74DofWqUVcwz2orwri/jil0/HiRuBHRLA1YYiKOjicWiic+
Jn1Qzji0nUUBJKT+vwa80xOkf19iaNQP3A/Z8F/l7iIHkQNSr2spOscxMZ0VM69rMNhB8x7QFPkn
nZuL1QMIUkSGTUqapBI1w10S33XTazcPNvCBUP2tWmNHDDIJlHSHDO1dq9OWyxhCCMmSxDnHig/t
xvV1ybGCYlmjIbChOK5iVFuNoj8eqWHUgTWjMU8fKHHePbNm/qc2+eWDmiq+MDj0d1HXIsGuFTCf
t2FWptQdsvGNsPzT6WpvUesUmemRsXyawp7l5oOfT1Jbed9kn7TA7lXnYVOTpPFBQjFPnf3VV4PG
uguMPpm0w+PTqYa/lCu1l14tg8ygQhy2ZVJt/xW3Mxd5K7gds/+V8Cr6XhL0bwRaewT+6hDu47zl
QgRBVc4Oe0ikrbC3d0qMdTJoPvT+qcZR7XYFvjTYR/zyuo1KIIZGs12kKoLzNURZQfFIzzCeqch5
82sZK6Ep8smQBxtDpQMKlN5m+AXJd3V/lcEvXx+OWPAmNcxQd/uBHCP5C1pLU7VadUBvMbNvb95z
mluI3xWP3prq4BmRNKDMJiGMyGaCNY3mTQxqjR8mvxTE1A5Aw/DVFctq/pYev8eIplhaTQfczpS7
SibNLI98crdq0u4aeKP4loaIBHG0thBIScs5ZoHUFCSBWlmPFm1HkPXr+13sd7RGUQiOoOjZR0cS
lavKpKrXVsp2tUqhMCjfpZ5IcENUv9Vd+h5qRPH7ikveg2knolU8UHJm7I58nrZsu0AZqLCGfsum
FkWz/fhK97GhH5URsjh4b9kISDyU8tFiCehtCr1/ABoOCOjZo9yRaDb0lONUnyUtm0ylNpfpRxVf
NfuKRu710bCVJL2PHK+rUIB5N2pGj0o+07ALu/vYuP4o+DSWftdj9PIXhGdn8nuj3QuXBQlg6BQb
6kgg7u6tpS0WfGSYeXZwTaUw8KRjzOWbb79sEy76W+5+P/zbRrJyAwJXdNrDEoP1+TRIAcgSkAlC
NfFQxESKJenRqIkDHl3gpYGwBGOaSxY9YJaUic3oRs9yAXQpQVYv/6m1Cn61t/Q4LpdVHjzO3oBZ
wTrPi5FXg75GlV1yxUaB2Yizou2R8bHVBQOyo2eeQ5ARglblh24HoExJ/zCxMix4865uhtRkLjPi
2fn/eqILWu/slDFEKf3UQwe4mRlV2tsXBZaetpU/0VGVLV8k8OQw0kARp1ch4S4pYRGF03T6WOmX
G2OwbcS8sLj7+LcSUsLdu0u9vKsz1DwBBAyHVe2qBFR/2iRfpQtZalfNjxQZMJot8LtgQjT1tlrT
fZmTZ96rPm6cWxvUCKJGcHTTMHq0SF7jbRGskFxzVtnvlPEhnMPUaC6/uJMrYqoHYNiTDIU8HFsU
9AOTvbYU5XO7sPoZENKKiQNIg5gCtwZGv1FXqGvF0QnNBakQ1bBTlaM7FiRZKE0NLe0WsQnUGFTk
Lr3q0kcsgh0cGvM2U6YpHczjLC/qM3Z5Uz6ZrLU1VZJc+tYniZXC4gRW9o0/STRfavygNU/jFtW7
bFDVaT8/AJFazxnmYuGLNTidmiBhuckdI543P0sRWQeWQ456KVXqaOmMvHXbJpaLTzhySPSDu24/
Y2r1eNRLRFzLttUhWrkMUolu0DKMV2smxeO0PCO1M8w/P56NunNstndcsS+/rMN1Zi5BB2WyjLj4
jQdAj/rPVZonXx++MXv57yaUdwwaPIIYOkLsi5CsnGrtRyQVcuNgoUt7pcPb4ZJJSkogOPu8MsjN
okPOumofscZ9Bx+joII0KkNnRSxaEgyETun3DrqfS9feszT1gu9w76ceu8PdD0N6eN/T0Kge41db
enGFhVQU42AvwZ1Mpkii0Cy4hAwYQLe1YtiPT5dbVKy/865xow4NdRn5o3Roa8npC0xPwC5KwzVw
sSl/0oWKl6zrQ61TKxXdfGvqVBgL/GQM/j5OwiQQYHvy8HjXJe5/T7uLKEPsL4hpzyggx+K//o9W
T/9uqn+2NX2ncvZN8wh5T962zm5413jgGNbUHTqoJXqEC0n04Ml8x1tcfZX/FyyZXAHbe0ZaTFGd
2RZEkEc1c3hYp3JYMAnYaRSG7Nn2nbnSJP/mZkq3D+9OVRSyRULTpyNB24MfqvLvPEsjzVuiMmjX
Hp6hXEr9Ny9EJfuSAonQBN3H4+oZETddVKF7nNuG7cKS/5Wp77eSQwxef7jipQznXJb/c8ZqT9LL
KhBU9gvl14JOJV9Q8SbmkWHXVlCVfbroW+h92MRIlpu8SSvnqbcaOx9Cpc1sd8WzVyUsf0U/swr9
OVnL1Mp+UXNyZYGdwCU2GBtZXIHUFWUa3xWIpflpqTdnN42fcyHsuBHM9SsLMz72LPylL9Whqc3C
0Chz+cLh6M5j+PHbaJ5NsJcVxXiAXPJFW6A1oi/dbXLu8nWhTSFl38VPyn1m8M4tPJ/uSpBWWlbb
aFqMIMc1ucG6wHCKTmBfZ4YqIAqCVVfXvE77+GJ4Wp0kydkiIxkfC3klAe5pPPDmJCA/9OwxQDBu
0alPIQd77hwJQtisrE6P7EHavsG9LtjyxbnAJiynEGhmczPJM2ugqAwxp7U2ccoQ9cTo7SKy/EER
pJ7Y+jL2c4h2WFnNVXJnzU2aRkQYtK6rkhpQIBAOg+znV5g9qbDBjdQ1N+7t4d1cMwVyqtAhY5Sw
tKrkEWhKdQUx12iJJoeUEL31hojqLk78GAPVTnrM470l5KL85ZNywgNoHGkL1oLtXXDZVIFiuYKg
waFf3cr1BLGv0WdBwEjMT+9bFHFBHAcfFjwtpfloC+avPQbJ/S34H89B9GkfOkyFhD0xgf7AHXYb
S95rsa877fNWMbJCJAc9vilnBfD/TfBHsslWq7Taogq0X6fLABRIzqqCnUQa8X+C+pVNFNH0cxuU
FcEqzOOR+ff4mvSyndtJXOeZQEsL4tI0WnabYj+qtnZ4oIEeZhDEkvCczYF7Zp8XgvS/dgyon054
jzPKL4RBB4LyvIeFejcMGaOzP9AVKNf67Zr3kAz5hJU5SIhohxFSDCQ1OrX+mY/kA5vFvnpq8h6F
kUGwrxw2jK/YqQsy+z/4+dhJXFTFwY0045XFbTicEZNp7YUCPiIvUXYvd8fsTAs+DIQC0GWdPHmz
64E3Z5X1lMsgORn6S0tZ37aqfD3+kYd6G9AIoBhPweeSEdA7j0rm/30FZrvWOtkCOGZYA7y6uyQJ
y2rvTjj0/kGSgmwMoJq5I/z7x0Uli8KZDALAVzoGNaGD1K8nh61X2ZdiKts2p3v8PBwCtl3TxppR
0CcrshUcgRCm+NWwCO7LO3Z9AcZBQBBRupwelwjan/Tyd7JDxbGno7Zm4J1UWA/Yx7dfmEikZKrR
04iSK2UlxCgSvA8jO4EetmSlD6VsNtksgwDzkqX5EG1lL1uYQqpF48NKNO3PPeQuWk96Qm0I+VIC
Va7ExFFM5C6n1I3nMqHbwJqP6LKVpkR61z4LgKxjpfb1H8SQva4p7M1nNVvLzRb5Q5N9MS7KwZ3m
VWT1/v/XduIwCA1QHTRIx10UpHv9gcknN79gei8X0i8riUt37ky3E+HkOxn166xjBAUL5Si0b1Vn
U8Lnt6pUfRcVPO+mvG+akPnrsEwSYZoLwaKvbPrNLdJzQGQVibpXCZpqf6mRt4TAp9Wo1bicN+ti
zq+XWMeB5HYhsNMFxzkkT/Rout4zCv4genvtItDw4Dm0dz7caJenmf+KYHLQuD+d1kE8IaglCZr2
Zm71tNSLcd8HBhtgFTqdchdr7TMhv2zEaleUMPqDONM1CECfjmb4o3Lw7pytInB0zlOWAzVopqQB
BAi/0FpleWRzoa3ko+Y9zd8LrvcXCg+9QSgSHkIGyqG+lgkxcC52rhzje5UFyeLAEB8BiKFqwQIO
94vCsy5t3Ev+EBIZlAmAdDoNOS+D1IOsfV64bZFF39FsfJeJPvXe1+tluWmWeOll1qIWlrlNya5g
MIGBohG6MQOtj7L2YnvnQJ447IMviK93Rar3u6tXPiOyYzBW5zszd+WYYxIu4h8FV28+3w8G/vTv
ZhJ0C57i+zUlc0/LyulINvZCi6bX2cKOfJIVbbJL2FPtzgFELm4dcmSBAw0y26qa+vfhax23uggM
NleF818hScFMGccfHn3qbDCai7b4Kj/Ulay56FU+N0VT728ybEPsMvY1eVo3ZV5JbQbotTmYER54
Hcz9YRQMsVxhk+ZisMZc96QF90EGBqipmWEpskSgOVf1rDkPdY8uhR6AvoN9ZseW/94cumQKrt13
4keCI5SsCv/LGAnqQ3weqLmFXEn15AeI/yvN5sAZuEQ/rP9ogT2z3T3vCDIp1G7ptUbX7ORE1iIV
DJeImkNumcspJCMNCiw9QHQcCN79OVEH/SxE+9sE36AQtmmaBfKD+OqYHjETbHZXdFf0fxkS0U8k
/shFlE+bfTD0G4hft8B6dsfvwWkP+VkJgZ4XnLOGAHYvUgncNHb1CBXlTZ7YTmtM2Rh1Y+3+ETYY
NWXBZMRKdgrzbt9Lt3AoPUbZHaIkjm/34wXLA8qWv5ccvMqwdf4WDUMcUcDKg0CAN3vtMhBQlw+d
BbetY8f0eXqnZNmWSEEURIZqzHPCoL4RGVIbouwEHdrUhrD5FTKOdJSgVwqpv01Y87tKMZB7zh5O
qtXPwPuRq/trD1O9KE2oenQed/cFfY6W22+0d+xqrDT/98fkFyWPPoBTG48HojTmeTAKo751RowL
2rwB3wJCRCm8KzeiNl2DoZZUVy0vwyoWPAqZzJyGtxH3jyZIKi02XoKBqJ+BnEP/tQrOG8rA0iO1
+qB2+i0cC8CCiNIBSBza7DWZFJeEWoplIxBqJLFx/Fs64RrCTlng8nH56jZ/xRxX92ZuuduNjXmX
R2jYdORewq5s+5K9wiJfA2wr7xs2aJAxYGxuU80HbDqjP9w9cDn4azoF9yynavw716zR0fZ5TO9T
i1KCHftV2hecQyhbecoK2PVV/zccfUw5BqWm5lrQaneqZWgWWmZVyGJH6gWw1zeZryKMhG+keaCv
eCzZCyhNt5IcgqxLxYkGlivtQw3vPQzvvCiZ2nVB6q52GRSC65RlKY7+6PkjFwEKVSbECxjCQn9/
3WBDgsYf3/xjrkW+4qxXtHf0KxSdO+JIl8AtVqVv+vp5EbC14dR0hYz2yqdJJY4kS1QAGrPjJe54
ThSeWGdhuRIPY67pQDem02x4dx0TeqcuSDHuGoJpPiH+/BnhaTEcy9852P6/LmAxOdUe7epj1B8X
QXm0TaI4+i58x7O4zFOo2LdmLbDYoAAdGeTWKKvXHg7LLj6cJ7BDL9KgRMpU/MQKu5FAQGSVjSLg
SD/L0kdd0wdlVfxjxtI5BwI1BpOG6Em7+keVFWaBXzU+hiO6TSgQJxAbk4gJB974BASIJtj7QFqd
7xncmo9Zb0j12BTalwnx4dJyqmYxnfaDN1HGvJk3fc2/kEtx9PaqDzM00ARpuQz7gO48kMj08uHH
atweATrtip5xE3upiPqNTJzBeATHT4ULeIV0Vedy8kewGMvswbImxQshkM+A6vgR4xjFD1fFEciu
ls990I+9xIbFQ0bStnOrGK9EG5r5+yoXroYyZyZZqGkb+sq+NLiyMbTNk4v191qon8r2uf4YCqji
ribgAuZ+27q0tTYZIeXX6OtbNZhzM9Tk0sdjhrDhy3R+3tUqoC2G7674R+T61YFYauFPGl/id7nQ
apehOn18gxtV7f26dkBFlgzxM0wjwCFLYVKxzIU5l1ttAqngGn1/7pIeutNBUJFn4AsyPUt1x99W
9vDRZk5joGyEo+8a6FlXRi+Zqp4sR0u5H70GF6uuLv42yoG+f5uN/hIIr7RSakFMkQxYKK3NTFfR
Px7thqrDoFZ/DF1NzgabSiMmMENEuYvpYeJ3s4X0XvfwNFgEIw/IKp6pUnYLEca/t8q+1HMT1+2u
oR9F1M/NMLv7H0dEBZ9JupNciegYL9EeXnoy4V/yAnViOORkfak3RGwqrOouBSK1dksVG8R3JxJi
6aAGx1/ZJ3qw5fpm8uUWhiOBA5sEj8OSIA5ULrtLeysAr3j63fQfv75xpJu03A4iIYToXjfDcVRI
fTTkX6QXj/IPv4c/4Q8t2YIgOvqHJghBEEY4bHBQPJCVPBZiO83uq/MYa/u82nq/JeQbJAmWA5a8
2Rv6z9pCI0g+YRBvWqG47QBU6Wzuu5EdFjLqAeMyK+NBHPgXSS26SpMCYz1RkpGHRBHWK8enjbve
/upuUnalEg/Td6lwYnNOn0/3qDQY4PDeW01RmM+QhSHHCJi8SmAGPBi0uriI01nlaf9eZ0AoWvP9
aobGrNESI2PMTO5JopR6CiHHVLRwjdSpiTKDkBKbY5+FDgFTkJnYdlRbJz9etC0N+L+w0T3lI0gn
iSVHGyPqhqFhAn84QNavez7jj/xcgTYnS1alF87wALXJArZHMqFPTxrQ7/EiZm0ZBpHYmMNSBTI7
3m9UqRbsAI/Lg8n1oxh57OWTbNzRt/yLUoBnsCuPtCer1UMHhfXLESBvWY585acfkUmzu+XIRdSg
nlFgkh46XDzGlUNtvFsNq5PSZUMAejaJHdSvCVvpmYDM/qfpZFNE8rm3rvIH785D7jDHbAwbf4A2
JSbz/enuH8UHxXs1qDzLZuVu8l273pYay12P3jwFP8bErtgaVhBv/P1g6R6P1fsJuSd1p9WCKS/T
7G48UoW6Uyhe07ypVpSkyBhiZ6p70HWkUP8KrF3MupIfRNaH2b5Q6ffwerUoHZSMTOkF4h87K9U1
tWhhpd/zvvjjYn/2yGnCIiMdMVHPffCaGyLnpHmlwryIt+VgZL79ciYGPg9kVBf6n11yJMH/pwpg
98WG0AqeWWiGqOMQdCkKJSCFTdYIomatcac+LWaqOIfoqsWxxpkpS+ldRKcnXD8L3SiEW2J21QJT
CC0VguBREkeQc7UoFPbQHz5KlwXz1pJm/q2aQocYQgpwqbMoweMSJIfadu/CXS6e7RdDceuio4+I
ru/SozgJWjh3R0/+yQ2KaIYYUHGfI8mLmN8h9w3WhMHNu3t9d1aFqxrY4QPS4JoROYx4aWJ9nsvb
VdmJ9X8Jicel//xyL9MDEO3taoFWIpG1Fm/kSCtAIlzHNoFkxmh20ydg/3q8TNf5FvFpX65d85uL
yOOUK8vXSQkIRogjaOkmiSnqT3BRqMC10mWogUkv6EuUObR2MPGd0J8GjboCUNSJZ2f8ZgsYWhhJ
B567bi4++WjxS5Em49LMODHbTD94C5L6SY2jCadIm4OcRIJx3qxTp1OXoznPa0qUTNm9IILOwM22
+IAg5laVy4c93a6zRGkVtFqpUrn1nqqC0MybkoFLtuQ0ExkxMXrVDMwkJSnukzB8DTjo1JPOvB3O
SfI5xL3qSbqsAqDZq9WaleQHxAMB2elf3Xsf2N70uhBIES1KIbLTXqGJZQrNsEu6Hqt170rPHt0S
pkgbjj+/eFFHKcnk8epyLy06YEOkoGCpM0Fovvn3cSJbrRo/0IJcNIp32xcs03d0Os/IkrYKGOIw
vT0Kd31+em5BC4OTlyc3HyBW1vRE6gce7771X0xF8NYD5RSvlStUQoXLB/C/mbo3JIH3X+dFANo5
AR/PYcxosv82hOGYrsC8MYyRW7o/xbL/uXVFxN67YqdovTGxXZKT8xqNd4vjdecLWhCbQVboAL0u
I1LRqP/g7vfDCRCFSc2K8s4vi9pZ6vkg/sgWiA6AFl6Okj38HcyYrINOZmpTZFjKHGkheMVt75kc
VD6NWesa3L7c0Hi1sBTP4EduT6vqgdL290ETA7Sam0DtlBPkaAz6oyM8jLjUAFosKLkjlS3evr3b
mCof5SolhXZ2dAcqeS6t9nl0pUfqPbGNUmsyBRIyj4rLWx2wKLUkVqy3qWgwJzQnUnDmay1NRwKi
vJz1oe5Xl7HZ514wq8oiFPCh07NWqkreZncr8LF/DVwR1yIGBluULVlba4U8puZ0YM8MzMFJKQE6
kOpCcc6xedoPDsff/aI0Gk//miKLzqt7VGRn9hxa8++yy7HFmYRR7nVOhE3O+8cVfm4QSfrhU/78
L5KY8+8AbKV3X7nUTJJBdstHhmmUuzIVR8bxBWP4x7Jqmi19vC0gqOgXxhwLH/9/zb1Xay2x5Pdy
ODKSsi2/2tgs+krW8BY+DuThtMOFqSYdH8QmWt7ybkWdPujUdYswnllST6MIG/JpVHWqjdskhXby
o/WF8lZnl3hrcscgPhO5PdLkTBSzdaNgg+ODAsQlqiv+xNMFpj8rdjtnsfQTaXikeBHQrGvlTGs7
0wCv+kV/bG2cNo6UEP4TCRbv8bNkXfE3Tc8gt/zXxVFV6+dnFrH2+JXef9lHp/EOau/h0R1yzFlZ
WppDEqpwrZraJpGBCPuIvSa+xHk1SERI9wDq65m4jxJ5aYEHqUfSkYwu7hH9V26oMXitdct479r+
27iH1hSyMLwgTe7XVzonkKvIA5i9uT8/cGGym63kIesBgIIPtlc9qZFCEfVjdavZNASdSpGDMLRV
kDi0sh7KwbxqcJqlz/xyWi1Lcofdj+0OJ/Sz9wBzggXgM4uTVAN/Rx7Wv59Fy4wcy1TII97hDBlX
ZluwK0QHqilTvQFFrJeeD0QZLaB/9Xwkof4hhoZPF8JgMc4tHI/A3yMCsTUJPYSRdVCwK7GVZIZN
DG3NFPv2aiJz0TNf7/liFMo4v5PXOcU1fERt+BVz9VCeIUjRrQAsUSfS7psG7DKMbusw/GkZB3nj
rFXtmwBgbMMoA+BPjtI92yPAVvcqGXeV+X8f6ZBM/PULud+pZZHw2RiR9GuL1p+2cou1m35NE5sn
+xIvxIBiRngdDnWUe/LirDVpKXPNCPYbszJNV/hEMVjxV/5U+/95+sIkaYlUudvI1skheAQ3gELm
E0seoJ9pZkFaTmvzyx7W+RYvWDKkrcNSFkC6784wGVzu9KNh7JiEbPadyNx4w8HCaQyAml+BUBGg
Z7cm45C7Cbaog5QwaNzVf2gKvAxxmrGyavdrkULZkEsHbtAU9FDP0Pf2ZmyW3N6WExnjPk/D9JRf
xVwmr2jCrifZWwdVdOGC8hBe6rHq8dfwziNiJCZ0fY1FEoY146HpuzvQttHtaDgETGGqjKoiqln+
/hzW6Gs95fUwUoQQYWNjhNnvUTzpynx/ZB5K6thMnwyq1yvnDP6PN88DQ6jWq97+MH1Ejm7KYQQe
RAmylv4L25QGFrglBb4vQ9GflJ+ccyFjhNITAogr+XLlIsvta5XNbl+GK3Ifmkw+o82ChQ0BGAzh
g/72Rb0Te/V5VJqMC/X4vv0flIN0iHqv5HWs4+w41hjvcLKsJaFlTHPMvjB8m9I9DhbB2/jUJDmA
QH5IikXMJZLmTD7fnx94Nq8QjAxhNM0ULXj5y5V+ylIiTDYVBTC4jKgiuRJZmwwzaw0ZMLiPYoQC
ky8j7gH0Rb2Ih7D9DDMLdegBgYhJbsG3307ACj4pvaqGIePqrONZfUHNiNnEwygCuUrAsi+Tbo+0
+FMD+IQ+O4AA5vH5NJHa2tnFR6D9yuikBEY2/KrzkOOxDJHB88KbTU/irWeSc7fLzoM3dmkkI3VF
ISbTu87bAUJwgHsDE2dieSeshuRcS+oFrPfCmDzd1zn1S7LgUghzNKg97TZsYWd2Sg2qP+lGCLTJ
SOckdreQyiCql6OBcpUF/pP409PQETuZWmmYO8UpFhx5eVJ4caAmxM4RfyHGtOmxFe8p9JvDeXM6
KUrJEm7V4FgEquVWkAQq7zxggwwBf51y9AlrGmUOpW4Z6a4Fwv/Jbv+P3HoJTEmB+itSPZO3f1ue
NogcFszT/oa2pgRbGOhNsasXx0N2o0D1QV+DD9YuIyE2BTVtrkpiTUSMVimH/jH+qOUSgocVQsfg
FcrqNbgmfrEuenqzp9/Ya0jT0FzL+6GiokCqqAAZKt2MQm+BWpT/ZEFmP2MZt+wWvz/BtPdDED02
GHVIH9iFua2lom9fpqksvcmgIm/o7tAmfG2P9/AmLbPyp/YmNJqVJwKZ8eIQOdGkJhN/u/4OCmdg
0nzCDDrhfd/ls6dsspzxyr3hjRNll30WTCJPqbdULgqpXJkh4Yt0e4rcJK5KJPF8WzTu6kBsxHKo
d8qiUiuvyaCA+gDVwsBGYRwYtPg5yTYKalC8NX+fJJeR8dV/XpPPrT8AQ/gidW3KNkYa3jAL1hrL
m19w61l8K00PceCvO2MnDeMvzJkXbiMbCrhFXIo3Ql9BZgq2fcLF12SEv6dtkGnGRuE5Xcky245M
NTmHujWn00jOSSXw1J2j7IiucS91mhWFzT3wg7khAmM3GRYIgibszW6Hr9Kl6hMX2IH9jMXo7DPX
eUh3Jlx0Mx/Hm1yXcvgOUEin4esNokAWlTG0F9Ba3FctPzaYhyImGe+1tBihUxRPa7uqxJZYI/T0
fz/uq2BR//+7ZoqczJGwpvO2sjBXQCAXsvuDftvKhjQ4cL4QQ7n6wszixHBt+Sty0dWzUz2aq47f
FGM8fVmh8QeW6pDdBu0kWJfRRGqOXXuM2UKt5infrk9WKp6UT+TXr8cgHobSJpeoHgFMQsEC3OA/
JpuSuLiRJ7pREF2HT6QH/IU9TqghsnnLuV/0LbStCWGySTpm0v+wXzUpAhI+7lKBc5xgT1HjpanB
yBaWfmpjBra27Jbg5YL620B44yx0AtjOXny+0Mlc+0Kfqttiw6vI6T8v5i6+qeozHb2Z6zng9+pc
qGXKgLhBs3eoFCjuI4Sc6UGLqFGvr3bZFLxx8+TG5Qj46rkfqgvQ43Etuc1zvul42x/Q0fznyox1
vfappbdQgaqi0+K4MvCWaJRWp7IEiSS30IvkFRxReLWA3Kv+GoZjCAWSqy0Dl3YjF0nLzYCEM2Cg
g3yjCpAe3OVpXfg6pnq41k+hvxhjzPo1HmTowfH8+CGII+XM7qfptrOYJwWuEaoEDLBWBjZCSvAS
P8p6yjfPCeZfubK2u+PMyIuAFZvWqA0J3Z+D2Bipz7mkvdiYYNLwN5YUxLucUxSU5va2FZafhArM
THOxk6Oh0R4da3mQX8Li20U2xSPyBXuzvJBHSgf0C5amGV8x2CpYdj50no4Fq0et4KV4Yra2lFZD
ITfOU4KE291ZVy4hYD/Pgvigo30O9jdgrxj4lt2lDbXUvC6/+5yJd7cCPw/DL9+kzVhG5ncifasN
kuJZKAH4SyUMoFQHWt5v7occTUS66BMG10E9qqEyuraxT8UMQ7enGkgQcs+CYYeDsIus5MW/cHVh
1je/0qjSVXbnMJwhot9B6pN3LMHQ2PdRMY6CByIcp4OPC6pE/O8eK7R6a/EnlNebwSB9yBX5jNf5
1zEXLFsmCRaZyE/6C/5c1YhKqvTfnLkHmn4iNCRPqeEca1CQXts5r8i9HSgeKFY1ei6okswQPx93
FhqTXaXBlmA4J9t3ODERY6zTkqUYYUSHuceFFhYpemMfMYh3TX7efGNPhWa9P7KDdnapyhdCLCvk
VNDLvd4ZOboXdHCwlVNEAu/0CiGpjmdKT4SsxJjoWN2oD5e5/HHMYA487OLpeFvlXXRMcvHAnpw7
whw/KWnKWmG/oEsTagTcXIJuhNP1q7T57MiXTSo27hWW2t8YhppNjZVNIi+yM2m+OvK6p84Gt8VX
Nb8VFgdflDJaIrJ+H6nG+k/fYgo7skcvNiK2bxQ/m9NooVaZjJwyKRTEI9ubERog6gnCAX4u124h
Gb3anRuBN+YgLRbX7FhEOQE76LkIJA0g1PU1LSP9iwd13N7k1JCc23CTPBOJD4x3Q1aZa1e5b4B+
g7BpOFIa0sAEn6Gpq1W/Q3wS2v4kMdK4uyXLsEMTl6aJukLp5i6CSMgj4WQWV5McRLhj2s/UdJKY
nXDgG93/UctfHc4TI5lBvUzfaQasERy2ku248aLswGFzjVO5kR6LBcQYXxxCKocpdsiggqPGHJnp
uXKsDjufprHldN4ijXVvsWWsO+eKLIZ3oXPRdc5J8tqXbWBaMcM5pnra9aRJh5tcSRAKo4CfOl0C
aVwTRlFp/PPmUruuaTDwQrsiKJiEBFB2wUyrCTjtFwpZh2PZu7L/euts8U2dbNKsWxIp7ih6TMvB
eC7n68/X+J4HF34bUAjk9ckmJIdyp3QFl7tcBGT+GzDajcHu0Q+GdcqgfMcSffEw3ixNt03A7jhb
ai0y2Drb2p9lD4cf8ZxCqDvChFn6kJ5AHc6ccZtotGFS1HQ0LXwFLVMXJebY9Y1AU9W00C2/KBKE
dWPBtKwjFLjGTOyDJg2zJ368Vd0WFnamcvZzumPqdiIKdVFW+rgSzvwacQkUx770JdUGeViF7u7T
/eC194M4KdA8W3W4GfVSJ171SQj7suoAQo0PtUoK1g7rW8ldNpW28MWX0S49scVB7O98AcyYmJz2
v2mheeTpEdEgO+h7HYXLe+pY7dEqLdGqpk2Njh5Yvvnyc9k6ZXCdmCRTYBKeiMxyC01Nrva4aJMH
vnXqsXLtGo8AlAYIk4EfCyLSI/Zev//yzdVLeSqoudcLnKrzMjszwihUWShrQ14OQzIb9Xxl341/
EjHNidaN+H01zz8+rDZtM0ETELNRgIKaOZsHgUUgRXS6rOTSpnAlkFuS2tXFljc8yJt/5UycCkx7
wKRUl/F7MmzB3wUPvvkYDmQeue3UsXGmQZc89yaZsZE3Fnk6KcIJ4GuzKjz6MSNVf4W9sydiSSG9
KwdmX5FPMCVbltXdp9j/+baxD0g5Tu5bTzrLlWDrK9iaqBtovvqHTbDUuQ69wFuN7mk72PTNJWvX
Nbsmg9p4AqUiaeSn963lxkmW40L+hoFfav4p3I0JGV3Zwd4SrieWK3rfT+G+W45I/72u1lul8wFe
JflgqbGNcCMPRD+1DGUR2p5eBk9x/TIQPo7a1En8cfrNq3lfRKGp1GiQBaovpFt8dzBhrstPLLXL
ILTl4a2Wyj7yS2/+tzdeDIxnBb4C64VSOtKxnUf/ij0QC01y6eGC7hQlohTlif44GtMl76H1t9bL
T4adK/FaQj3Hr4UWhZIeTRGeGvFnxIIUO40hA60op8hR5ckVdjErIWKre9fNruS+RqQfscH6i/mm
OAYYKNtLmvcrK2dl2kYSz4v525yLTFYMGtpVfS5MTIT9Sw4XuHE3bphmdNIp/9Ox7dqTg8tnVmZR
j3FhIqpkmwlxyFRorBNhjO8R28YvZEq9JKMKROovYaYa8l28bugyhmMys2F4ZWdVb2oC1mycI7ko
S64fftjyR8piWRzWtTvmh5Su1YdzZdzlzckzvfT33dn+p1GSHzPreSpIQePnZhXKxTlV9hPcX5Os
FXBQhs5xTkPjk1RkCZ3rMintZ0czPLRmWmUjwcECeE2y1lIvF74T6IdHRCx0HCFDF3fPFi0HdDCj
Fekd1TSBXvANHdNCtVEQWCNYKLKALmseEKPoQsJRXhow0qRaENzdpKXNBHuwCtyOMj65wD5Gs2uZ
ee56WGFL0KRO8ze0oLFBE+dPrmGCbsaE4yiHjUkMOTKVehbhuekhwHB70MIxAlfLWYH4HaXd8f5Y
FCGIHu3/VdtNhlePNbWIoXPHu9lN6nQibruidPOec5UQn+fMnE23hXCV8aAAJZT8hHqDyXDoM0rz
N0+LX98uv4gUxgEHBGtdILmHf9k/vq/0fIuVFvYwN1NEcY1mkOfdXI+vXh4/6MJhDMuXDgPtfJWE
H0J8vB65hlWduJIsa8Rnz640kyi8ZW9AQ9NCN9l/nkeB6AZVUeipRnnkZy+kFj++zuFunErjvcEk
3VkPTVdcLFy35cnlHrmSqu6TCexaFdtdRL6gHk6SGQ5yRuayLBxoddexEPH1V3SCuxEwemPguLC7
51Iw1dO7sE2mccFxvBVq+xFqi0BLK4Oo80KIrIlFjw3pv/jXspDfVyY9iv2HiqPutr7hBMG2h8/l
7j1Gwy5BxOhHmQx3Z5q3QbS2NhZxFiIDtbaEHmcsoIO9JUMqGt/H7uYB/it2IonfsDvlq+TL+tUH
LYHS8wjahiW6QlDQ7pGbvh1xX6etIcbMNpoeLqlqFqtwlW8gSRWu17jYhk39xyvy75qRrmxT9eIh
mrbOg3xbcqRLPoJdfGnqIWzSqMDrzA0+T3pobd1WVUlqgSOkrAr3xjWf8oVuSu2jHDSHazUuBu8i
zRnEjVzIhp9hSC2GiwyVaZXcw2acbtIAscPbGQbNH8lL8YOFEQLQ2ulBHaBLHAox2Xd9USueG9VZ
i/lC3j0HAjP072l8tJ/UF/ZOTnBTpJhnhS9G3ClfYCayGljZeWKCvXvUaU6zQvdFYsW4k+UnmQy7
WPupnVfQJJ2RI8L9BAeCCrJnJLsd4GAe5olN/3yYjFQrMb4EgiwXO/rFi46p6cCwKKlD/gyeju6S
bMEZBfPgTNx/O0BLQf54jRhVwQ9yKN73HyOeVfrOa1XyJbSKGhBnvk7uY/0dyUPs6nUyWuALp49u
aXGz7Ph3tSEGF2P7KMkaAKWt/rYvb1XEifXOoAmKeeo8VQjjuR3OnZh7bFmdfPfVRC7nRkE+6cM0
TQfPByKe1VhOxfahietkWq49Smlw15oI081UY2ucM+iiimJR9YYKv5oMF6IflB3oGhOCLh0sLoZ5
ZGF0F5chHWd3PHiHhu7aU7xtGAweo2uYqcj4+TNGshr4uuqfCB4RhKzVX1TAbvV2nEdLzbbkuuMT
4Of881HB1BhZkLKDna3LbmuaQu8jM4hAgTa7/istNOtgB1YjhJPFBOOv2TykdhmicVckyj7Xhgzm
tZ29ghE6dU+hFyK4R0FuLgCs8GBfX/LGLWEMks2SozjpkfvXmft7AobAwsN4qAz2hhAhIGt0RfSv
BssX9ow8AeIvtgXv60NWUoOi9O/IsqX1Ju7ieZIgHmoU+JQJFhNWsg37lq9FMCD0C7QYT2WMGlCG
OLY3c0qcdQAJ5zcYu1n1MyYf6lQalxjowJl4VbGNiDN/kh16gcugrPoXgNTnWq6Y6IU6W5pQglVq
W7E530LlW3wCQNEjEdPydYgk7M38gIEVuVN6S2FIGN8O6bGMlXrzv1EHyVY9FiegLFGrkr5IZsmP
8n5/YRIlGi9TTMut8wXw5S9RnP8yiW+rWbc5HujPVw5/Xt5SEyAXIDEGf2Kuc3f+KMh0BJo2ifQi
n+d23sGFwMQWPFcKcCd7PpZawkohGX0umWJ2jWnRvz7Rjtet+C5oRupg+r32c6TDSuLN8WUJ8Tkr
Lg3bKOg9tNS37zSCOvy1l4yBNF6KaEKXKSZPCLVmie+UTYkyn5HMEqwjumiMXNWWp727DUMlCeZZ
Vhu5He5aPBVkEMj1cJk39cfw/GrWGrob9nJYMd4ghSpi3ulcZ3GdRaa8gB/x/d8XUZCWgzcOmhPb
0v7duWqNxnTLU02XFsH8xoCJEsA5OMycfdOZ3kOMxBrAkDaMm9CGBLflDcuifjrk8p0qwsampPq6
ngIdEMRJbfvCDNWxUzIiffLXgWx1dDi+5wBPl1JlXMfRcP/dPZlVtVhK9WUPE5jH0LioYfVNqsIE
eO0p18ht8iyOvD02aDacXLzbYaHa/zu8oi+yqEAvt+frs6jsX0urSAYDmw5sgWaaNb1Rw5ebpJyO
Ri09QgF/h+DGAoylSZg1WLPbyg+0bxoO+QnyFJoSZQujH482bJUtLNMgrFcfueVtFzwnnMhuHwB2
MaAgQrmxcvgAxnTrf+a9FEs7hvEYmbIXWe7z3zFQ0Id5lML54ClT8AUbWMfwlkfTDEinEJ64a48V
Be9lnq6kgioiU9nogka4cX4+fMLAU0jSWtXFOITXNrzzfcFRh/0gtCPMLQ42/E8n1aIB5Mqh4czI
adHlFXdTwAe0V18jiwQGlY/2W2lyJKuebK7YX7KHa4DI94cPWhhXbYvn1AovgnxB3pryuQdQoYMz
Y24SR9IIqwQP/E/r1MM7o5thcuYs5e22DmRd+7srdB7v+NaMBhEK+BKahgmojVIsexhRcD3Qp1bF
vhcWH+doCQ09ZWNRLfY7gigBeSp4zdGuO61orMF1Kt4vt0m6er5XUEDU11GnHM8VXrilv5q9yPzp
5lFjuIqu/RH5r5TNNv2mvl4HPNSWo2mzNIb/ChluHYfYw5Bp8sCqKGvtHC3gfpyNKDwmuf4PgSH9
aTv27V7F9uDNrsSk53q0RXZ0VAO2Pq1JhKIchh8POjz6v8t6Go7wdQDlape1ic9iWaERSy1jbQZ0
6J132lO6zoQ8PDhwjIH3V1wSpVW9pwmnuSdt9Q5bT6Cbp5l3fd4ihzVAWIMtHhwZxbrmQHsOqsrb
PMbS2KGxNuaXguFIpT+Na6iUdQEt6YHil9GYjnXzbZI9NDLVNRzzsoCYcvEsIgIbcSwviU/pjFte
V2nikqsX49wKzbK/YaTGYa819RXA2bzSEituSjRZvOoPsrXv24e7gRjMdF6HDo41K1ROX+3zDBFe
lnUhK17ib2NL9Q6TVnAwQYPVnDItPy7XN72gXFsQs2Us0PLw7rRlGs8f3KrNoAHJ6VI+DibzZ+fi
sh0dv8n5u9h8Ys8BLRvmWIhbow6Wvbk4yfwAdqwM0O+OzMI0Rto7mSgK5pwN/OUNcT2KZG2maRHN
iFl7DAtfS/M+x+Jsc9WX1XFM5qzf1+XCxLwlt/xPgaZ+krZEceOnRd19KmpAzi1c9PntIZ7wUL3x
WxYyPd6yIhUla96ssjjzJ/tlQWqOBG46b7KQpPVYi+nxVlnUUxmCDpcpKBGz0P4eFDy/+ZnIVLb/
KpIy+kR61yhSQcCW9S24ght2S8m+ODLZEbcyN2fzrnv/Xw1YfQBuSCWF9li//CYoJJ0OWkT+eNKW
vDYpBYfGkLokc5sVrEIQkWPrPgZNh8miOfCBT25etdUmrg4400ru8WfQvIRaj1WKvXywfCJDVaXD
xs51nV0WwuosR/MQxg4qY/l4V1ok62NCr8E6U/7x65GKkqzQvUdb1zJXR+2Wi63vSnZIuWWLWLAy
k72p6wBFKB+76Mg04996YUhbSEp76PazRooNndItt6958yz1PjtvdGfhnywrUl79MFM0erBPnUYd
KxaqQfiITk46fgq6nmpsaohl6yAYy6gfneuI4UhiS1JQm9nQY+qkSGWnc4TK1vHK1rbO+0WszMqm
Hp1bnDNvfKVGyCJFCN9TL5/NB/4Gt8FUsU32/5blePZ9YO3Y+2kFaTfU0dIxL3+CH0Y9vc72NaL9
UyHh7Kygrk/GS2c60NeatnfYpBdrMZ3XZfIh89Zet78Q6/HZS3Vn6UEIyqWR2wExFOjXX7heAIyG
mc4ski3T0TFWU8PDY7gayxxu4m1qoxOfUeBG1NxOMdqr5YGvzqw0T9rxAhbyKMabKZZc9sYAEuNx
KvLM6h8hWTuA5S/x9gg1oOufC8K9DZFlObDCarD0QbbZ42qXE56IB7s800AC6hg68Ow7/gan/djw
GjlscX+4TBdX3EF7niN2nTZFbary/afNY3zp1W1A9p818wpUOtYAO3Ifyy+kTmVL/u8w384YheLw
1CWjV8zD0qUOEilcUARJS5EKucoXGqJ97wHHqNATNGAAqzDJWD6HuFSFZvdSnM+wKYHEUvxfDECF
vyTTowLCnAVcG8b1UDbwddihvecOw/ZXRAHD9hKvOEYOdbdU3j9LSy7bQjQsD5dMxyKQYY5Pfrib
uR9DRZ24OSAewVM8L058jnIb4bBgVD4MMdcNi8pi5DVgMOAvJoxvMko5k/h6IugkZLWSTEftVRqR
HRteyFXPjo6/OpRn5u9Ckwlpv5pc9xz3tp32N+ZxhMse2l1pFp5dDQNLAIO5FPS8ood7IQ2pVJvV
pxy5GlS4OBSGxFvae1UvtJz7Km8238sEHeW229GdRk2cdXdmSdECrjK8iFmxZO0VsxbashNPMVpO
DlTV3dc9GFy9Fnr6skHV3q3jnpHwU1P5mIs+fne4y7owZS+ZCZcuoJGREMssPAwNUeNX+eQtS63G
cYIXCJWr3EIYjgyGUegQIvEyNal4Yi8AbeG9QqWlpqUwcjBX8ir0WAPiK3hvSufDH8y9bm9zpsb5
UZ3hxZRb9Rss7vBAdlNiINh1nMlLpV6oM7wg/twYXYj1ghrHG7htEbePtQ8fpbtIoepyKKl+IGkP
tIIz+OMA11kNNzwIDqZRvGSI5OWAQimMkUuyyqsmO8vz9V7uPf1PyupQq+vy2fBTnJ7dWlO888W7
sjsSiVxby259Tf22ziZnXcVI19Sg1Jro5ebSeCVls53B8IMY3IGXUoVrqpdgpGWJmhX7At67wkEx
w8kQ0YwI9UXipQYOSD1b1SWl+WBklEmA25Qb9BTitISgnClUGvDWsFSIu2ap2geLTWQh88o+3rDg
yq/KSXb7u45XZm9W7W0GoASpfdGQA/GG+EGiGRDdOSnopVuboBRFNA8/f/oN4nxWI06Qlt5u/L4h
SasiDjXOoZVi98SGUsZinJML0HktMFcGgT61IxbMxj/YaFIT0/aKH/ZwDb038jqWthgtRVMP6Cgq
nASX/fqHMEYK6j+vDMsFLa/7bmkA8gyDqksf/JFrRBzn1jVsVdb2hiuqHzK2DKUMQMV3EYPnwplf
1zKsymjNnxNMVdb2R5mAiWkF/ywx8ChltIAmQCtYdFbgKtoDkcfIXzZRV4yROUUyyTcHmUfaBQyY
J2xD3JlNIDHDMieoM3SF5HeAJigf8zuAsL8Lf+XKRNCGEDbbWNQSgPquO+snZsbmSDqDWIeap03M
O21tM31ogSm2JTZ9JuItPlHhBDG9YLeZCBxRiSVcg/UE7vaOznC8jn0x8CLiccRFQ2185u+2TzKA
C3w5CFWVuu0fOQwDFWnSF/jArtr9RvzJ5LRmdQ+s62DAfYY0jks53auamWPnpKYJWf6r/SYiAGEe
/07BrMe8MQdJ8ezuFS4ubK8al3Fc9yV51N8G6x/OrfFhT/JqXaIUmJa3QJ0zuCwmLYLrUU0TtoL7
0+vUGDee4vaguhsq0SSDf91jsqmJJ/GN2/ijuSxOhA8TC6bZeQ5lG+MEiKFFMXUILJCdi6aNSiBc
s9rFydzJKc3C79FAa6LvCsiTpSgs1MEBGsubhlP1rTfPhSYkLvYfcJSBLIl3XSYf17124LEWRc5z
T9MA1X1/3l+qgtrJb7IMaTzf2ti+OD/gXrEgcipoWe/fx47RKfE2y7DICgoXeMV49MJrIOYYNzS6
tbh5yYJyD6Zuc/rBCq3guXfE4U4OiqRv583yVHuZFR2ysZal3H7h7vlymLVr5MLSOEbj4TMQH6Fj
rWXKLX2EsuSzFvXLVf7+g9yn+Jj5fqstFCW3oc622JYY5xO5A9H1ab/dl27TYs5AKGTyWT7Jrkxs
RE5ez87INDLzwYlgsAR7yyS/SLlyvVha3zrrCh1l5eXMsMOxykC5vtb2RIYxZVQfaL4zX1ffRaTv
9Wf9ALEDK/leQz2mlki2UB9CZjI8CC5XNqX8/WIIhkmMyTkdLtYHbpdn1OJjKvx2vKj8htYE2s1H
UosIv0LvZBiDm5MFxkhOW+LKjOPhghGDjAGQxjgeyWMvzYzbwNKBbjY8Pl31OYMJuBdki/LTDpAv
BctpAgmY6boRpPWSf2I9mXax0Qjxi199PAMDxBi4oMaSQ0dtZFfBK+6fNp0bK6/2a6DiaWeos8eg
flARqSKgIEQFJ1DrV4cDG0Dl+aeyXJjdGBxxDmiJEVMxdXDNuvSClN180/sgs9l2KUYLNNr3hwhk
IlGqxtzc33yiPq1LlplIs9TAEekeSuXcgmyS1rxY2qMh/ujWwEdT0McdQmFZcrn5TuLwDIdyY2EE
sfd0So+2ff4bPamSxK0ChDn2FBUcKWIHr3j/xyFl4IcjmbDszkgKtgw2P2uSRbh3ZMrPJ1ZGMY0/
fX+GD7ZH3fBnLY4I2PxwB8s/jy6YT7y2g5hP7I+PDZGT21s+07Xz2QRBuy1mUTC2ngLnpKQ0D2b3
yBmmwESQtK4EZNWWst7nLoYBKlHptwOR/GSjKJMmWCFSNscWz0jyAfG2DNUWGDtfx+sg/0yRujhU
2Lnff2aP5ie71qNdhWpQB/I3n2HjDP6Dyt/H8QGnVL46dwHznY8yTvBX3MFGG9RqQESkv/vuQLa1
rw6hHh2f7U2mq/Fq3zaCeKhdGPIvyr1dT3zQT6kDygcVgMIZSPb5dLlCnG3WqbIXtCCFiisg2a0E
V1dk1nPO+5V391YBQUt+RAM6NQpLPL+NcTPqUjoef9JVm1pXCBH5Dpo9yc814sKuQk4QSaWecPr4
e6t6yhoAgrSvlX6mXuwDRsm0nLmo5cK6UxVarWsOBiksJ0spkICvCyHrko/Ow56yS5g++9e4xpVz
KtULUDQw6dPBlQ/EknYc9Khrr7RHSpPzjt8lus67jcbCWgxGFmqBTrmZ4LhcOgtsWvtAar3gMrAB
ehpHzVKcpsuyVNm2HbHRo4fWoDto1UU7ZnnuksJj3TBGlr0X3uKER7T2Y/TY0cUKBPcrKaTMXIx7
sNx7vSVNAcFld7dZjRzAo460XBBOkELJ3YPF/JZxZO6fids7dMbdzWbytyv+AwRps/UsdwsMkNAx
62W+iYgBnmt/MpDPXjKpUMsb5oZVzHWN0hG3Misw5hghDbG9zgvToyfDU62XPyIL/yvR76+Pg0SS
A+CLiOzCj0yYW86TUy5ZsYyYjRzONB6F44Maledkt4/iTS3yYKs+RanOTJIBict0cTJnl7xgf1Gk
QejduC9muvS1GGur3QI6SLWsUuw92qkFHiRDCOqwcot0yQgpLvedfednMxyReEr9+zcqzNhrTTPx
7MvCG0d5pwPpm5dHyrazXZDmaxTmnlyxokpBAYHMjNWEgKcFPJ8mUuRzVGNWv1SPySLlYi/hYi1z
4pbxzt0ht6CfXT/LYp58OsLk+A2JaXDnXWZBVjbWTqfxjiwRgAvdr7y+iL4jMOZbJDUUdk7RtD49
UYEvWi/48fW5kVODthkqSmngIiDLGdVxL0f5UVnT5m6oojLGROoohPR3xmE7vMmg3SUQ97GjRIHq
vlfMOWc3KMVP2UBjYCYdg25Nsbi0JFH4YSsHCDjC4GJ5UWDr/RCjTZ1z5qb0/zTUlcd3wv9+eVaQ
WzfHcSRlV5A8OlSWULGIDWuwWT7pBWz59DwDa1cjPc2hdcyXc0Ifxd4aCzdKBzE+vGDeSskEx3O6
J8eSKHn8m76EsQHjw60H5rkKCp6wMReXSJG0UUp9G50wdEbHDRfhCl0IFgSEtEIIOTLUMyq0LK6Z
9ts2qWeqJO79lUCSSyxVHvyyjk2Y1+A98gjJ6tBLnnCHgvXWRPLR4+tp0NVsaapJbVJKuEURWoJo
ocONBxTYmTXmoTGnoYdBi4mW/epTcKzfKN9voprTrwHzy1ylBB/qS249Yg8UNrN0LrS1TdkEctQj
HCt4k9cVgkzv2vC46mqlWm3oFVPgYgjQrIK4S+bqv/S8Go4ApjPr4SrEPU0ZyP3fqgHsKQWyD+xo
RhBh4OBaL/MgPK41irGV9TGDO/+Ch7d0zIDHuP+gKLO7izr7tx6NSfbtNAnHYwSfS/dEdT09vuDI
w3lVo/qCB9VeIbvFQmT1Cd0cv6WNskZH923OUg6bOuJuz6R+U1lcy8HhPH+Z1dQv4qWt0e4Q3RVx
WrZJgTa4Ln07Rm/nHU/Z+QnNmdCJh4L+i3dATsqqr38MBxovEVVvbA08ox7ZW+TbQcoFNy+GbfIK
tWXvG1bHk42JbZ4F1NFQD9v7hASdDbdLHNKsJnx6/QcD7YMux6xUBGTsdJRA9lGejyjuOPROZcDh
hE/6Job6uRHt76DSoHhELcg8DLExV7Uu6NzrtpawBD/DHdb4R6qq0I3jcuSih87y0frdpbTntMcA
5koxK6Vrmj+qk2wL8esmHZ+jGCdJOQVGD1PHI0LdL5eKGi72Pt3un7tuP836E3M50ZL0V0Z1duRH
NtAq+fUJ8jUnzD3Dbrc/OypAQkqEJoK9O+xQTKWs9gXwHDn+jMY7xKU1bAZxPfY8FYGIO4o2gwaC
Cz2X3uALaKXkg7leC9tR6pAmdAFOMeegqzixyQbxIlrl4wfTlWxJVVPaKk/RUyw54kQ/vPoCQbZy
1C/nINKHJwAWrh/OnX1BZqOXeg+EV2jUZ2RSVKYY3COe1CWqppwMALRrWjq3uK/Zz9rzIZS2zc0p
KgzgOxbBekjPTVMxt9Iivaa2GYRAzNgJDH+psSzWlQxfVMVjjpxwlRHGRb78iJ4xMUunDcyuvXbP
RCkk63MzkRojvkY2Pn9tQKNL5pzyOF3fY6ab9whXh336w6OOBW2+cvcEvFhG+Xe/ggWhP6Z1VNcF
Pbxvxws9XB9u8VBHU+4Z+1vpltd3UsK6fwTPFgaeYKMOTPgdb8aGwZB5uXXgSC294DjbYpoqU+SS
saR7aHLUOWZUQPx7/pkfGchRCJ+iOCkvidQwILBKmqu/PK4aBF4TX11YskjVbdxvez2P7VtFjfmW
wXgnQjKxFJw04JvhYjYhWzgH1XhU5nDMB6yPiDv+gvimheKWk97LC13BMX8u/8twcqKIhMKtNkf+
x3/bK4LNOVACIF7lyl2czF1k0W0lUm6WVlJZuPpgM7wvuBDEdDurx01Qe/56EFsvZFizQHIgxO0w
CycZz9SeEV09IG4Fr9j85P452RKtfGmSsrUZUWAac7pNYNT4FjP/nsgfBcl0EEwinn42eIi2PgcB
4YCyvV9wOFMQdFQhItd86+XRSKBgBm6WFDC4oHVXFFO4meZFtk3DUyTDs1UdlTO1MzheJArEiDhe
Na4520ipmBFaJQ3Q0D5VzJvm2oJOs5nhTnbDjzVfsfw809GcRqkJgQnNJ/h/kdql91kImf1Yv0vS
fiIVnm6ivhJBvxVtrbqV4pPRrnz3w8a0EHq3H92ZP8jQXXPM+RqjXWL0CZule8m3TmpZFVXnvFyu
Qd6T63rnJ3M87zysIKU15gynGqILliJiMJADPyRjHJDT+Lptrw4ocDH/eHhwbQOSx/YIPVykCl8K
irJr/rK7tU6Qjh2V47PiLx4/wx1dPwptRC4apBqc7XX4qhoqbMArpoZYM24TBYYCalqiOmN/eEaB
clmbiLyEFCC8JWXOF1yWXKrCDZBlGGMsc2jrjbrTi+wFkkHE92ccaG0ZOSJbSHPt82M8wB1gcvUz
xayArJzTfNlsffK8yuOs/7rcNffYQ71X61AGUX9/Si0SlkpKFIItFo8Z+8F2Bowgg3vjs6ROEwfL
HZtKMzaPoleEWI4PH0NpCYyhBR91Ov6ftBPm7afuhhSS1f9RJEwV8KrC1n0EtP/o6bU4KL/D0Ax2
/P4aDiyPlHkJnVN3dR36DEEjYRFayBdooNOn3e3Ga66XWhZcp0b2umQKK2f7SgH9ZQEhxEyJeMhX
ksi3J+QSVCKV8TCa97IY5hPp2pS/LY2Rv8ER3TQ3/5lWOET4Bl5EgwTx6df+tBcCIEXF8bIM5hTr
th9xKuP3SCK9/pumKdprVOTRkfS9V6H8PWgf6z9Iwxyvg2sVimL4eJgICzvpQIN0oxU0g+kbnu/Z
VEx/U9CeIEmo+UnHxK0l/ImopVoYFpEHzaXyYumL/G0HGe3H2ZdkveiyLrjSIG2XvI7y6wONxa6Z
LkZD4vp8qDV0N3u5+9uqp3z28fbzYl8cYh8AcTuUm1dMtVnPC4RJoNEncqZa0GcrC+UdlZE2JHYU
FuOG9cnz07cHeiGgeXNnm+DVTUd2GVvl832f9A7X7YKINFb6v2hCwn/HBO2rrK6/WvoRAm1M5/9w
E/gFLQKj3MSebIA6Irw5i32KiUogsClI8OsYjjRfwnVtAbDPp3MtZcET1TPK3Otk5jUp11jOlL9K
KZOHQF1JTITuyoMermTOaX4f5mNpuUgYB6qPo1LCjJmvSPQNj7SsR80EtQ4PbH+kD1VFR/CgGTAt
imTuMy0tPNSKT5HaX6+QDUF3LscwVNz9+s9t1hm1y8HG7HPLTD9hRYNVvFvaVex8LM0tWHTCVMbc
TETbR5KDHHalgJlHYbNPljcHVoSlg6hSIWtIHA/ypdgMj8eAtUOKZZDgx9j7NpHZB3dnnSJKFSqs
UkR6wK1UExPX/NHIqNN5mMugue9JNT9xihCpzOg0GcUQ0MmqJUSZDN6kHupC2yp2fsU5yUwRcHU5
/gPO76CcKWZdrpYnegXmAB8vxfeLpntHXBxPM7TjpWbnFicdlTS7BjVDn8ll3Rz48ss8mqjhdV+8
gD9WUVu7Wj7YtHKSRSIH4BH3hpVLWLnrU1Upy2AmxzrB0+wjZ3RqGHOkQUpySQRpRAFUfU5XXZtr
YsfRMA/4noLSv+vZFALBDW8r1uF3KxOa1SNmsGtHFXialTzayCGAau30egHypi3459LMprwxKn4u
xBpEAZJ45mfnhWWZKrZh/gijA6cdw+5IYMAG5FgCpXM1QGiwrupRClrts9tShBuMqJGxNECcs859
kubw0ItPjdgD+ZhykcLT3nP0ouLZeC3AWgEK+BcackUkmINjxtemY1ftzJXvPKnrXfG2QYzUx4NJ
NMSDgbsEWrNFi96weVarLUjfRVtHirQ4WWnCoDBKwWS0mCFOx4bm+cL2YKM84WRwufeHUNH3c2D/
XzsVCLhtGA6j5uGq6qgedT2cqRXCl8gLuSJEY6xp1irtFoPNIT+EMq01H4TJf3YcLyC5m9ROMmGW
qLdU7GqDBsFi/bk4ia5sPb0fet1h3JfAp62RijdeaWLvWV8D+nU6ifgB8ZcIZ9UQSX9hnDfaIm6n
bNoBqYWTQfWuJb2po741M22Lw19SO80HUqWOj1GCpVxo2AmglgwQ4QJ/w7eS0gVjlp1tTMT+bako
JzTu7UaEYD/yLCvU7UqzUd3EplMoWm7tAPGl/vo6jIdg9OceRjUw2H6PpEw+AdfyweEOdYJMbE7J
xl5s6NgD/6Uh1fOviii6KpjsYjqD4rkQXxCGlcaspogEskIBaBX1v5rnO1BeSvzptj9MkEytYxMb
ibpIPR2/FndxFMRLMpLzmpXUD0A8mzb7DgY/coNYAyiu803Ff9SQsus/vRV5xQlEipsQozchHz0y
nfWI4ZOZyZSAjZBWSPauWrnQhZ73zax5eLkZwFpSttBEKNhyW3SvVaucymaVsgfB5ZjYz7nYOGOz
r4IBn0x8tX4gl423NpFMpwJqMzbvnk7rUM+gA77GKdaP+Il6EcYR+QWfQ5xMrLYYTi6AKpRYuPz+
0A1lUnM3QMq1Mk8A127JOGCqAZMSKAziHxC/KIqc+V2lFjtzKb53cjVVuFivyGqNPFZsUH+4mKqg
iSxP2jWtIE0OD42w1188q4AbyfCHOyqhGl5WUymqz/9L8v+nwT7r+pssTvJGDCqOkobwRgzw4lvm
Pd3v2YO+LoSgnf+9jh0FKVwIFyXZ8NnFGrreTUG3u7MXvBS6bqxwzMyQUsu7t5M2iZX7Rn51+nEo
YOHSO04sshq9BV7dXSsmq86nfAL92P0lWP9BQmj9/qxvRmbZnq86gDEXYrA9IzTgzSc5mL3VWs47
a+UVfDZA04of0Ff13YZTB7JeFkrHosYOTeab6eGB3Oama0lTSs4M+w9J5c4CbRkXdjC7iE4ugkqx
5+RYpd8u0y3cuPK1XYKJFFKxIFlSASEY/HzkEBsWfmWwy/MIQNDSFx+nGpqQTQgWhvZxgmVrXWQd
jkxez0rBM5F3PdaYnQpeQWAUuk02em4h1whZIscAG6WBcuJsJ9YaEm7FymX/qbzUpc3C0o7zLLr9
+huBMb62VvDUcOAhVb5iXFVs5SR6cqdmIBzN7kZ3exRAgKaLeYGWKDObiTEH7mNnF/LRMlbU/iae
ehz6COWcQrCDRiH06D7MocRht8u0YgaH64cF1jlQdNRbZ/95di3BFlkjPH8SdtheuvPfGqe0txPt
1xCoIM7jbXva0XP3xfsAJ0H+dCeRPnNrneSgu4RuhbCEbvLX/xaPcDB5LE7Gc8B0hRT5QmMTjgTu
ky3JmPfPFmKiFmqrcmeqa63rFYmzTP99Gt4pSieaLfBfq3TzaWOmVtDkmXYl1MMfhNMOPn7/JeoV
nHRDQWjSS6kzUAuwNYywKgclfd5PMHy0fI3tthuQ/t+H2P6LXeZvZxvqX0yNx4JefAHYoxYW8IUC
SmzoUmPBqfoDrK4taTNZAJkD3lKhXy0rgfU7WOGepGkW/fJnImT/9OQ12Y+zLniw6omQQNQ2ddcN
8wPMV9H0zbZtjZyAeAGVNQZ48K8V0Abw04dyA+nPqo1YkJCwP+xcBi068U9U3Imb458wIwQwjaUa
y6jOGQ7Yh/jusgGb7irid0BnICwSLGvR8kpkANswBdjjHN828c4SPp17a3agkk43gJyBV69inrGg
9O6XP6CQ79JmQeJavdyXn6KwdDYQby9nn1Wf+GbHbCBzNgkBhktgS60xWM6Qe46dg7Add6TZJRd2
xuSulo/K2EAPdwVgcNNK3767WEPNzgq45qXnsQzVvGqH7RBzqxnQIYnDkty0oO42VXlHcUqbjTkk
tFKERo3ii8F2P2G5jyN1H9n7AWew6tNTv8MzOrZ1SHhB5nVz33jarZR9zVLfy8WUWQXlm7m4N/rG
TL2O5oNIkMK4Ow25DTBbXD6uex5+lbTDSRvyXCZWZDUy9+qxhywtSZ803qT2a+x3dNP2I5/12kaS
JWR529PzjEBnT8KZYgh3op5A7ZknftinQ0cWDk8omzxO51HXs2W2Ne3jAGVVwK0oZ+VDVyvhSTUt
LlC6eBBA/PNtmOLNetjuCvGYMw+yFQhWzGKFpTMEP5zwKUNsI529uJbrNqoeADWpthdslEJ2dWdO
+M8m1J8aLsMTcf5ay90cW1dBDzf9GPCLeHVSMk+qK0Mrdhdgg0r2xG8n4tQgN/ciNulDNw1vcv8X
WDKx///9iLqDBtNpW5B6E3kkeuKINYB37fVPa2fMuDoeFiVwUZGAVCpxTlO8RwJOPkdICsGwY4CF
OqF/pG1ZbftnqgxwC+fV4vGab7AwhLyq4m6BOZbAEPZiYgynNccZXByPVhcBbhicYww5hwcKuohW
+jakJJqseYLdLMVEzoEg65I9MCCzrrFNe/cdtiUlMmNJJcflbcNyCWKmlzPr3CGdsgUy09lxA0hs
e3s5/FJtzhM9THara+cM3SdJzjhY9diiGepnjMV8zPMXnAV/Yr6kxulNzdikzWmJQvQQMcaF8MfY
3STVATtHIm7tqNcHDtGAp5InEzmBzdBcuY0zRmd89mCD4QvoLK/9GEvfpAn6vFG73iCrYPUEvQ1o
IdPjbzEOpgLoJS0Dqh8/pwMVs0npzUq8KFJkak7tXZyRwhDZ8CQxoXUMI+7vffoHrQJz6jQYrl/b
LMlVky2vqxsVfaD9nJNJ9yJd+6khOXjsZHzqPGpdJJYx1C//9Yy2ZJ+XsTlsAPhduICNabypouH9
myQxg2vSU8UFpmlhCJL3bUQnmVwVOGNImVRvjlUlj6ZrmIPHzXh4raywCqTe8srABe0E4jLdWacz
2tCl9HWC38tzbbNBQLkpaM8+WuLkvLM+a987eeqtmSnH5GKxWonZQaF0xZQe7I779NmKziKoxBcs
F4/SermDcy2uTZWjhHhcFgQBk6vx4RccxhObz7VdAG9gEkAyZN4c2Gh7J1M1eRmHeo4cYl6/mY/F
D6P73awxhyybEY0xi3gb0qCXqJCH3GwAZzxYfiKTgsmYs1+xvZDcLgsC5SdK9t+yxf9E0C7ysKPe
xJPu219LmzIDUdPwvdre4uCv5D3ekI7Sff9dW7FGD5JlnvO+9/8MOQ9ySDYHLB+cQZCCnsvFFC/K
nBUuhf/Ec69i38tMxCE3DY56mxJySThT2JGCIeEkhQIOr97GMqGVa0BxtGzoNgk31VUhHR5iRMVk
9vpbgZvWMVlvT3y1YiHD9jv36alJB95Xxym9LNZFvbZ6PGokXT5GjHnOzp7RCWQtODXHoVdV9T5t
ZxCGGGJExKmXRN/Chj4NYWhK+hF20kIkgqvbqBTW/jiKdOH93phJcd3N0gppM6UIBAM1WS9iuEEv
BY1kCH5r5dcE7c9e9HAfVMC0lxv5JXkQcma6Ig7xML3/ZGkWT0m4V61fv+PSR3+oW71KA6YDjdiT
UMOdTy67Cx9hCOy35+hn2+l/xAe1jIzNnqhoJ+myRcY57TrmY8XvRWzyiO40EUoTt41iysEELA4u
DfffX5VJjf6Pn+wCYnnCviTeS4jJHsYYz2XNEzBUTf8Kf9ZYTi7KYbnKg0QcsOumCHAsNigAWUau
F8R0XvZPzRUUgszVWLA7lp2ob6W/qRmIV8tHYd3asgmNxVk2qk9Vg8vp5uDBepOxnndDTw86DCPW
Zz9GfMqeQQknLDRqb/o+na5Id/i05KF/sEtmZ9qw2WX0FCRKdUer/bIs2YL5XVNjhDM1HJGt3PSh
H8SPgCF3lHdeJH9evuyNsSHbz6EFfW1eSRpKNrQueHYMBKEYpiivaBLFJ1HlrMAU0GjVeu8+2rRn
S0dOHGGoS6QVzTupW2D+CLYZftLaDX1+OAcP9nuzMrjMpICH5PaYJkJ8ahyhgaXK/yowtMfsRGKu
m72Z6HzRtZnvZHyuXTXBV7XbJwR46fRfo79jcD9oOphLGVsXkSLvg8WsSIpxzqluapaZD9mbsg1J
awa/Zu6bG03tp5Sajpoy6ibZg4oHMKFMJUxPg9GSYYys6RNQ/lif2G/Ln9hLz1a7Iez5Zo8RDghu
0x1KUue49ajds6xFfH2XAEHvtSy68kG6o7lxiyzfPvSgEDHBslQ2e74lETIcdXqxNj3OheNJw5kI
hL3Sd+qBAiMasdxkCPro6RQrmWntsnDD3jBrG+A8R9ewOXOv4mRGGQFLyNREjbQK/OZSRwMC6iYe
EHRRcMuaRd1nO3wyxWP7sKdtXffRS3Bpc73hAMp5kbX6WugHjw2Tu9MA25uBjtUgRbo4gzwgXVIx
6Fd1DztBw+R7uhY/6XvUHvYolXqTH4siEVsOY0WSTgCMnvh/r2Sa69nouQuhxeWDQeY+04nGMJRr
YPXgQcmNwwW+uCubQJQj3dPoEvP8NJW53mXHe2qFElUFhXPGi0nvcfFZ6p8x4NMjCeiduMMQh5Rd
hjVLdMVxDUStj1KaYbTS/h9go9Y9r/jiZXCh71xcz+Q3J/KYqZO2/LwpuDvP8L/Nfuy+IEcUelnc
yzGtIb9t1kQdBdlG5E6QWmmkJu1+GUv8LOZgtPy9LQCF5hbQ9lDvCH+1Lcb4PeY1YM0q3EIhbjzO
SvK8JXUyXFwwknwr7egqzLD3Kf7UomdIwsl+agSa3qycpUoxziVchQQPMjQeE4yoMIhwc4/0MsZN
YuUjMUIWLnVTLQ1pceTz5bw/Rlzw3NZaf2I6pT0+V1IyJSvpmZlSi2Lb1lxk0jNVHlr/ETZYjQGn
YoPEcLRvD+oH0VwZfHC6GxagrvAcxbwePUsJZxUDYHEH9RIN5iw05Un1jmNLtVlQRJCv85WBKKst
dU59/GACyqbnIm5YXMXJfrxZqkdI0N3TK9OGxf7FMnRi10juNsMfwGvBuy5m7sR/qwmzY5icdrqr
4HrEqoduLjbmsedxpVomM+CPvpVjYG6Yfn41f823XS7NUzU9rIHHwIMPftbaSLnronyJYiMW5C//
/EwV6L8X/lBH7rflhNH1faK0u1QkBnj0wTPZc97RAxe02306msul9VKc0hbxQWoZhwIfhnDkEVSH
Y4ckSSB1mYX4gKkKnSoAInnfVsejZp4kIUXXEmt/Eo+EMgJtMFtYi1UCj1L6ZICsQ9Rfs+pbFcE7
lv+mm7xVosXjgD6UWlUTS6fTSzai6HC7CpKQX3cUwm/dISozgBhOzxhihjRqkHpOA1jRlUklvjcp
lZKfqPpeldMRcO1QVFIzsviyjs4QqB2n7SjA3/liu2kNsfpYurYOHvXPbAzEgthV6JjkvhIjISIR
Cxgfhlaq8YNUAITP3YqhOYATgXnFe+cfG+Exlbp/ihq9h0RXdfK9Vocrg8HZpnVxo+i1l6IdK3L+
I2in6lye8pobA9a3EFhD32/ODhqippzqfQH0Nto6hTmyrpbz/BVXgMg463SFkeMGrrmiRZBitpoy
rfMRPPW26MMz58W/hU533d8XuH79plDbXs2uVBhSPLCCPQ6nGb6nDyAooNlSYlbMXdnX1+O8TDVJ
z0ZCJDFMWBo8sGSR9dmxbf81uuf78JFBVui0xSEl2CTtODnAeAnbzBjzWixfHv5iU+Q6QXkrK4Y8
kLge1zF3KZjSW02soFqXLgXaJDTSW7MdCguQV52WeMeN6jjA+jqLHHnziHcugqLfLYbLBRGmBmCO
QfZKGsQ4HvjYxSLwNfpdViBzCXj+CcsMzIh7sQGsM8G0TMa9YoI9gO+WZ308wL20OPClP0ecl0ZN
fEnGPorFVMg+plnBguOks82A7ohCHZT1q/3TA9BIqO7PXIho/zw5FzmiS3CLgHwsyzjcGM3N5T8x
2LKfaEXUJzAsNF5itGBvLA240tBLI8nYcETG0EYTR0FQO9b7THgMef+s4ra10FwkThIVvWG6ISr1
z3Dl9RdcBKRJOEFpAkRhOQtFIMcg8rKiqy9aGMcjje2+xDPSqw6xkLvXi/9aZNe64YLxAzX0PySd
09m5kvKV4VkIBg==
`protect end_protected

